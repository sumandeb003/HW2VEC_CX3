//****************************************************************
// TRIT-ASIC Generated Trojans.  The design generated below is for academic use only.
// Please cite the following if using the benchmark provided:
// J. Cruz, Y. Huang, P. Mishra, S. Bhunia, 
// "An Automated Configurable Trojan Insertion Framework for Dynamic Trust Benchmarks", DATE, 2018
//****************************************************************

module s5378( GND, VDD, RST, CLK, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat, n3070gat, 
		n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat, n3077gat, n3078gat, n3079gat, n3080gat, 
		n3081gat, n3082gat, n3083gat, n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat, 
		n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat, n3099gat, n3100gat, n3104gat, 
		n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat, n3111gat, n3112gat, n3113gat, n3114gat, 
		n3115gat, n3116gat, n3117gat, n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat, 
		n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat, n3132gat, n3133gat, n3134gat, 
		n3135gat, n3136gat, n3137gat, n3138gat, n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, 
		n3145gat, n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat);

	input GND, VDD, RST, CLK, n3065gat, n3066gat, n3067gat, n3068gat, n3069gat,
         n3070gat, n3071gat, n3072gat, n3073gat, n3074gat, n3075gat, n3076gat,
         n3077gat, n3078gat, n3079gat, n3080gat, n3081gat, n3082gat, n3083gat,
         n3084gat, n3085gat, n3086gat, n3087gat, n3088gat, n3089gat, n3090gat,
         n3091gat, n3092gat, n3093gat, n3094gat, n3095gat, n3097gat, n3098gat,
         n3099gat, n3100gat;

	output n3104gat, n3105gat, n3106gat, n3107gat, n3108gat, n3109gat, n3110gat,
         n3111gat, n3112gat, n3113gat, n3114gat, n3115gat, n3116gat, n3117gat,
         n3118gat, n3119gat, n3120gat, n3121gat, n3122gat, n3123gat, n3124gat,
         n3125gat, n3126gat, n3127gat, n3128gat, n3129gat, n3130gat, n3131gat,
         n3132gat, n3133gat, n3134gat, n3135gat, n3136gat, n3137gat, n3138gat,
         n3139gat, n3140gat, n3141gat, n3142gat, n3143gat, n3144gat, n3145gat,
         n3146gat, n3147gat, n3148gat, n3149gat, n3150gat, n3151gat, n3152gat;

	wire n656, n1146, n1892, n1147, n1118, n674, n1114, n1148, n1113, n177, 
		n1111, n178, n1119, n1911, n1120, n1908, n1121, n1122, n652, n660, 
		n1170, n1169, n1893, n1228, n1888, n634, n614, n187, n1222, n189, 
		n650, n1117, n617, n657, n1223, n1007, n1123, n626, n1115, n633, 
		n621, n1124, n655, n1125, n1126, n665, n1151, n1150, n632, n1152, 
		n1127, n200, n201, n644, n1204, n1110, n620, n1202, n639, n1207, 
		n615, n1208, n1205, n638, n1200, n1128, n1221, n645, n1129, n637, 
		n1220, n1130, n205, n206, n1224, n1217, n1225, n1198, n1197, n1900, 
		n623, n1157, n1131, n659, n1154, n1155, n1158, n1159, n1156, n1153, 
		n1901, n1160, n1132, n1161, n636, n1165, n1133, n1162, n663, n1149, 
		n666, n648, n1164, n672, n1163, n1134, n226, n649, n1218, n1214, 
		n1219, n1216, n643, n1215, n618, n1210, n641, n1211, n646, n1209, 
		n642, n1212, n619, n1213, n1898, n1186, n628, n1187, n669, n1135, 
		n629, n1193, n1188, n1194, n673, n1166, n640, n1136, n1899, n654, 
		n1196, n1184, n667, n622, n1185, n1195, n1183, n1167, n675, n1137, 
		n1138, n1168, n676, n1896, n1172, n653, n1139, n630, n1173, n670, 
		n1140, n1174, n668, n1175, n631, n1141, n647, n1171, n1176, n1897, 
		n1179, n664, n1142, n671, n1143, n1177, n1144, n246, n635, n1116, 
		n658, n1876, n1180, n1902, n1192, n1189, n616, n1191, n1190, n251, 
		n625, n1145, n627, n1206, n624, n1181, n1182, n661, n1178, n1203, 
		n662, n1201, n651, n1199, n1112, n1771gat, n256, n2446gat, n1226, n258, 
		n2021gat, n2084gat, n1227, n2102gat, n260, n2458gat, n2121gat, n2025gat, n2044gat, n1363gat, 
		n1433gat, n2179gat, n1332gat, n2029gat, n261, n262, n2266gat, n9, n607, n6, 
		n681, n689, n688, n690, n694, n700, n699, n703, n705, n702, 
		n710, n712, n709, n714, n708, n697, n695, n717, n716, n719, 
		n722, n724, n723, n728, n721, n732, n733, n731, n720, n718, 
		n735, n738, n737, n741, n742, n740, n743, n736, n744, n729, 
		n730, n726, n727, n725, n704, n746, n749, n701, n745, n751, 
		n754, n755, n756, n753, n760, n762, n761, n763, n759, n764, 
		n766, n765, n767, n768, n774, n779, n781, n783, n785, n787, 
		n789, n791, n793, n773, n772, n796, n794, n792, n804, n807, 
		n809, n806, n813, n771, n814, n815, n816, n819, n778, n820, 
		n780, n823, n782, n825, n826, n784, n828, n786, n830, n831, 
		n788, n834, n821, n835, n802, n795, n790, n838, n839, n776, 
		n810, n818, n775, n777, n805, n808, n817, n812, n811, n801, 
		n840, n692, n853, n684, n858, n857, n30, n29, n28, n27, 
		n25, n15, n10, DFF_9_N3, n869, n836, n871, n870, n837, n876, 
		n875, n844, n797, DFF_99_N3, n803, n878, n877, DFF_98_N3, n846, n880, 
		DFF_97_N3, n845, DFF_95_N3, n882, n883, DFF_94_N3, n693, n885, n886, n884, 
		n888, n887, DFF_93_N3, n891, n892, n893, n890, DFF_92_N3, n898, n897, 
		DFF_91_N3, n899, n706, n901, n903, n902, n900, n905, n904, DFF_90_N3, 
		n907, DFF_89_N3, n908, DFF_88_N3, n909, DFF_87_N3, n910, DFF_86_N3, n911, DFF_85_N3, 
		n912, DFF_84_N3, n913, DFF_83_N3, n914, DFF_82_N3, n915, DFF_81_N3, n916, n918, 
		n920, n919, n917, n922, n921, DFF_80_N3, DFF_79_N3, DFF_78_N3, DFF_77_N3, DFF_76_N3, 
		DFF_75_N3, DFF_74_N3, DFF_73_N3, DFF_72_N3, n906, n929, n930, n713, n707, n928, 
		n932, n769, n923, n934, n683, n874, n936, DFF_70_N3, n680, DFF_69_N3, 
		n868, n938, DFF_67_N3, n855, DFF_66_N3, n859, DFF_65_N3, n687, DFF_64_N3, DFF_63_N3, 
		n940, DFF_96_N3, DFF_62_N3, n851, DFF_60_N3, n850, n849, DFF_59_N3, DFF_58_N3, n946, 
		n606, n879, n848, DFF_57_N3, n824, n950, n952, n954, n953, n951, 
		n956, n955, DFF_56_N3, n961, n13, n958, DFF_55_N3, n966, n963, n967, 
		n970, DFF_54_N3, DFF_53_N3, n974, n17, n972, DFF_52_N3, n978, n26, n976, 
		n979, n980, DFF_51_N3, n983, n19, n981, n969, n957, n968, n962, 
		DFF_50_N3, DFF_49_N3, DFF_48_N3, n960, n965, DFF_47_N3, n822, n989, n991, n993, 
		n992, n990, n995, n994, DFF_46_N3, n997, DFF_45_N3, n1000, n1001, n1002, 
		DFF_44_N3, n1003, DFF_43_N3, n1005, DFF_42_N3, n1008, n1009, n1004, n1006, n998, 
		n996, n984, n860, n1010, n854, n988, DFF_37_N3, n829, n1011, n1013, 
		n1015, n1014, n1012, n1017, n1016, DFF_36_N3, n959, n925, DFF_35_N3, n964, 
		n867, DFF_34_N3, n866, n971, DFF_33_N3, n973, n926, DFF_32_N3, n924, n977, 
		DFF_31_N3, n982, n927, DFF_30_N3, n865, n985, DFF_29_N3, n864, n986, DFF_28_N3, 
		n987, n1018, n863, n842, DFF_27_N3, n827, n1019, n1021, n1023, n1022, 
		n1020, n1025, n1024, DFF_21_N3, DFF_20_N3, DFF_19_N3, DFF_17_N3, DFF_178_N3, DFF_177_N3, DFF_176_N3, 
		n862, n1028, n1030, DFF_175_N3, DFF_174_N3, n1032, n894, DFF_173_N3, n679, n685, 
		DFF_171_N3, DFF_170_N3, n941, DFF_16_N3, DFF_169_N3, n1039, n711, n889, n931, n933, 
		DFF_168_N3, DFF_167_N3, DFF_166_N3, DFF_165_N3, DFF_164_N3, DFF_163_N3, DFF_162_N3, DFF_161_N3, DFF_160_N3, DFF_15_N3, 
		n1041, n832, n1042, n833, n1044, n1046, n1048, n1047, n1049, n1045, 
		n1043, DFF_159_N3, DFF_158_N3, DFF_157_N3, DFF_156_N3, DFF_155_N3, DFF_154_N3, DFF_153_N3, DFF_151_N3, DFF_150_N3, 
		DFF_149_N3, DFF_148_N3, DFF_147_N3, DFF_146_N3, n757, DFF_145_N3, DFF_144_N3, DFF_142_N3, n1033, n1036, 
		n1052, n1055, n1054, n1057, n1059, n1061, n1060, n1058, n1063, n1056, 
		n1065, n1067, n1068, n1066, n1062, n947, n948, n1064, DFF_141_N3, DFF_140_N3, 
		DFF_139_N3, n1070, n1072, n800, n1071, n935, n861, n873, n799, n1069, 
		n852, n856, n1073, n798, n843, n872, n841, DFF_138_N3, DFF_137_N3, DFF_134_N3, 
		n1075, DFF_71_N3, DFF_133_N3, n1051, DFF_131_N3, n937, n939, n1077, n758, DFF_130_N3, 
		DFF_129_N3, DFF_128_N3, DFF_127_N3, n1078, n895, n1081, n1080, n1079, DFF_126_N3, DFF_125_N3, 
		DFF_124_N3, DFF_123_N3, DFF_122_N3, DFF_121_N3, DFF_120_N3, DFF_119_N3, DFF_118_N3, DFF_117_N3, n847, n949, 
		n1026, n1035, n1029, n1083, DFF_116_N3, n31, n1040, DFF_143_N3, n691, n752, 
		n734, n748, n750, n1082, n1086, n1038, n739, n770, n975, n1037, 
		n999, n32, n1076, n1085, n1087, DFF_115_N3, n1088, n1053, n1089, n1034, 
		n1090, DFF_114_N3, DFF_113_N3, DFF_112_N3, DFF_111_N3, DFF_110_N3, DFF_109_N3, DFF_108_N3, DFF_107_N3, DFF_106_N3, 
		DFF_105_N3, n33, DFF_104_N3, n698, DFF_101_N3, n696, n1092, n1093, n1091, n1094, 
		DFF_100_N3, n945, n1096, n1097, n1099, n1101, n1084, n1100, n1103, n1102, 
		n1098, n943, n1031, n1105, n747, n715, n1104, n1027, n1095, n896, 
		n881, n682, n1074, n1108, n1107, n1050, n1106, n1109, n942, n686, 
		n944, troj47_0_n2, troj47_0_n1, tempDFF_46_N3, Trigger_en_47_0;

	dfxbp_1 DFF_0_Q_reg( .D(DFF_33_N3), .CLK(CLK), .Q(n656), .Q_N(n1146) );
	dfxbp_1 DFF_178_Q_reg( .D(DFF_178_N3), .CLK(CLK), .Q_N(n1892) );
	dfxbp_1 DFF_177_Q_reg( .D(DFF_177_N3), .CLK(CLK), .Q(n1147) );
	dfxbp_1 DFF_176_Q_reg( .D(DFF_176_N3), .CLK(CLK), .Q(n1118), .Q_N(n674) );
	dfxbp_1 DFF_174_Q_reg( .D(DFF_174_N3), .CLK(CLK), .Q(n1114) );
	dfxbp_1 DFF_173_Q_reg( .D(DFF_173_N3), .CLK(CLK), .Q_N(n1148) );
	dfxbp_1 DFF_172_Q_reg( .D(n30), .CLK(CLK), .Q(n1113) );
	dfxbp_1 DFF_171_Q_reg( .D(DFF_171_N3), .CLK(CLK), .Q(n177) );
	dfxbp_1 DFF_170_Q_reg( .D(DFF_170_N3), .CLK(CLK), .Q(n1111) );
	dfxbp_1 DFF_167_Q_reg( .D(DFF_167_N3), .CLK(CLK), .Q(n178) );
	dfxbp_1 DFF_163_Q_reg( .D(DFF_163_N3), .CLK(CLK), .Q_N(n1119) );
	dfxbp_1 DFF_162_Q_reg( .D(DFF_162_N3), .CLK(CLK), .Q_N(n1911) );
	dfxbp_1 DFF_161_Q_reg( .D(DFF_161_N3), .CLK(CLK), .Q_N(n1120) );
	dfxbp_1 DFF_160_Q_reg( .D(DFF_160_N3), .CLK(CLK), .Q_N(n1908) );
	dfxbp_1 DFF_159_Q_reg( .D(DFF_159_N3), .CLK(CLK), .Q_N(n1121) );
	dfxbp_1 DFF_158_Q_reg( .D(DFF_158_N3), .CLK(CLK), .Q(n1122), .Q_N(n652) );
	dfxbp_1 DFF_157_Q_reg( .D(DFF_157_N3), .CLK(CLK), .Q(n660), .Q_N(n1170) );
	dfxbp_1 DFF_156_Q_reg( .D(DFF_156_N3), .CLK(CLK), .Q_N(n1169) );
	dfxbp_1 DFF_155_Q_reg( .D(DFF_155_N3), .CLK(CLK), .Q_N(n1893) );
	dfxbp_1 DFF_154_Q_reg( .D(DFF_154_N3), .CLK(CLK), .Q_N(n1228) );
	dfxbp_1 DFF_151_Q_reg( .D(DFF_151_N3), .CLK(CLK), .Q_N(n1888) );
	dfxbp_1 DFF_150_Q_reg( .D(DFF_150_N3), .CLK(CLK), .Q(n634) );
	dfxbp_1 DFF_149_Q_reg( .D(DFF_149_N3), .CLK(CLK), .Q(n614) );
	dfxbp_1 DFF_147_Q_reg( .D(DFF_147_N3), .CLK(CLK), .Q(n187) );
	dfxbp_1 DFF_145_Q_reg( .D(DFF_145_N3), .CLK(CLK), .Q_N(n1222) );
	dfxbp_1 DFF_143_Q_reg( .D(DFF_143_N3), .CLK(CLK), .Q(n189) );
	dfxbp_1 DFF_142_Q_reg( .D(DFF_142_N3), .CLK(CLK), .Q(n650), .Q_N(n1117) );
	dfxbp_1 DFF_141_Q_reg( .D(DFF_141_N3), .CLK(CLK), .Q(n617) );
	dfxbp_1 DFF_140_Q_reg( .D(DFF_140_N3), .CLK(CLK), .Q(n657) );
	dfxbp_1 DFF_139_Q_reg( .D(DFF_139_N3), .CLK(CLK), .Q_N(n1223) );
	dfxbp_1 DFF_137_Q_reg( .D(DFF_137_N3), .CLK(CLK), .Q(n1007), .Q_N(n3148gat) );
	dfxbp_1 DFF_136_Q_reg( .D(n33), .CLK(CLK), .Q(n1123) );
	dfxbp_1 DFF_135_Q_reg( .D(n9), .CLK(CLK), .Q(n626) );
	dfxbp_1 DFF_134_Q_reg( .D(DFF_134_N3), .CLK(CLK), .Q(n1115) );
	dfxbp_1 DFF_133_Q_reg( .D(DFF_133_N3), .CLK(CLK), .Q(n633) );
	dfxbp_1 DFF_132_Q_reg( .D(n6), .CLK(CLK), .Q(n621), .Q_N(n3106gat) );
	dfxbp_1 DFF_131_Q_reg( .D(DFF_131_N3), .CLK(CLK), .Q(n1124), .Q_N(n655) );
	dfxbp_1 DFF_130_Q_reg( .D(DFF_130_N3), .CLK(CLK), .Q_N(n1125) );
	dfxbp_1 DFF_128_Q_reg( .D(DFF_128_N3), .CLK(CLK), .Q(n1126) );
	dfxbp_1 DFF_125_Q_reg( .D(DFF_125_N3), .CLK(CLK), .Q(n665), .Q_N(n1151) );
	dfxbp_1 DFF_124_Q_reg( .D(DFF_124_N3), .CLK(CLK), .Q(n1150) );
	dfxbp_1 DFF_123_Q_reg( .D(DFF_123_N3), .CLK(CLK), .Q(n632), .Q_N(n1152) );
	dfxbp_1 DFF_121_Q_reg( .D(DFF_121_N3), .CLK(CLK), .Q(n1127) );
	dfxbp_1 DFF_119_Q_reg( .D(DFF_119_N3), .CLK(CLK), .Q(n200) );
	dfxbp_1 DFF_118_Q_reg( .D(DFF_118_N3), .CLK(CLK), .Q(n201) );
	dfxbp_1 DFF_117_Q_reg( .D(DFF_117_N3), .CLK(CLK), .Q(n644), .Q_N(n1204) );
	dfxbp_1 DFF_115_Q_reg( .D(DFF_115_N3), .CLK(CLK), .Q(n1110) );
	dfxbp_1 DFF_114_Q_reg( .D(DFF_114_N3), .CLK(CLK), .Q(n620), .Q_N(n1202) );
	dfxbp_1 DFF_113_Q_reg( .D(DFF_113_N3), .CLK(CLK), .Q(n639), .Q_N(n1207) );
	dfxbp_1 DFF_112_Q_reg( .D(DFF_112_N3), .CLK(CLK), .Q(n615), .Q_N(n1208) );
	dfxbp_1 DFF_111_Q_reg( .D(DFF_111_N3), .CLK(CLK), .Q_N(n1205) );
	dfxbp_1 DFF_110_Q_reg( .D(DFF_110_N3), .CLK(CLK), .Q(n638), .Q_N(n1200) );
	dfxbp_1 DFF_109_Q_reg( .D(DFF_109_N3), .CLK(CLK), .Q_N(n1128) );
	dfxbp_1 DFF_108_Q_reg( .D(DFF_108_N3), .CLK(CLK), .Q_N(n1221) );
	dfxbp_1 DFF_107_Q_reg( .D(DFF_107_N3), .CLK(CLK), .Q(n645), .Q_N(n1129) );
	dfxbp_1 DFF_106_Q_reg( .D(DFF_106_N3), .CLK(CLK), .Q(n637), .Q_N(n1220) );
	dfxbp_1 DFF_105_Q_reg( .D(DFF_105_N3), .CLK(CLK), .Q_N(n1130) );
	dfxbp_1 DFF_103_Q_reg( .D(n32), .CLK(CLK), .Q(n205) );
	dfxbp_1 DFF_102_Q_reg( .D(n31), .CLK(CLK), .Q(n206) );
	dfxbp_1 DFF_101_Q_reg( .D(DFF_101_N3), .CLK(CLK), .Q_N(n1224) );
	dfxbp_1 DFF_100_Q_reg( .D(DFF_100_N3), .CLK(CLK), .Q_N(n1217) );
	dfxbp_1 DFF_99_Q_reg( .D(DFF_99_N3), .CLK(CLK), .Q_N(n1225) );
	dfxbp_1 DFF_98_Q_reg( .D(DFF_98_N3), .CLK(CLK), .Q_N(n3126gat) );
	dfxbp_1 DFF_97_Q_reg( .D(DFF_97_N3), .CLK(CLK), .Q_N(n3127gat) );
	dfxbp_1 DFF_96_Q_reg( .D(DFF_96_N3), .CLK(CLK), .Q_N(n3128gat) );
	dfxbp_1 DFF_95_Q_reg( .D(DFF_95_N3), .CLK(CLK), .Q_N(n1198) );
	dfxbp_1 DFF_93_Q_reg( .D(DFF_93_N3), .CLK(CLK), .Q_N(n1197) );
	dfxbp_1 DFF_91_Q_reg( .D(DFF_91_N3), .CLK(CLK), .Q_N(n1900) );
	dfxbp_1 DFF_90_Q_reg( .D(DFF_90_N3), .CLK(CLK), .Q_N(n623) );
	dfxbp_1 DFF_89_Q_reg( .D(DFF_89_N3), .CLK(CLK), .Q_N(n1157) );
	dfxbp_1 DFF_88_Q_reg( .D(DFF_88_N3), .CLK(CLK), .Q(n1131), .Q_N(n659) );
	dfxbp_1 DFF_87_Q_reg( .D(DFF_87_N3), .CLK(CLK), .Q_N(n1154) );
	dfxbp_1 DFF_86_Q_reg( .D(DFF_86_N3), .CLK(CLK), .Q_N(n1155) );
	dfxbp_1 DFF_85_Q_reg( .D(DFF_85_N3), .CLK(CLK), .Q_N(n1158) );
	dfxbp_1 DFF_84_Q_reg( .D(DFF_84_N3), .CLK(CLK), .Q_N(n1159) );
	dfxbp_1 DFF_83_Q_reg( .D(DFF_83_N3), .CLK(CLK), .Q_N(n1156) );
	dfxbp_1 DFF_82_Q_reg( .D(DFF_82_N3), .CLK(CLK), .Q(n1153) );
	dfxbp_1 DFF_81_Q_reg( .D(DFF_81_N3), .CLK(CLK), .Q_N(n1901) );
	dfxbp_1 DFF_80_Q_reg( .D(DFF_80_N3), .CLK(CLK), .Q(n1160) );
	dfxbp_1 DFF_79_Q_reg( .D(DFF_79_N3), .CLK(CLK), .Q_N(n1132) );
	dfxbp_1 DFF_78_Q_reg( .D(DFF_78_N3), .CLK(CLK), .Q(n1161), .Q_N(n636) );
	dfxbp_1 DFF_77_Q_reg( .D(DFF_77_N3), .CLK(CLK), .Q_N(n1165) );
	dfxbp_1 DFF_76_Q_reg( .D(DFF_76_N3), .CLK(CLK), .Q_N(n1133) );
	dfxbp_1 DFF_75_Q_reg( .D(DFF_75_N3), .CLK(CLK), .Q(n1162), .Q_N(n663) );
	dfxbp_1 DFF_74_Q_reg( .D(DFF_74_N3), .CLK(CLK), .Q(n1149), .Q_N(n666) );
	dfxbp_1 DFF_73_Q_reg( .D(DFF_73_N3), .CLK(CLK), .Q(n648), .Q_N(n1164) );
	dfxbp_1 DFF_72_Q_reg( .D(DFF_72_N3), .CLK(CLK), .Q(n672), .Q_N(n1163) );
	dfxbp_1 DFF_71_Q_reg( .D(DFF_71_N3), .CLK(CLK), .Q_N(n1134) );
	dfxbp_1 DFF_70_Q_reg( .D(DFF_70_N3), .CLK(CLK), .Q(n226) );
	dfxbp_1 DFF_69_Q_reg( .D(DFF_69_N3), .CLK(CLK), .Q(n649) );
	dfxbp_1 DFF_67_Q_reg( .D(DFF_67_N3), .CLK(CLK), .Q_N(n1218) );
	dfxbp_1 DFF_66_Q_reg( .D(DFF_66_N3), .CLK(CLK), .Q_N(n1214) );
	dfxbp_1 DFF_65_Q_reg( .D(DFF_65_N3), .CLK(CLK), .Q_N(n1219) );
	dfxbp_1 DFF_64_Q_reg( .D(DFF_64_N3), .CLK(CLK), .Q_N(n1216) );
	dfxbp_1 DFF_63_Q_reg( .D(DFF_63_N3), .CLK(CLK), .Q(n643), .Q_N(n1215) );
	dfxbp_1 DFF_62_Q_reg( .D(DFF_62_N3), .CLK(CLK), .Q(n618), .Q_N(n1210) );
	dfxbp_1 DFF_61_Q_reg( .D(n606), .CLK(CLK), .Q(n641), .Q_N(n1211) );
	dfxbp_1 DFF_60_Q_reg( .D(DFF_60_N3), .CLK(CLK), .Q(n646), .Q_N(n1209) );
	dfxbp_1 DFF_59_Q_reg( .D(DFF_59_N3), .CLK(CLK), .Q(n642), .Q_N(n1212) );
	dfxbp_1 DFF_58_Q_reg( .D(DFF_58_N3), .CLK(CLK), .Q(n619), .Q_N(n1213) );
	dfxbp_1 DFF_57_Q_reg( .D(DFF_57_N3), .CLK(CLK), .Q_N(n1898) );
	dfxbp_1 DFF_56_Q_reg( .D(DFF_56_N3), .CLK(CLK), .Q_N(n1186) );
	dfxbp_1 DFF_55_Q_reg( .D(DFF_55_N3), .CLK(CLK), .Q(n628), .Q_N(n1187) );
	dfxbp_1 DFF_54_Q_reg( .D(DFF_54_N3), .CLK(CLK), .Q(n669), .Q_N(n1135) );
	dfxbp_1 DFF_53_Q_reg( .D(DFF_53_N3), .CLK(CLK), .Q(n629), .Q_N(n1193) );
	dfxbp_1 DFF_52_Q_reg( .D(DFF_52_N3), .CLK(CLK), .Q(n1188) );
	dfxbp_1 DFF_51_Q_reg( .D(DFF_51_N3), .CLK(CLK), .Q_N(n1194) );
	dfxbp_1 DFF_50_Q_reg( .D(DFF_50_N3), .CLK(CLK), .Q(n673), .Q_N(n1166) );
	dfxbp_1 DFF_49_Q_reg( .D(DFF_49_N3), .CLK(CLK), .Q_N(n640) );
	dfxbp_1 DFF_48_Q_reg( .D(DFF_48_N3), .CLK(CLK), .Q_N(n1136) );
	dfxbp_1 DFF_47_Q_reg( .D(DFF_47_N3), .CLK(CLK), .Q_N(n1899) );
	dfxbp_1 DFF_46_Q_reg( .D(DFF_46_N3), .CLK(CLK), .Q(n654), .Q_N(n1196) );
	dfxbp_1 DFF_45_Q_reg( .D(DFF_45_N3), .CLK(CLK), .Q(n1184), .Q_N(n667) );
	dfxbp_1 DFF_44_Q_reg( .D(DFF_44_N3), .CLK(CLK), .Q(n622), .Q_N(n1185) );
	dfxbp_1 DFF_43_Q_reg( .D(DFF_43_N3), .CLK(CLK), .Q_N(n1195) );
	dfxbp_1 DFF_42_Q_reg( .D(DFF_42_N3), .CLK(CLK), .Q_N(n1183) );
	dfxbp_1 DFF_41_Q_reg( .D(n17), .CLK(CLK), .Q(n1167), .Q_N(n675) );
	dfxbp_1 DFF_40_Q_reg( .D(n19), .CLK(CLK), .Q_N(n1137) );
	dfxbp_1 DFF_39_Q_reg( .D(n13), .CLK(CLK), .Q_N(n1138) );
	dfxbp_1 DFF_38_Q_reg( .D(n15), .CLK(CLK), .Q(n1168), .Q_N(n676) );
	dfxbp_1 DFF_37_Q_reg( .D(DFF_37_N3), .CLK(CLK), .Q_N(n1896) );
	dfxbp_1 DFF_36_Q_reg( .D(DFF_36_N3), .CLK(CLK), .Q_N(n1172) );
	dfxbp_1 DFF_35_Q_reg( .D(DFF_35_N3), .CLK(CLK), .Q(n653), .Q_N(n1139) );
	dfxbp_1 DFF_34_Q_reg( .D(DFF_34_N3), .CLK(CLK), .Q(n630), .Q_N(n1173) );
	dfxbp_1 DFF_33_Q_reg( .D(DFF_33_N3), .CLK(CLK), .Q(n670), .Q_N(n1140) );
	dfxbp_1 DFF_32_Q_reg( .D(DFF_32_N3), .CLK(CLK), .Q_N(n1174) );
	dfxbp_1 DFF_31_Q_reg( .D(DFF_31_N3), .CLK(CLK), .Q(n668), .Q_N(n1175) );
	dfxbp_1 DFF_30_Q_reg( .D(DFF_30_N3), .CLK(CLK), .Q(n631), .Q_N(n1141) );
	dfxbp_1 DFF_29_Q_reg( .D(DFF_29_N3), .CLK(CLK), .Q(n647), .Q_N(n1171) );
	dfxbp_1 DFF_28_Q_reg( .D(DFF_28_N3), .CLK(CLK), .Q_N(n1176) );
	dfxbp_1 DFF_27_Q_reg( .D(DFF_27_N3), .CLK(CLK), .Q_N(n1897) );
	dfxbp_1 DFF_26_Q_reg( .D(n25), .CLK(CLK), .Q(n1179), .Q_N(n664) );
	dfxbp_1 DFF_25_Q_reg( .D(n26), .CLK(CLK), .Q_N(n1142) );
	dfxbp_1 DFF_24_Q_reg( .D(n27), .CLK(CLK), .Q(n671), .Q_N(n1143) );
	dfxbp_1 DFF_23_Q_reg( .D(n28), .CLK(CLK), .Q_N(n1177) );
	dfxbp_1 DFF_22_Q_reg( .D(n29), .CLK(CLK), .Q_N(n1144) );
	dfxbp_1 DFF_21_Q_reg( .D(DFF_21_N3), .CLK(CLK), .Q_N(n246) );
	dfxbp_1 DFF_19_Q_reg( .D(DFF_19_N3), .CLK(CLK), .Q(n635), .Q_N(n1116) );
	dfxbp_1 DFF_18_Q_reg( .D(DFF_19_N3), .CLK(CLK), .Q(n658) );
	dfxbp_1 DFF_17_Q_reg( .D(DFF_17_N3), .CLK(CLK), .Q_N(n1876) );
	dfxbp_1 DFF_16_Q_reg( .D(DFF_16_N3), .CLK(CLK), .Q(n1180) );
	dfxbp_1 DFF_15_Q_reg( .D(DFF_15_N3), .CLK(CLK), .Q_N(n1902) );
	dfxbp_1 DFF_14_Q_reg( .D(n25), .CLK(CLK), .Q(n1192) );
	dfxbp_1 DFF_13_Q_reg( .D(n26), .CLK(CLK), .Q_N(n1189) );
	dfxbp_1 DFF_12_Q_reg( .D(n27), .CLK(CLK), .Q(n616) );
	dfxbp_1 DFF_11_Q_reg( .D(n28), .CLK(CLK), .Q(n1191) );
	dfxbp_1 DFF_10_Q_reg( .D(n29), .CLK(CLK), .Q_N(n1190) );
	dfxbp_1 DFF_9_Q_reg( .D(DFF_9_N3), .CLK(CLK), .Q(n251) );
	dfxbp_1 DFF_8_Q_reg( .D(n19), .CLK(CLK), .Q(n625), .Q_N(n1145) );
	dfxbp_1 DFF_7_Q_reg( .D(n17), .CLK(CLK), .Q(n627), .Q_N(n1206) );
	dfxbp_1 DFF_6_Q_reg( .D(n15), .CLK(CLK), .Q(n624), .Q_N(n1181) );
	dfxbp_1 DFF_5_Q_reg( .D(n13), .CLK(CLK), .Q_N(n1182) );
	dfxbp_1 DFF_4_Q_reg( .D(n19), .CLK(CLK), .Q(n661), .Q_N(n1178) );
	dfxbp_1 DFF_3_Q_reg( .D(n17), .CLK(CLK), .Q_N(n1203) );
	dfxbp_1 DFF_2_Q_reg( .D(n15), .CLK(CLK), .Q(n662), .Q_N(n1201) );
	dfxbp_1 DFF_1_Q_reg( .D(n13), .CLK(CLK), .Q(n651), .Q_N(n1199) );
	dfxbp_1 DFF_169_Q_reg( .D(DFF_169_N3), .CLK(CLK), .Q(n1112) );
	dfxbp_1 DFF_168_Q_reg( .D(DFF_168_N3), .CLK(CLK), .Q(n1771gat) );
	dfxbp_1 DFF_153_Q_reg( .D(DFF_153_N3), .CLK(CLK), .Q_N(n256) );
	dfxbp_1 DFF_138_Q_reg( .D(DFF_138_N3), .CLK(CLK), .Q(n2446gat) );
	dfxbp_1 DFF_92_Q_reg( .D(DFF_92_N3), .CLK(CLK), .Q(n1226) );
	dfxbp_1 DFF_126_Q_reg( .D(DFF_126_N3), .CLK(CLK), .Q_N(n258) );
	dfxbp_1 DFF_116_Q_reg( .D(DFF_116_N3), .CLK(CLK), .Q(n2021gat) );
	dfxbp_1 DFF_104_Q_reg( .D(DFF_104_N3), .CLK(CLK), .Q(n2084gat) );
	dfxbp_1 DFF_94_Q_reg( .D(DFF_94_N3), .CLK(CLK), .Q(n1227) );
	dfxbp_1 DFF_68_Q_reg( .D(n607), .CLK(CLK), .Q(n2102gat) );
	dfxbp_1 DFF_175_Q_reg( .D(DFF_175_N3), .CLK(CLK), .Q_N(n260) );
	dfxbp_1 DFF_166_Q_reg( .D(DFF_166_N3), .CLK(CLK), .Q(n2458gat) );
	dfxbp_1 DFF_152_Q_reg( .D(n10), .CLK(CLK), .Q(n2121gat) );
	dfxbp_1 DFF_146_Q_reg( .D(DFF_146_N3), .CLK(CLK), .Q(n2025gat) );
	dfxbp_1 DFF_144_Q_reg( .D(DFF_144_N3), .CLK(CLK), .Q(n2044gat) );
	dfxbp_1 DFF_129_Q_reg( .D(DFF_129_N3), .CLK(CLK), .Q(n1363gat) );
	dfxbp_1 DFF_127_Q_reg( .D(DFF_127_N3), .CLK(CLK), .Q(n1433gat) );
	dfxbp_1 DFF_122_Q_reg( .D(DFF_122_N3), .CLK(CLK), .Q(n2179gat) );
	dfxbp_1 DFF_120_Q_reg( .D(DFF_120_N3), .CLK(CLK), .Q(n1332gat) );
	dfxbp_1 DFF_20_Q_reg( .D(DFF_20_N3), .CLK(CLK), .Q(n2029gat) );
	dfxbp_1 DFF_165_Q_reg( .D(DFF_165_N3), .CLK(CLK), .Q_N(n261) );
	dfxbp_1 DFF_164_Q_reg( .D(DFF_164_N3), .CLK(CLK), .Q_N(n262) );
	dfxbp_1 DFF_148_Q_reg( .D(DFF_148_N3), .CLK(CLK), .Q(n2266gat) );
	inv_2 U711( .A(1'b0), .Y(n3152gat) );
	inv_2 U713( .A(1'b0), .Y(n3115gat) );
	inv_2 U715( .A(1'b0), .Y(n3112gat) );
	buf_1 U717( .A(n3142gat), .X(n3141gat) );
	buf_1 U718( .A(n3140gat), .X(n3139gat) );
	inv_1 U719( .A(n679), .Y(n9) );
	inv_1 U720( .A(n680), .Y(n607) );
	a211oi_1 U721( .A1(n1124), .A2(n1125), .B1(n681), .C1(n682), .Y(n6) );
	inv_1 U722( .A(DFF_146_N3), .Y(n681) );
	o211ai_1 U723( .A1(n3085gat), .A2(n683), .B1(n684), .C1(n685), .Y(n3151gat) );
	o22ai_1 U724( .A1(n650), .A2(n616), .B1(n686), .B2(n687), .Y(n3150gat) );
	nor4_1 U725( .A(n688), .B(n689), .C(n1222), .D(n1223), .Y(n3146gat) );
	nor2_1 U726( .A(n3106gat), .B(n690), .Y(n689) );
	nand4_1 U727( .A(n657), .B(n614), .C(n634), .D(n617), .Y(n688) );
	and2_0 U728( .A(n690), .B(n691), .X(n3145gat) );
	nand2_1 U729( .A(n692), .B(n178), .Y(n690) );
	or3_1 U730( .A(n693), .B(n694), .C(n695), .X(n3144gat) );
	or3_1 U731( .A(n695), .B(n694), .C(n696), .X(n3143gat) );
	o32ai_1 U732( .A1(n697), .A2(n698), .A3(n644), .B1(n699), .B2(n700), .Y( n694) );
	nand2_1 U733( .A(n1210), .B(n701), .Y(n700) );
	mux2i_1 U734( .A0(n702), .A1(n703), .S(n1209), .Y(n699) );
	nor2_1 U735( .A(n704), .B(n705), .Y(n703) );
	xor2_1 U736( .A(n1206), .B(n706), .X(n705) );
	o221ai_1 U737( .A1(n707), .A2(n708), .B1(n619), .B2(n709), .C1(n710), .Y( n702) );
	a22oi_1 U738( .A1(n1156), .A2(n711), .B1(n1158), .B2(n712), .Y(n710) );
	inv_1 U739( .A(n713), .Y(n712) );
	inv_1 U740( .A(n714), .Y(n709) );
	mux4_2 U741( .A0(n1155), .A1(n1154), .A2(n623), .A3(n1157), .S0(n1211), .S1(n642), .X(n714) );
	mux2i_1 U742( .A0(n1159), .A1(n659), .S(n1211), .Y(n708) );
	mux2_1 U743( .A0(n626), .A1(n1115), .S(n715), .X(n697) );
	o32ai_1 U744( .A1(n656), .A2(n3106gat), .A3(n633), .B1(n716), .B2(n717), .Y(n695) );
	nand2_1 U745( .A(n1110), .B(n618), .Y(n717) );
	mux2i_1 U746( .A0(n718), .A1(n719), .S(n1209), .Y(n716) );
	o221ai_1 U747( .A1(n704), .A2(n720), .B1(n1212), .B2(n721), .C1(n722), .Y( n719) );
	o21ai_0 U748( .A1(n723), .A2(n724), .B1(n725), .Y(n722) );
	o22ai_1 U749( .A1(n726), .A2(n622), .B1(n727), .B2(n671), .Y(n724) );
	inv_1 U750( .A(n728), .Y(n723) );
	a22oi_1 U751( .A1(n729), .A2(n1144), .B1(n730), .B2(n1183), .Y(n728) );
	mux2i_1 U752( .A0(n731), .A1(n732), .S(n1213), .Y(n721) );
	o221ai_1 U753( .A1(n1179), .A2(n727), .B1(n726), .B2(n654), .C1(n733), .Y( n732) );
	a22oi_1 U754( .A1(n1195), .A2(n730), .B1(n1177), .B2(n729), .Y(n733) );
	o22ai_1 U755( .A1(n726), .A2(n629), .B1(n727), .B2(n670), .Y(n731) );
	mux2i_1 U756( .A0(n1175), .A1(n1194), .S(n698), .Y(n720) );
	o221ai_1 U757( .A1(n713), .A2(n734), .B1(n704), .B2(n2084gat), .C1(n735), .Y(n718) );
	a221oi_1 U758( .A1(n725), .A2(n736), .B1(n737), .B2(n1213), .C1(n738), .Y( n735) );
	a21oi_1 U759( .A1(n704), .A2(n713), .B1(n739), .Y(n738) );
	mux2i_1 U760( .A0(n740), .A1(n741), .S(n1212), .Y(n737) );
	a221oi_1 U761( .A1(n1186), .A2(n730), .B1(n1172), .B2(n729), .C1(n742), .Y( n741) );
	o22ai_1 U762( .A1(n726), .A2(n628), .B1(n727), .B2(n653), .Y(n742) );
	a221oi_1 U763( .A1(n730), .A2(n640), .B1(n1171), .B2(n729), .C1(n743), .Y( n740) );
	o22ai_1 U764( .A1(n726), .A2(n669), .B1(n727), .B2(n630), .Y(n743) );
	o221ai_1 U765( .A1(n727), .A2(n631), .B1(n726), .B2(n673), .C1(n744), .Y( n736) );
	a22oi_1 U766( .A1(n1136), .A2(n730), .B1(n1176), .B2(n729), .Y(n744) );
	nor2_1 U767( .A(n1211), .B(n698), .Y(n729) );
	nor2_1 U768( .A(n3149gat), .B(n1211), .Y(n730) );
	nand2_1 U769( .A(n1211), .B(n698), .Y(n726) );
	nand2_1 U770( .A(n1211), .B(n3149gat), .Y(n727) );
	inv_1 U771( .A(n707), .Y(n725) );
	inv_1 U772( .A(n711), .Y(n704) );
	mux2_1 U773( .A0(n745), .A1(n746), .S(n747), .X(n3142gat) );
	o32ai_1 U774( .A1(n177), .A2(n748), .A3(n644), .B1(n1111), .B2(n749), .Y( n746) );
	a211oi_1 U775( .A1(n1112), .A2(n750), .B1(n3149gat), .C1(n701), .Y(n749) );
	inv_1 U776( .A(n734), .Y(n701) );
	o22ai_1 U777( .A1(n1113), .A2(n1148), .B1(n1114), .B2(n751), .Y(n745) );
	a21oi_1 U778( .A1(n1148), .A2(n752), .B1(n3149gat), .Y(n751) );
	nand2_1 U779( .A(n753), .B(n754), .Y(n3140gat) );
	nand3_1 U780( .A(n621), .B(n655), .C(n755), .Y(n754) );
	a21oi_1 U781( .A1(n635), .A2(n756), .B1(n3098gat), .Y(n755) );
	nand3_1 U782( .A(n757), .B(n758), .C(n3097gat), .Y(n756) );
	mux2i_1 U783( .A0(n759), .A1(n760), .S(n747), .Y(n753) );
	nand2_1 U784( .A(n761), .B(n762), .Y(n760) );
	nand3_1 U785( .A(n750), .B(n260), .C(n1204), .Y(n762) );
	mux2i_1 U786( .A0(n763), .A1(n1892), .S(n1147), .Y(n761) );
	a21oi_1 U787( .A1(n1204), .A2(n734), .B1(n626), .Y(n763) );
	o22ai_1 U788( .A1(n626), .A2(n674), .B1(n1115), .B2(n764), .Y(n759) );
	a21oi_1 U789( .A1(n765), .A2(n1148), .B1(n766), .Y(n764) );
	nor3_1 U790( .A(n698), .B(n1118), .C(n1204), .Y(n766) );
	nor2_1 U791( .A(n691), .B(n767), .Y(n765) );
	nor4_1 U792( .A(n1211), .B(n707), .C(n646), .D(n618), .Y(n767) );
	nor4_1 U793( .A(n768), .B(n769), .C(n713), .D(n618), .Y(n3138gat) );
	or4_1 U794( .A(n646), .B(n770), .C(n1219), .D(n1214), .X(n768) );
	o22ai_1 U795( .A1(n771), .A2(n772), .B1(n773), .B2(n774), .Y(n3137gat) );
	a222oi_1 U796( .A1(n775), .A2(n675), .B1(n776), .B2(n1203), .C1(n1133), .C2(n777), .Y(n774) );
	o22ai_1 U797( .A1(n778), .A2(n772), .B1(n773), .B2(n779), .Y(n3136gat) );
	a222oi_1 U798( .A1(n1137), .A2(n775), .B1(n776), .B2(n1178), .C1(n777), .C2(n663), .Y(n779) );
	o22ai_1 U799( .A1(n780), .A2(n772), .B1(n773), .B2(n781), .Y(n3135gat) );
	a222oi_1 U800( .A1(n775), .A2(n676), .B1(n776), .B2(n1201), .C1(n777), .C2( n636), .Y(n781) );
	o22ai_1 U801( .A1(n782), .A2(n772), .B1(n773), .B2(n783), .Y(n3134gat) );
	a222oi_1 U802( .A1(n1138), .A2(n775), .B1(n1199), .B2(n776), .C1(n1132), .C2(n777), .Y(n783) );
	o22ai_1 U803( .A1(n784), .A2(n772), .B1(n773), .B2(n785), .Y(n3133gat) );
	a222oi_1 U804( .A1(n775), .A2(n1196), .B1(n776), .B2(n664), .C1(n1165), .C2(n777), .Y(n785) );
	o22ai_1 U805( .A1(n786), .A2(n772), .B1(n773), .B2(n787), .Y(n3132gat) );
	a222oi_1 U806( .A1(n775), .A2(n1195), .B1(n776), .B2(n1177), .C1(n1164), .C2(n777), .Y(n787) );
	o22ai_1 U807( .A1(n788), .A2(n772), .B1(n773), .B2(n789), .Y(n3131gat) );
	a222oi_1 U808( .A1(n775), .A2(n1185), .B1(n776), .B2(n1143), .C1(n777), .C2(n666), .Y(n789) );
	o22ai_1 U809( .A1(n790), .A2(n772), .B1(n773), .B2(n791), .Y(n3130gat) );
	a222oi_1 U810( .A1(n775), .A2(n1183), .B1(n776), .B2(n1144), .C1(n1163), .C2(n777), .Y(n791) );
	o22ai_1 U811( .A1(n792), .A2(n772), .B1(n773), .B2(n793), .Y(n3129gat) );
	a222oi_1 U812( .A1(n775), .A2(n667), .B1(n1142), .B2(n776), .C1(n777), .C2( n3116gat), .Y(n793) );
	a21oi_1 U813( .A1(n3088gat), .A2(n794), .B1(n795), .Y(n773) );
	mux2i_1 U814( .A0(n794), .A1(n796), .S(n3088gat), .Y(n772) );
	nor3_1 U815( .A(n797), .B(n798), .C(n799), .Y(n796) );
	nor2_1 U816( .A(n800), .B(n801), .Y(n794) );
	o21ai_0 U817( .A1(n792), .A2(n802), .B1(n803), .Y(n3125gat) );
	inv_1 U818( .A(n804), .Y(n792) );
	o221ai_1 U819( .A1(n706), .A2(n805), .B1(n1188), .B2(n806), .C1(n807), .Y( n804) );
	a222oi_1 U820( .A1(n1174), .A2(n776), .B1(n808), .B2(n809), .C1(n1189), .C2(n810), .Y(n807) );
	o21ai_0 U821( .A1(n1146), .A2(n811), .B1(n812), .Y(n809) );
	inv_1 U822( .A(n775), .Y(n806) );
	o21ai_0 U823( .A1(n771), .A2(n802), .B1(n813), .Y(n3124gat) );
	xnor2_1 U824( .A(n1160), .B(n3116gat), .Y(n813) );
	a221oi_1 U825( .A1(n1154), .A2(n777), .B1(n1193), .B2(n775), .C1(n814), .Y( n771) );
	inv_1 U826( .A(n815), .Y(n814) );
	a21oi_1 U827( .A1(n776), .A2(n1140), .B1(n816), .Y(n815) );
	o32ai_1 U828( .A1(n817), .A2(n811), .A3(n656), .B1(n627), .B2(n818), .Y( n816) );
	o21ai_0 U829( .A1(n778), .A2(n802), .B1(n819), .Y(n3123gat) );
	xor2_1 U830( .A(n1153), .B(n706), .X(n819) );
	a221oi_1 U831( .A1(n1155), .A2(n777), .B1(n775), .B2(n1194), .C1(n820), .Y( n778) );
	o22ai_1 U832( .A1(n818), .A2(n625), .B1(n668), .B2(n821), .Y(n820) );
	o21ai_0 U833( .A1(n780), .A2(n802), .B1(n822), .Y(n3122gat) );
	a221oi_1 U834( .A1(n1157), .A2(n777), .B1(n1187), .B2(n775), .C1(n823), .Y( n780) );
	o22ai_1 U835( .A1(n818), .A2(n624), .B1(n821), .B2(n653), .Y(n823) );
	o21ai_0 U836( .A1(n782), .A2(n802), .B1(n824), .Y(n3121gat) );
	a221oi_1 U837( .A1(n623), .A2(n777), .B1(n1186), .B2(n775), .C1(n825), .Y( n782) );
	inv_1 U838( .A(n826), .Y(n825) );
	a22oi_1 U839( .A1(n810), .A2(n1182), .B1(n776), .B2(n1172), .Y(n826) );
	o21ai_0 U840( .A1(n784), .A2(n802), .B1(n827), .Y(n3120gat) );
	a221oi_1 U841( .A1(n659), .A2(n777), .B1(n1135), .B2(n775), .C1(n828), .Y( n784) );
	o22ai_1 U842( .A1(n818), .A2(n1192), .B1(n821), .B2(n630), .Y(n828) );
	o21ai_0 U843( .A1(n786), .A2(n802), .B1(n829), .Y(n3119gat) );
	a221oi_1 U844( .A1(n1159), .A2(n777), .B1(n640), .B2(n775), .C1(n830), .Y( n786) );
	o22ai_1 U845( .A1(n818), .A2(n1191), .B1(n821), .B2(n647), .Y(n830) );
	o21ai_0 U846( .A1(n788), .A2(n802), .B1(n831), .Y(n3118gat) );
	xnor2_1 U847( .A(n832), .B(n833), .Y(n831) );
	a221oi_1 U848( .A1(n1158), .A2(n777), .B1(n1166), .B2(n775), .C1(n834), .Y( n788) );
	o22ai_1 U849( .A1(n818), .A2(n616), .B1(n821), .B2(n631), .Y(n834) );
	inv_1 U850( .A(n776), .Y(n821) );
	o21ai_0 U851( .A1(n790), .A2(n802), .B1(n835), .Y(n3117gat) );
	xnor2_1 U852( .A(n836), .B(n837), .Y(n835) );
	inv_1 U853( .A(n795), .Y(n802) );
	a21oi_1 U854( .A1(n799), .A2(n797), .B1(n798), .Y(n795) );
	a221oi_1 U855( .A1(n1156), .A2(n777), .B1(n1136), .B2(n775), .C1(n838), .Y( n790) );
	inv_1 U856( .A(n839), .Y(n838) );
	a22oi_1 U857( .A1(n810), .A2(n1190), .B1(n776), .B2(n1176), .Y(n839) );
	nor2_1 U858( .A(n811), .B(n808), .Y(n776) );
	inv_1 U859( .A(n818), .Y(n810) );
	nand3_1 U860( .A(n812), .B(n817), .C(n811), .Y(n818) );
	nor2_1 U861( .A(n812), .B(n808), .Y(n775) );
	inv_1 U862( .A(n805), .Y(n777) );
	nand3_1 U863( .A(n811), .B(n812), .C(n808), .Y(n805) );
	inv_1 U864( .A(n817), .Y(n808) );
	o22ai_1 U865( .A1(n840), .A2(n841), .B1(n799), .B2(n842), .Y(n817) );
	o22ai_1 U866( .A1(n840), .A2(n799), .B1(n842), .B2(n797), .Y(n812) );
	a21oi_1 U867( .A1(n840), .A2(n843), .B1(n801), .Y(n811) );
	inv_1 U868( .A(n844), .Y(n801) );
	inv_1 U869( .A(n3095gat), .Y(n840) );
	nand2_1 U870( .A(n845), .B(n1162), .Y(n3114gat) );
	nand2_1 U871( .A(n1161), .B(n846), .Y(n3113gat) );
	or2_0 U872( .A(n847), .B(n1165), .X(n3111gat) );
	nand2_1 U873( .A(n848), .B(n648), .Y(n3110gat) );
	o21ai_0 U874( .A1(n849), .A2(n850), .B1(n1149), .Y(n3109gat) );
	nand2_1 U875( .A(n851), .B(n672), .Y(n3108gat) );
	nor2_1 U876( .A(n3106gat), .B(n692), .Y(n3107gat) );
	and2_0 U877( .A(n1124), .B(n1771gat), .X(n692) );
	o221ai_1 U878( .A1(n852), .A2(n853), .B1(n3087gat), .B2(n854), .C1(n855), .Y(n3105gat) );
	nand2_1 U879( .A(n856), .B(n841), .Y(n853) );
	o221ai_1 U880( .A1(n683), .A2(n857), .B1(n858), .B2(n684), .C1(n859), .Y( n3104gat) );
	nand3_1 U881( .A(n797), .B(n841), .C(n860), .Y(n684) );
	inv_1 U882( .A(n3094gat), .Y(n858) );
	nand2_1 U883( .A(n861), .B(n843), .Y(n857) );
	inv_1 U884( .A(n862), .Y(n30) );
	inv_1 U885( .A(n863), .Y(n29) );
	inv_1 U886( .A(n864), .Y(n28) );
	inv_1 U887( .A(n865), .Y(n27) );
	inv_1 U888( .A(n866), .Y(n25) );
	inv_1 U889( .A(n867), .Y(n15) );
	inv_1 U890( .A(n868), .Y(n10) );
	nor2_1 U891( .A(RST), .B(n869), .Y(DFF_9_N3) );
	xor2_1 U892( .A(n837), .B(n836), .X(n869) );
	xor2_1 U893( .A(n870), .B(n871), .X(n836) );
	a21oi_1 U894( .A1(n3084gat), .A2(n3083gat), .B1(n872), .Y(n871) );
	or2_0 U895( .A(n873), .B(n874), .X(n870) );
	mux2i_1 U896( .A0(n875), .A1(n876), .S(n3089gat), .Y(n837) );
	xor2_1 U897( .A(n3086gat), .B(n3085gat), .X(n876) );
	o21ai_0 U898( .A1(n797), .A2(n843), .B1(n844), .Y(n875) );
	nand2_1 U899( .A(n843), .B(n797), .Y(n844) );
	inv_1 U900( .A(n3086gat), .Y(n797) );
	and2_0 U901( .A(n33), .B(n803), .X(DFF_99_N3) );
	xor2_1 U902( .A(n877), .B(n878), .X(n803) );
	xor2_1 U903( .A(n1198), .B(n3128gat), .X(n878) );
	xnor2_1 U904( .A(n3127gat), .B(n3126gat), .Y(n877) );
	nor2_1 U905( .A(n879), .B(n846), .Y(DFF_98_N3) );
	xnor2_1 U906( .A(n880), .B(n1150), .Y(n846) );
	nand2_1 U907( .A(n1151), .B(n1152), .Y(n880) );
	nor2_1 U908( .A(n845), .B(n879), .Y(DFF_97_N3) );
	nor2_1 U909( .A(n1151), .B(n1152), .Y(n845) );
	a21oi_1 U910( .A1(n881), .A2(n882), .B1(RST), .Y(DFF_95_N3) );
	xor2_1 U911( .A(n2266gat), .B(n883), .X(n882) );
	nand2_1 U912( .A(n1151), .B(n632), .Y(n883) );
	nor2_1 U913( .A(RST), .B(n693), .Y(DFF_94_N3) );
	xor2_1 U914( .A(n884), .B(n885), .X(n693) );
	xnor2_1 U915( .A(n641), .B(n886), .Y(n885) );
	xor2_1 U916( .A(n1209), .B(n1210), .X(n886) );
	mux2i_1 U917( .A0(n887), .A1(n888), .S(n1197), .Y(n884) );
	o21ai_0 U918( .A1(n1212), .A2(n619), .B1(n707), .Y(n888) );
	o21ai_0 U919( .A1(n642), .A2(n619), .B1(n889), .Y(n887) );
	a21oi_1 U920( .A1(n890), .A2(n891), .B1(RST), .Y(DFF_93_N3) );
	xor2_1 U921( .A(n1893), .B(n892), .X(n891) );
	nor3_1 U922( .A(n615), .B(n849), .C(n893), .Y(n892) );
	inv_1 U923( .A(n894), .Y(n893) );
	nor2_1 U924( .A(n895), .B(n896), .Y(n890) );
	a21oi_1 U925( .A1(n897), .A2(n898), .B1(RST), .Y(DFF_92_N3) );
	nor4_1 U926( .A(n3090gat), .B(n1899), .C(n1896), .D(n1897), .Y(n898) );
	nor4_1 U927( .A(n1902), .B(n1900), .C(n1901), .D(n1898), .Y(n897) );
	nor2_1 U928( .A(RST), .B(n899), .Y(DFF_91_N3) );
	xnor2_1 U929( .A(n1153), .B(n706), .Y(n899) );
	xnor2_1 U930( .A(n900), .B(n901), .Y(n706) );
	xor2_1 U931( .A(n902), .B(n903), .X(n901) );
	xor2_1 U932( .A(n1154), .B(n1155), .X(n903) );
	xnor2_1 U933( .A(n623), .B(n1131), .Y(n902) );
	xor2_1 U934( .A(n904), .B(n905), .X(n900) );
	xor2_1 U935( .A(n1156), .B(n1157), .X(n905) );
	xnor2_1 U936( .A(n1159), .B(n1158), .Y(n904) );
	nand2_1 U937( .A(n906), .B(n907), .Y(DFF_90_N3) );
	inv_1 U938( .A(DFF_36_N3), .Y(n907) );
	nand2_1 U939( .A(n906), .B(n908), .Y(DFF_89_N3) );
	inv_1 U940( .A(DFF_35_N3), .Y(n908) );
	nand2_1 U941( .A(n906), .B(n909), .Y(DFF_88_N3) );
	inv_1 U942( .A(DFF_34_N3), .Y(n909) );
	nand2_1 U943( .A(n906), .B(n910), .Y(DFF_87_N3) );
	inv_1 U944( .A(DFF_33_N3), .Y(n910) );
	nand2_1 U945( .A(n906), .B(n911), .Y(DFF_86_N3) );
	inv_1 U946( .A(DFF_31_N3), .Y(n911) );
	nand2_1 U947( .A(n906), .B(n912), .Y(DFF_85_N3) );
	inv_1 U948( .A(DFF_30_N3), .Y(n912) );
	nand2_1 U949( .A(n906), .B(n913), .Y(DFF_84_N3) );
	inv_1 U950( .A(DFF_29_N3), .Y(n913) );
	nand2_1 U951( .A(n906), .B(n914), .Y(DFF_83_N3) );
	inv_1 U952( .A(DFF_28_N3), .Y(n914) );
	nand2_1 U953( .A(n906), .B(n915), .Y(DFF_82_N3) );
	inv_1 U954( .A(DFF_32_N3), .Y(n915) );
	nor2_1 U955( .A(RST), .B(n916), .Y(DFF_81_N3) );
	xor2_1 U956( .A(n1160), .B(n3116gat), .X(n916) );
	xnor2_1 U957( .A(n917), .B(n918), .Y(n3116gat) );
	xor2_1 U958( .A(n919), .B(n920), .X(n918) );
	xor2_1 U959( .A(n1149), .B(n1161), .X(n920) );
	xor2_1 U960( .A(n1132), .B(n1133), .X(n919) );
	xor2_1 U961( .A(n921), .B(n922), .X(n917) );
	xor2_1 U962( .A(n1162), .B(n1163), .X(n922) );
	xor2_1 U963( .A(n1165), .B(n648), .X(n921) );
	o21ai_0 U964( .A1(n923), .A2(n924), .B1(n906), .Y(DFF_80_N3) );
	o21ai_0 U965( .A1(n923), .A2(n925), .B1(n906), .Y(DFF_79_N3) );
	o21ai_0 U966( .A1(n923), .A2(n867), .B1(n906), .Y(DFF_78_N3) );
	o21ai_0 U967( .A1(n923), .A2(n866), .B1(n906), .Y(DFF_77_N3) );
	o21ai_0 U968( .A1(n923), .A2(n926), .B1(n906), .Y(DFF_76_N3) );
	o21ai_0 U969( .A1(n923), .A2(n927), .B1(n906), .Y(DFF_75_N3) );
	o21ai_0 U970( .A1(n923), .A2(n865), .B1(n906), .Y(DFF_74_N3) );
	o21ai_0 U971( .A1(n923), .A2(n864), .B1(n906), .Y(DFF_73_N3) );
	o21ai_0 U972( .A1(n923), .A2(n863), .B1(n906), .Y(DFF_72_N3) );
	nand4_1 U973( .A(DFF_119_N3), .B(n1219), .C(n928), .D(n929), .Y(n906) );
	a211oi_1 U974( .A1(n1209), .A2(n930), .B1(n618), .C1(n1214), .Y(n929) );
	o21ai_0 U975( .A1(n1211), .A2(n707), .B1(n713), .Y(n930) );
	nand2_1 U976( .A(n1211), .B(n931), .Y(n713) );
	nand2_1 U977( .A(n1212), .B(n619), .Y(n707) );
	mux2i_1 U978( .A0(n769), .A1(n932), .S(n1134), .Y(n928) );
	nand3_1 U979( .A(n1216), .B(n643), .C(n1218), .Y(n932) );
	inv_1 U980( .A(n933), .Y(n769) );
	inv_1 U981( .A(n934), .Y(n923) );
	o32ai_1 U982( .A1(n852), .A2(n3088gat), .A3(n856), .B1(n683), .B2(n935), .Y(n934) );
	nand4_1 U983( .A(n3086gat), .B(n936), .C(n874), .D(n621), .Y(n683) );
	nor2_1 U984( .A(n841), .B(n3087gat), .Y(n874) );
	inv_1 U985( .A(n800), .Y(n936) );
	nor2_1 U986( .A(n937), .B(n680), .Y(DFF_70_N3) );
	nand3_1 U987( .A(n1190), .B(n33), .C(n1117), .Y(n680) );
	nor3_1 U988( .A(n256), .B(n938), .C(n868), .Y(DFF_69_N3) );
	nand2_1 U989( .A(n33), .B(n1888), .Y(n868) );
	inv_1 U990( .A(n939), .Y(n938) );
	nor2_1 U991( .A(n855), .B(n940), .Y(DFF_67_N3) );
	xor2_1 U992( .A(n1130), .B(n941), .X(n855) );
	nor2_1 U993( .A(n859), .B(n940), .Y(DFF_66_N3) );
	a21oi_1 U994( .A1(n942), .A2(n1128), .B1(n943), .Y(n859) );
	nor3_1 U995( .A(n940), .B(n686), .C(n687), .Y(DFF_65_N3) );
	and2_0 U996( .A(n637), .B(n944), .X(n687) );
	nor2_1 U997( .A(n685), .B(n940), .Y(DFF_64_N3) );
	inv_1 U998( .A(n940), .Y(DFF_63_N3) );
	nand2_1 U999( .A(n945), .B(DFF_96_N3), .Y(n940) );
	inv_1 U1000( .A(n879), .Y(DFF_96_N3) );
	nor2_1 U1001( .A(n851), .B(n946), .Y(DFF_62_N3) );
	xor2_1 U1002( .A(n639), .B(n849), .X(n851) );
	nor3_1 U1003( .A(n946), .B(n849), .C(n850), .Y(DFF_60_N3) );
	a21oi_1 U1004( .A1(n1200), .A2(n947), .B1(n1202), .Y(n850) );
	nor3_1 U1005( .A(n638), .B(n620), .C(n948), .Y(n849) );
	nor2_1 U1006( .A(n949), .B(n946), .Y(DFF_59_N3) );
	nor2_1 U1007( .A(n848), .B(n946), .Y(DFF_58_N3) );
	inv_1 U1008( .A(n606), .Y(n946) );
	nor2_1 U1009( .A(n879), .B(n895), .Y(n606) );
	nand2_1 U1010( .A(n881), .B(n33), .Y(n879) );
	xor2_1 U1011( .A(n948), .B(n1200), .X(n848) );
	and2_0 U1012( .A(n33), .B(n824), .X(DFF_57_N3) );
	xor2_1 U1013( .A(n640), .B(n950), .X(n824) );
	xor2_1 U1014( .A(n951), .B(n952), .X(n950) );
	xor2_1 U1015( .A(n953), .B(n954), .X(n952) );
	xor2_1 U1016( .A(n1193), .B(n1194), .X(n954) );
	xor2_1 U1017( .A(n1187), .B(n1188), .X(n953) );
	xor2_1 U1018( .A(n955), .B(n956), .X(n951) );
	xor2_1 U1019( .A(n1166), .B(n1186), .X(n956) );
	xor2_1 U1020( .A(n1135), .B(n1136), .X(n955) );
	o221ai_1 U1021( .A1(n957), .A2(n958), .B1(n959), .B2(n960), .C1(n961), .Y( DFF_56_N3) );
	nand2_1 U1022( .A(n962), .B(n13), .Y(n961) );
	inv_1 U1023( .A(n925), .Y(n13) );
	xor2_1 U1024( .A(n1911), .B(n963), .X(n958) );
	o221ai_1 U1025( .A1(n964), .A2(n960), .B1(n867), .B2(n965), .C1(n966), .Y( DFF_55_N3) );
	nand3_1 U1026( .A(n967), .B(n963), .C(n968), .Y(n966) );
	nand3_1 U1027( .A(n969), .B(n652), .C(n1120), .Y(n963) );
	inv_1 U1028( .A(n970), .Y(n967) );
	a21oi_1 U1029( .A1(n652), .A2(n969), .B1(n1120), .Y(n970) );
	o22ai_1 U1030( .A1(n866), .A2(n965), .B1(n971), .B2(n960), .Y(DFF_54_N3) );
	o221ai_1 U1031( .A1(n972), .A2(n957), .B1(n973), .B2(n960), .C1(n974), .Y( DFF_53_N3) );
	nand2_1 U1032( .A(n962), .B(n17), .Y(n974) );
	inv_1 U1033( .A(n926), .Y(n17) );
	xnor2_1 U1034( .A(n1121), .B(n975), .Y(n972) );
	o221ai_1 U1035( .A1(n957), .A2(n976), .B1(n977), .B2(n960), .C1(n978), .Y( DFF_52_N3) );
	nand2_1 U1036( .A(n962), .B(n26), .Y(n978) );
	inv_1 U1037( .A(n924), .Y(n26) );
	xor2_1 U1038( .A(n1908), .B(n979), .X(n976) );
	nand2_1 U1039( .A(n975), .B(n980), .Y(n979) );
	o21ai_0 U1040( .A1(n1122), .A2(n1120), .B1(n1121), .Y(n980) );
	o221ai_1 U1041( .A1(n957), .A2(n981), .B1(n982), .B2(n960), .C1(n983), .Y( DFF_51_N3) );
	nand2_1 U1042( .A(n962), .B(n19), .Y(n983) );
	inv_1 U1043( .A(n927), .Y(n19) );
	xor2_1 U1044( .A(n1122), .B(n969), .X(n981) );
	and2_0 U1045( .A(n1121), .B(n975), .X(n969) );
	inv_1 U1046( .A(n968), .Y(n957) );
	nor3_1 U1047( .A(n984), .B(RST), .C(n962), .Y(n968) );
	inv_1 U1048( .A(n965), .Y(n962) );
	o22ai_1 U1049( .A1(n865), .A2(n965), .B1(n985), .B2(n960), .Y(DFF_50_N3) );
	o22ai_1 U1050( .A1(n864), .A2(n965), .B1(n986), .B2(n960), .Y(DFF_49_N3) );
	o22ai_1 U1051( .A1(n863), .A2(n965), .B1(n987), .B2(n960), .Y(DFF_48_N3) );
	nand2_1 U1052( .A(n984), .B(n33), .Y(n960) );
	nand2_1 U1053( .A(n873), .B(n988), .Y(n965) );
	and2_0 U1054( .A(n33), .B(n822), .X(DFF_47_N3) );
	xnor2_1 U1055( .A(n622), .B(n989), .Y(n822) );
	xor2_1 U1056( .A(n990), .B(n991), .X(n989) );
	xor2_1 U1057( .A(n992), .B(n993), .X(n991) );
	xor2_1 U1058( .A(n1195), .B(n1196), .X(n993) );
	xor2_1 U1059( .A(n1183), .B(n1184), .X(n992) );
	xor2_1 U1060( .A(n994), .B(n995), .X(n990) );
	xor2_1 U1061( .A(n1167), .B(n1168), .X(n995) );
	xor2_1 U1062( .A(n1137), .B(n1138), .X(n994) );
	o22ai_1 U1063( .A1(n996), .A2(n866), .B1(n997), .B2(n998), .Y(tempDFF_46_N3) );
	xnor2_1 U1064( .A(n999), .B(n1169), .Y(n997) );
	o22ai_1 U1065( .A1(n996), .A2(n924), .B1(n998), .B2(n1000), .Y(DFF_45_N3) );
	xor2_1 U1066( .A(n262), .B(n1001), .X(n1000) );
	nand2_1 U1067( .A(n999), .B(n1002), .Y(n1001) );
	o21ai_0 U1068( .A1(n1119), .A2(n660), .B1(n1169), .Y(n1002) );
	o22ai_1 U1069( .A1(n996), .A2(n865), .B1(n1003), .B2(n998), .Y(DFF_44_N3) );
	xnor2_1 U1070( .A(n1004), .B(n1119), .Y(n1003) );
	o22ai_1 U1071( .A1(n996), .A2(n864), .B1(n1005), .B2(n998), .Y(DFF_43_N3) );
	xor2_1 U1072( .A(n1006), .B(n1170), .X(n1005) );
	o22ai_1 U1073( .A1(n996), .A2(n863), .B1(n998), .B2(n1008), .Y(DFF_42_N3) );
	xor2_1 U1074( .A(n261), .B(n1009), .X(n1008) );
	nand2_1 U1075( .A(n1004), .B(n1119), .Y(n1009) );
	nor2_1 U1076( .A(n1006), .B(n660), .Y(n1004) );
	nand2_1 U1077( .A(n999), .B(n1169), .Y(n1006) );
	nand2_1 U1078( .A(n996), .B(n33), .Y(n998) );
	a21oi_1 U1079( .A1(n3087gat), .A2(n1010), .B1(n984), .Y(n996) );
	nor3_1 U1080( .A(n841), .B(n860), .C(n852), .Y(n984) );
	inv_1 U1081( .A(n856), .Y(n860) );
	inv_1 U1082( .A(n854), .Y(n1010) );
	nand2_1 U1083( .A(n988), .B(n3088gat), .Y(n854) );
	nor4_1 U1084( .A(n935), .B(n800), .C(n3086gat), .D(n3106gat), .Y(n988) );
	and2_0 U1085( .A(n33), .B(n829), .X(DFF_37_N3) );
	xor2_1 U1086( .A(n647), .B(n1011), .X(n829) );
	xor2_1 U1087( .A(n1012), .B(n1013), .X(n1011) );
	xor2_1 U1088( .A(n1014), .B(n1015), .X(n1013) );
	xor2_1 U1089( .A(n1175), .B(n1176), .X(n1015) );
	xor2_1 U1090( .A(n1173), .B(n1174), .X(n1014) );
	xor2_1 U1091( .A(n1016), .B(n1017), .X(n1012) );
	xor2_1 U1092( .A(n1141), .B(n1172), .X(n1017) );
	xor2_1 U1093( .A(n1139), .B(n1140), .X(n1016) );
	o22ai_1 U1094( .A1(n842), .A2(n925), .B1(n1018), .B2(n959), .Y(DFF_36_N3) );
	inv_1 U1095( .A(n3078gat), .Y(n959) );
	nand2_1 U1096( .A(n3069gat), .B(n33), .Y(n925) );
	o22ai_1 U1097( .A1(n842), .A2(n867), .B1(n1018), .B2(n964), .Y(DFF_35_N3) );
	inv_1 U1098( .A(n3079gat), .Y(n964) );
	nand2_1 U1099( .A(n3070gat), .B(n33), .Y(n867) );
	o22ai_1 U1100( .A1(n1018), .A2(n971), .B1(n842), .B2(n866), .Y(DFF_34_N3) );
	nand2_1 U1101( .A(n3068gat), .B(n33), .Y(n866) );
	inv_1 U1102( .A(n3077gat), .Y(n971) );
	o22ai_1 U1103( .A1(n842), .A2(n926), .B1(n1018), .B2(n973), .Y(DFF_33_N3) );
	inv_1 U1104( .A(n3081gat), .Y(n973) );
	nand2_1 U1105( .A(n3072gat), .B(n33), .Y(n926) );
	o22ai_1 U1106( .A1(n1018), .A2(n977), .B1(n842), .B2(n924), .Y(DFF_32_N3) );
	nand2_1 U1107( .A(n3073gat), .B(n33), .Y(n924) );
	inv_1 U1108( .A(n3082gat), .Y(n977) );
	o22ai_1 U1109( .A1(n842), .A2(n927), .B1(n1018), .B2(n982), .Y(DFF_31_N3) );
	inv_1 U1110( .A(n3080gat), .Y(n982) );
	nand2_1 U1111( .A(n3071gat), .B(n33), .Y(n927) );
	o22ai_1 U1112( .A1(n1018), .A2(n985), .B1(n842), .B2(n865), .Y(DFF_30_N3) );
	nand2_1 U1113( .A(n3066gat), .B(n33), .Y(n865) );
	inv_1 U1114( .A(n3075gat), .Y(n985) );
	o22ai_1 U1115( .A1(n1018), .A2(n986), .B1(n842), .B2(n864), .Y(DFF_29_N3) );
	nand2_1 U1116( .A(n3067gat), .B(n33), .Y(n864) );
	inv_1 U1117( .A(n3076gat), .Y(n986) );
	o22ai_1 U1118( .A1(n842), .A2(n863), .B1(n1018), .B2(n987), .Y(DFF_28_N3) );
	inv_1 U1119( .A(n3074gat), .Y(n987) );
	nand2_1 U1120( .A(n3095gat), .B(n33), .Y(n1018) );
	nand2_1 U1121( .A(n3065gat), .B(n33), .Y(n863) );
	inv_1 U1122( .A(n3093gat), .Y(n842) );
	and2_0 U1123( .A(n33), .B(n827), .X(DFF_27_N3) );
	xor2_1 U1124( .A(n1177), .B(n1019), .X(n827) );
	xor2_1 U1125( .A(n1020), .B(n1021), .X(n1019) );
	xor2_1 U1126( .A(n1022), .B(n1023), .X(n1021) );
	xor2_1 U1127( .A(n1201), .B(n1203), .X(n1023) );
	xor2_1 U1128( .A(n1179), .B(n1199), .X(n1022) );
	xor2_1 U1129( .A(n1024), .B(n1025), .X(n1020) );
	xor2_1 U1130( .A(n1144), .B(n1178), .X(n1025) );
	xor2_1 U1131( .A(n1142), .B(n1143), .X(n1024) );
	nor2_1 U1132( .A(RST), .B(n2029gat), .Y(DFF_21_N3) );
	a21oi_1 U1133( .A1(n635), .A2(n658), .B1(RST), .Y(DFF_20_N3) );
	nor3_1 U1134( .A(n1876), .B(n3099gat), .C(RST), .Y(DFF_19_N3) );
	nor2_1 U1135( .A(n1180), .B(RST), .Y(DFF_17_N3) );
	nor3_1 U1136( .A(n1026), .B(n1125), .C(n1027), .Y(DFF_178_N3) );
	nor3_1 U1137( .A(n1028), .B(n1029), .C(n941), .Y(DFF_177_N3) );
	nor2_1 U1138( .A(n1028), .B(n862), .Y(DFF_176_N3) );
	nand2_1 U1139( .A(n943), .B(n33), .Y(n862) );
	nand4_1 U1140( .A(n1200), .B(n1202), .C(n1030), .D(n1208), .Y(n1028) );
	nor2_1 U1141( .A(n1205), .B(n1207), .Y(n1030) );
	nor3_1 U1142( .A(n1026), .B(n1221), .C(n645), .Y(DFF_175_N3) );
	nor3_1 U1143( .A(n1031), .B(n1032), .C(n1033), .Y(DFF_174_N3) );
	nor4_1 U1144( .A(n1208), .B(n639), .C(n620), .D(n894), .Y(n1032) );
	nand2_1 U1145( .A(n1205), .B(n638), .Y(n894) );
	nor2_1 U1146( .A(n1034), .B(n679), .Y(DFF_173_N3) );
	nand3_1 U1147( .A(n1035), .B(n685), .C(n1220), .Y(n679) );
	nor2_1 U1148( .A(n1129), .B(n1221), .Y(n685) );
	nor3_1 U1149( .A(n1027), .B(n1029), .C(n637), .Y(DFF_171_N3) );
	nor3_1 U1150( .A(n941), .B(n1036), .C(n1029), .Y(DFF_170_N3) );
	inv_1 U1151( .A(n686), .Y(n941) );
	and3_1 U1152( .A(n1037), .B(n33), .C(n1038), .X(DFF_16_N3) );
	nor4_1 U1153( .A(n1039), .B(n1219), .C(n1209), .D(n1214), .Y(DFF_169_N3) );
	nand3_1 U1154( .A(n933), .B(n711), .C(DFF_113_N3), .Y(n1039) );
	nor2_1 U1155( .A(n889), .B(n1211), .Y(n711) );
	inv_1 U1156( .A(n931), .Y(n889) );
	nor2_1 U1157( .A(n1213), .B(n1212), .Y(n931) );
	nor3_1 U1158( .A(n1218), .B(n1216), .C(n643), .Y(n933) );
	nor2_1 U1159( .A(n937), .B(n1040), .Y(DFF_168_N3) );
	nor2_1 U1160( .A(RST), .B(n2458gat), .Y(DFF_167_N3) );
	nor2_1 U1161( .A(RST), .B(n633), .Y(DFF_166_N3) );
	and2_0 U1162( .A(n33), .B(n1183), .X(DFF_165_N3) );
	nor2_1 U1163( .A(n1184), .B(RST), .Y(DFF_164_N3) );
	nor2_1 U1164( .A(RST), .B(n622), .Y(DFF_163_N3) );
	and2_0 U1165( .A(n33), .B(n1186), .X(DFF_162_N3) );
	nor2_1 U1166( .A(RST), .B(n628), .Y(DFF_161_N3) );
	nor2_1 U1167( .A(n1188), .B(RST), .Y(DFF_160_N3) );
	nor2_1 U1168( .A(RST), .B(n1041), .Y(DFF_15_N3) );
	xor2_1 U1169( .A(n833), .B(n832), .X(n1041) );
	xor2_1 U1170( .A(n1191), .B(n1042), .X(n832) );
	xor2_1 U1171( .A(n1189), .B(n1190), .X(n1042) );
	xor2_1 U1172( .A(n1043), .B(n1044), .X(n833) );
	a21oi_1 U1173( .A1(n1045), .A2(n1038), .B1(n1046), .Y(n1044) );
	mux2i_1 U1174( .A0(n1047), .A1(n1048), .S(n1181), .Y(n1046) );
	xor2_1 U1175( .A(n1182), .B(n1045), .X(n1048) );
	nand2_1 U1176( .A(n1182), .B(n1049), .Y(n1047) );
	inv_1 U1177( .A(n1045), .Y(n1049) );
	xor2_1 U1178( .A(n616), .B(n1192), .X(n1045) );
	a21oi_1 U1179( .A1(n1145), .A2(n1206), .B1(n1037), .Y(n1043) );
	nor2_1 U1180( .A(RST), .B(n629), .Y(DFF_159_N3) );
	and2_0 U1181( .A(n33), .B(n1194), .X(DFF_158_N3) );
	and2_0 U1182( .A(n33), .B(n1195), .X(DFF_157_N3) );
	nor2_1 U1183( .A(RST), .B(n654), .Y(DFF_156_N3) );
	and2_0 U1184( .A(n33), .B(n1197), .X(DFF_155_N3) );
	and2_0 U1185( .A(n33), .B(n1217), .X(DFF_154_N3) );
	nor2_1 U1186( .A(RST), .B(n2121gat), .Y(DFF_153_N3) );
	nor2_1 U1187( .A(RST), .B(n634), .Y(DFF_151_N3) );
	nor2_1 U1188( .A(RST), .B(n614), .Y(DFF_150_N3) );
	and2_0 U1189( .A(n33), .B(n1222), .X(DFF_149_N3) );
	and2_0 U1190( .A(n33), .B(n1198), .X(DFF_148_N3) );
	nor2_1 U1191( .A(RST), .B(n2025gat), .Y(DFF_147_N3) );
	nor2_1 U1192( .A(n1033), .B(n757), .Y(DFF_146_N3) );
	inv_1 U1193( .A(n1050), .Y(n757) );
	nor2_1 U1194( .A(RST), .B(n2044gat), .Y(DFF_145_N3) );
	nor3_1 U1195( .A(n189), .B(n1126), .C(n1051), .Y(DFF_144_N3) );
	nor4_1 U1196( .A(n1125), .B(n682), .C(n1033), .D(n617), .Y(DFF_142_N3) );
	or2_0 U1197( .A(n1036), .B(RST), .X(n1033) );
	and4_1 U1198( .A(n1207), .B(n1052), .C(n1053), .D(n3149gat), .X(n1036) );
	nand2_1 U1199( .A(n1054), .B(n1055), .Y(n1052) );
	nand3_1 U1200( .A(n1202), .B(n638), .C(n949), .Y(n1055) );
	mux2i_1 U1201( .A0(n1056), .A1(n1057), .S(n1200), .Y(n1054) );
	nor3_1 U1202( .A(n1058), .B(n662), .C(n1059), .Y(n1057) );
	mux2i_1 U1203( .A0(n1060), .A1(n1061), .S(n1178), .Y(n1059) );
	inv_1 U1204( .A(n1062), .Y(n1061) );
	a21oi_1 U1205( .A1(n1063), .A2(n615), .B1(n1205), .Y(n1060) );
	o211ai_1 U1206( .A1(n1063), .A2(n615), .B1(n620), .C1(n651), .Y(n1058) );
	inv_1 U1207( .A(n1064), .Y(n1063) );
	nor3_1 U1208( .A(n1065), .B(n1201), .C(n1202), .Y(n1056) );
	o21ai_0 U1209( .A1(n1066), .A2(n661), .B1(n1067), .Y(n1065) );
	o32ai_1 U1210( .A1(n1064), .A2(n1205), .A3(n615), .B1(n1199), .B2(n1068), .Y(n1067) );
	a21oi_1 U1211( .A1(n949), .A2(n1064), .B1(n1178), .Y(n1068) );
	a21oi_1 U1212( .A1(n1208), .A2(n1064), .B1(n1062), .Y(n1066) );
	o21ai_0 U1213( .A1(n947), .A2(n1064), .B1(n1205), .Y(n1062) );
	inv_1 U1214( .A(n948), .Y(n947) );
	nand2_1 U1215( .A(n1208), .B(n1205), .Y(n948) );
	nand2_1 U1216( .A(n1203), .B(n651), .Y(n1064) );
	nor2_1 U1217( .A(RST), .B(n657), .Y(DFF_141_N3) );
	and2_0 U1218( .A(n33), .B(n1223), .X(DFF_140_N3) );
	a21oi_1 U1219( .A1(n1069), .A2(n1070), .B1(RST), .Y(DFF_139_N3) );
	nand4_1 U1220( .A(n873), .B(n1071), .C(n1072), .D(n3086gat), .Y(n1070) );
	nor2_1 U1221( .A(n3106gat), .B(n800), .Y(n1072) );
	nand2_1 U1222( .A(n3093gat), .B(n872), .Y(n800) );
	inv_1 U1223( .A(n935), .Y(n1071) );
	nand2_1 U1224( .A(n3085gat), .B(n861), .Y(n935) );
	or2_0 U1225( .A(n3091gat), .B(n3092gat), .X(n861) );
	nor2_1 U1226( .A(n799), .B(n3088gat), .Y(n873) );
	inv_1 U1227( .A(n3087gat), .Y(n799) );
	or3_1 U1228( .A(n841), .B(n856), .C(n852), .X(n1069) );
	nand4_1 U1229( .A(n3094gat), .B(n3086gat), .C(n1073), .D(n621), .Y(n852) );
	nand3_1 U1230( .A(n1073), .B(n621), .C(n3087gat), .Y(n856) );
	inv_1 U1231( .A(n798), .Y(n1073) );
	nand3_1 U1232( .A(n872), .B(n843), .C(n3095gat), .Y(n798) );
	inv_1 U1233( .A(n3085gat), .Y(n843) );
	nor2_1 U1234( .A(n3083gat), .B(n3084gat), .Y(n872) );
	inv_1 U1235( .A(n3088gat), .Y(n841) );
	nor2_1 U1236( .A(RST), .B(n1074), .Y(DFF_138_N3) );
	nor2_1 U1237( .A(n1123), .B(RST), .Y(DFF_137_N3) );
	nor4_1 U1238( .A(n1075), .B(n1027), .C(n1128), .D(n1220), .Y(DFF_134_N3) );
	nand2_1 U1239( .A(DFF_71_N3), .B(n1130), .Y(n1075) );
	nor2_1 U1240( .A(n747), .B(RST), .Y(DFF_71_N3) );
	inv_1 U1241( .A(n1051), .Y(DFF_133_N3) );
	nand2_1 U1242( .A(n33), .B(n655), .Y(n1051) );
	nor2_1 U1243( .A(n937), .B(n1076), .Y(DFF_131_N3) );
	o211ai_1 U1244( .A1(n1116), .A2(n758), .B1(n939), .C1(n1180), .Y(n937) );
	nand2_1 U1245( .A(n3147gat), .B(n1077), .Y(n939) );
	inv_1 U1246( .A(n3100gat), .Y(n1077) );
	nand2_1 U1247( .A(n2446gat), .B(n1007), .Y(n3147gat) );
	nand2_1 U1248( .A(n246), .B(n658), .Y(n758) );
	nor2_1 U1249( .A(RST), .B(n1363gat), .Y(DFF_130_N3) );
	nor2_1 U1250( .A(n1126), .B(RST), .Y(DFF_129_N3) );
	nor2_1 U1251( .A(RST), .B(n1433gat), .Y(DFF_128_N3) );
	nor3_1 U1252( .A(n1078), .B(RST), .C(n945), .Y(DFF_127_N3) );
	o21ai_0 U1253( .A1(n1079), .A2(n258), .B1(n895), .Y(n1078) );
	and3_1 U1254( .A(n1080), .B(n1202), .C(n1081), .X(n895) );
	nor3_1 U1255( .A(n639), .B(n1200), .C(n949), .Y(n1081) );
	mux2i_1 U1256( .A0(n1208), .A1(n1205), .S(n747), .Y(n1080) );
	nor4_1 U1257( .A(n1150), .B(n632), .C(n665), .D(n2179gat), .Y(n1079) );
	a21oi_1 U1258( .A1(n1082), .A2(n734), .B1(RST), .Y(DFF_126_N3) );
	and2_0 U1259( .A(n33), .B(n3128gat), .X(DFF_125_N3) );
	and2_0 U1260( .A(n33), .B(n3126gat), .X(DFF_124_N3) );
	and2_0 U1261( .A(n33), .B(n3127gat), .X(DFF_123_N3) );
	nor2_1 U1262( .A(RST), .B(n770), .Y(DFF_122_N3) );
	nor2_1 U1263( .A(RST), .B(n1332gat), .Y(DFF_121_N3) );
	nor3_1 U1264( .A(n1034), .B(n944), .C(n1026), .Y(DFF_120_N3) );
	nor2_1 U1265( .A(n748), .B(RST), .Y(DFF_119_N3) );
	nor2_1 U1266( .A(RST), .B(n644), .Y(DFF_118_N3) );
	nor4_1 U1267( .A(n1083), .B(n1026), .C(n1027), .D(n847), .Y(DFF_117_N3) );
	inv_1 U1268( .A(n949), .Y(n847) );
	nor2_1 U1269( .A(n1205), .B(n1208), .Y(n949) );
	nand2_1 U1270( .A(n1035), .B(n637), .Y(n1026) );
	inv_1 U1271( .A(n1029), .Y(n1035) );
	nand2_1 U1272( .A(n1084), .B(n33), .Y(n1029) );
	nand3_1 U1273( .A(n620), .B(n638), .C(n1207), .Y(n1083) );
	or3_1 U1274( .A(n32), .B(DFF_143_N3), .C(n31), .X(DFF_116_N3) );
	inv_1 U1275( .A(n1040), .Y(n31) );
	nand2_1 U1276( .A(n1206), .B(n1085), .Y(n1040) );
	nor2_1 U1277( .A(n691), .B(RST), .Y(DFF_143_N3) );
	inv_1 U1278( .A(n752), .Y(n691) );
	nand2_1 U1279( .A(n748), .B(n734), .Y(n752) );
	nand3_1 U1280( .A(n1145), .B(n1117), .C(n1038), .Y(n734) );
	inv_1 U1281( .A(n750), .Y(n748) );
	nand2_1 U1282( .A(n770), .B(n1082), .Y(n750) );
	and2_0 U1283( .A(n739), .B(n1086), .X(n1082) );
	nand4_1 U1284( .A(n1206), .B(n1038), .C(n1117), .D(n625), .Y(n1086) );
	nor2_1 U1285( .A(n1182), .B(n1181), .Y(n1038) );
	nand4_1 U1286( .A(n1182), .B(n1037), .C(n1117), .D(n624), .Y(n739) );
	nor2_1 U1287( .A(n999), .B(n975), .Y(n770) );
	and2_0 U1288( .A(n1037), .B(n1087), .X(n975) );
	nor2_1 U1289( .A(n1206), .B(n1145), .Y(n1037) );
	and3_1 U1290( .A(n1087), .B(n625), .C(n1206), .X(n999) );
	inv_1 U1291( .A(n1076), .Y(n32) );
	nand2_1 U1292( .A(n1085), .B(n627), .Y(n1076) );
	and3_1 U1293( .A(n1087), .B(n33), .C(n1145), .X(n1085) );
	nor3_1 U1294( .A(n650), .B(n1182), .C(n624), .Y(n1087) );
	nor3_1 U1295( .A(n1034), .B(RST), .C(n1088), .Y(DFF_115_N3) );
	inv_1 U1296( .A(n1053), .Y(n1088) );
	nand2_1 U1297( .A(n1031), .B(n1089), .Y(n1053) );
	nand3_1 U1298( .A(n747), .B(n1084), .C(n686), .Y(n1089) );
	nand4_1 U1299( .A(n1200), .B(n1202), .C(n1090), .D(n1205), .Y(n1034) );
	nor2_1 U1300( .A(n1207), .B(n1208), .Y(n1090) );
	nor2_1 U1301( .A(RST), .B(n646), .Y(DFF_114_N3) );
	nor2_1 U1302( .A(n618), .B(RST), .Y(DFF_113_N3) );
	nor2_1 U1303( .A(RST), .B(n641), .Y(DFF_112_N3) );
	nor2_1 U1304( .A(RST), .B(n642), .Y(DFF_111_N3) );
	nor2_1 U1305( .A(RST), .B(n619), .Y(DFF_110_N3) );
	and2_0 U1306( .A(n33), .B(n1214), .X(DFF_109_N3) );
	nor2_1 U1307( .A(RST), .B(n643), .Y(DFF_108_N3) );
	and2_0 U1308( .A(n33), .B(n1216), .X(DFF_107_N3) );
	and2_0 U1309( .A(n33), .B(n1219), .X(DFF_106_N3) );
	and2_0 U1310( .A(n33), .B(n1218), .X(DFF_105_N3) );
	inv_1 U1311( .A(RST), .Y(n33) );
	nor2_1 U1312( .A(RST), .B(n698), .Y(DFF_104_N3) );
	inv_1 U1313( .A(n3149gat), .Y(n698) );
	nand3_1 U1314( .A(n205), .B(n206), .C(n649), .Y(n3149gat) );
	nor2_1 U1315( .A(RST), .B(n696), .Y(DFF_101_N3) );
	xnor2_1 U1316( .A(n1091), .B(n1092), .Y(n696) );
	xor2_1 U1317( .A(n1216), .B(n1093), .X(n1092) );
	xor2_1 U1318( .A(n1214), .B(n1215), .X(n1093) );
	xnor2_1 U1319( .A(n1219), .B(n1094), .Y(n1091) );
	xor2_1 U1320( .A(n1217), .B(n1218), .X(n1094) );
	a21oi_1 U1321( .A1(n1095), .A2(n945), .B1(RST), .Y(DFF_100_N3) );
	inv_1 U1322( .A(n1096), .Y(n945) );
	o21ai_0 U1323( .A1(n1127), .A2(n1031), .B1(n1097), .Y(n1096) );
	mux2i_1 U1324( .A0(n1098), .A1(n1099), .S(n747), .Y(n1097) );
	nor2_1 U1325( .A(n1100), .B(n1101), .Y(n1099) );
	inv_1 U1326( .A(n1084), .Y(n1101) );
	nor2_1 U1327( .A(n1130), .B(n1128), .Y(n1084) );
	mux2i_1 U1328( .A0(n686), .A1(n1102), .S(n1103), .Y(n1100) );
	nor2_1 U1329( .A(n201), .B(n200), .Y(n1103) );
	nor2_1 U1330( .A(n637), .B(n1027), .Y(n1102) );
	and2_0 U1331( .A(n943), .B(n1127), .X(n1098) );
	nor2_1 U1332( .A(n942), .B(n1128), .Y(n943) );
	nand3_1 U1333( .A(n1128), .B(n1104), .C(n1105), .Y(n1031) );
	nor3_1 U1334( .A(n747), .B(n1130), .C(n1220), .Y(n1105) );
	inv_1 U1335( .A(n715), .Y(n747) );
	o21ai_0 U1336( .A1(n649), .A2(n226), .B1(n2102gat), .Y(n715) );
	inv_1 U1337( .A(n1027), .Y(n1104) );
	nand2_1 U1338( .A(n1221), .B(n645), .Y(n1027) );
	nor2_1 U1339( .A(n1106), .B(n896), .Y(n1095) );
	inv_1 U1340( .A(n881), .Y(n896) );
	nor4_1 U1341( .A(n1107), .B(n682), .C(n1223), .D(n1222), .Y(n881) );
	a21oi_1 U1342( .A1(n1074), .A2(n1123), .B1(n3100gat), .Y(n682) );
	and4_1 U1343( .A(n1226), .B(n1227), .C(n1108), .D(n251), .X(n1074) );
	nor2_1 U1344( .A(n1224), .B(n1225), .Y(n1108) );
	and2_0 U1345( .A(n1050), .B(n187), .X(n1107) );
	nand2_1 U1346( .A(n2021gat), .B(n649), .Y(n1050) );
	xor2_1 U1347( .A(n1109), .B(n1228), .X(n1106) );
	o211ai_1 U1348( .A1(n1220), .A2(n645), .B1(n942), .C1(n1221), .Y(n1109) );
	nand2_1 U1349( .A(n1130), .B(n686), .Y(n942) );
	nor2_1 U1350( .A(n944), .B(n637), .Y(n686) );
	nand2_1 U1351( .A(n1129), .B(n1221), .Y(n944) );
	xor2_1 troj47_0_U1( .A(tempDFF_46_N3), .B(Trigger_en_47_0), .X(DFF_46_N3) );
	and2_1 troj47_0_U2( .A(troj47_0_n1), .B(troj47_0_n2), .X(Trigger_en_47_0) );
	nor3_1 troj47_0_U3( .A(DFF_33_N3), .B(n862), .C(n1006), .Y(troj47_0_n2) );
	and3_1 troj47_0_U4( .A(DFF_56_N3), .B(DFF_122_N3), .C(n810), .X(troj47_0_n1) );
endmodule
