//****************************************************************
// TRIT-ASIC Generated Trojans.  The design generated below is for academic use only.
// Please cite the following if using the benchmark provided:
// J. Cruz, Y. Huang, P. Mishra, S. Bhunia, 
// "An Automated Configurable Trojan Insertion Framework for Dynamic Trust Benchmarks", DATE, 2018
//****************************************************************

module s38584( GND, VDD, RST, CLK, g100, g113, g114, g115, g116, g120, 
		g124, g125, g126, g127, g134, g135, g35, g36, g44, g5, 
		g53, g54, g56, g57, g64, g6744, g6745, g6746, g6747, g6748, 
		g6749, g6750, g6751, g6752, g6753, g72, g73, g84, g90, g91, 
		g92, g99, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, 
		g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, 
		g12833, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, 
		g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, 
		g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, 
		g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, 
		g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, 
		g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, 
		g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, 
		g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, 
		g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, 
		g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, 
		g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, 
		g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164, g24165, g24166, 
		g24167, g24168, g24169, g24170, g24171, g24172, g24173, g24174, g24175, g24176, 
		g24177, g24178, g24179, g24180, g24181, g24182, g24183, g24184, g24185, g25114, 
		g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, 
		g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, 
		g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, 
		g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, 
		g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, 
		g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, 
		g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, 
		g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, 
		g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, 
		g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540, g7916, 
		g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, 
		g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, 
		g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, 
		g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, 
		g9617, g9680, g9682, g9741, g9743, g9817);

	input GND, VDD, RST, CLK, g100, g113, g114, g115, g116, g120, g124, g125,
         g126, g127, g134, g135, g35, g36, g44, g5, g53, g54, g56, g57, g64,
         g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753,
         g72, g73, g84, g90, g91, g92, g99;

	output g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447,
         g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422,
         g12470, g12832, g12833, g12919, g12923, g13039, g13049, g13068,
         g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906,
         g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201,
         g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673,
         g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624,
         g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744,
         g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320,
         g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607,
         g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711,
         g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787,
         g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096,
         g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357,
         g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176,
         g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612,
         g23652, g23683, g23759, g24151, g24161, g24162, g24163, g24164,
         g24165, g24166, g24167, g24168, g24169, g24170, g24171, g24172,
         g24173, g24174, g24175, g24176, g24177, g24178, g24179, g24180,
         g24181, g24182, g24183, g24184, g24185, g25114, g25167, g25219,
         g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588,
         g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030,
         g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214,
         g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327,
         g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793,
         g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975,
         g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935,
         g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201,
         g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238,
         g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597,
         g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923,
         g34925, g34927, g34956, g34972, g7243, g7245, g7257, g7260, g7540,
         g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291,
         g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783,
         g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916,
         g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555,
         g9615, g9617, g9680, g9682, g9741, g9743, g9817;

	wire n11944, n10166, n10890, n10167, n10886, n10884, n10885, n10888, n10883, n10889, 
		n11781, n6079, n10887, n5958, n11974, n6068, n6031, n5952, n11895, n5960, 
		n11876, n11945, n5953, n6032, n11963, n5882, n10601, n10600, n10210, n11799, 
		n10603, n11955, n11892, n11859, n11775, n5955, n5872, n11936, n6066, n11907, 
		n5899, n10611, n11943, n5903, n10614, n11956, n5902, n10608, n11972, n5900, 
		n10606, n11839, n10619, n11942, n5898, n10604, n11968, n5901, n10615, n11960, 
		n5904, n10617, n10224, n10221, n10225, n10228, n10227, n10226, n10223, n10222, 
		g341, n11937, n6092, n10881, n5919, n11913, n5905, n11912, n5887, n11940, 
		n5948, n10170, n10449, n10205, n11789, n5950, n11966, n5954, n11938, n6072, 
		n10501, n11843, n6080, n10877, n10357, n11761, n6085, n10428, n11763, n6084, 
		n10882, g496, n10662, n11857, n5888, n10664, n11858, n6082, n11819, n6053, 
		n11954, n6088, n5914, n10663, n5920, n11826, n6070, n10234, n11834, n5970, 
		n11914, n5907, n11939, n6062, n10450, n5944, n19679, n11807, n6069, g933, 
		n11957, n5884, n11828, n5932, n10455, n5945, n11829, n5934, n11959, n5908, 
		n11891, n6033, n11861, n19677, n11788, n5961, g1277, n10454, n11816, n5933, 
		n11862, n5881, n11866, n6074, n11864, n5866, n11865, n5969, n11867, n6076, 
		n11869, n6077, n11863, n5871, n11868, n6075, n10665, n10453, n11897, n6064, 
		n10666, n11964, n10211, n5940, n5938, n11952, n6014, n11951, n6016, n5923, 
		n5930, n5926, n5925, n5935, n5936, n11900, n6006, n11899, n5987, n5937, 
		n11823, n6018, n11856, n6019, n10500, n11874, n5976, n11873, n5977, n5921, 
		n11811, n5973, n11875, n6010, n11850, n6011, n11883, n5979, n11817, n5980, 
		n5924, n11815, n5978, n11806, n5986, n10495, n5929, n11871, n6002, n11870, 
		n6003, n5922, n11824, n5982, n11785, n5971, n10499, n11827, n6004, n11841, 
		n6005, n10493, n11800, n5985, n10498, n5927, n11894, n6008, n11893, n5974, 
		n5928, n11833, n6012, n11851, n6013, n10494, n11903, n5993, n11902, n5972, 
		n5939, n11803, n5992, n11793, n5999, n10497, n11812, n5994, n11783, n6015, 
		n10496, n10312, n10316, n10313, n10309, n10315, n10310, n10314, n10311, n11762, 
		n6030, n11852, n6025, n11784, n5984, n11825, n6001, n10488, n11773, n6027, 
		n11853, n6026, n11792, n5989, n11782, n6024, n11813, n5995, n10486, n11772, 
		n6036, n11786, n6021, n11796, n5990, n11846, n6007, n10489, n11764, n6029, 
		n11808, n5996, n11814, n5975, n11797, n5991, n10487, n11767, n6037, n11780, 
		n6023, n11809, n5981, n11822, n6000, n10490, n11776, n6028, n11830, n5983, 
		n11820, n5997, n11770, n6034, n11804, n6022, n11778, n5998, n11805, n6020, 
		n10491, n11771, n6035, n11854, n6017, n11855, n5988, n11848, n6009, n10492, 
		n11840, n5886, n11901, n5896, n11962, n5867, g111, n11946, n5894, n5869, 
		n11920, n6048, n11921, n5873, n11904, n5890, n5864, n11926, n6049, n11927, 
		n6097, n5918, n11877, n5892, n5943, n11924, n6046, n11925, n6095, n11795, 
		n5965, n11837, n5885, g85, n11950, n5893, n11794, n5963, n5868, n11928, 
		n6047, n11929, n6093, n11953, n5891, n11836, n5964, n11958, n5889, n11849, 
		n5966, n5863, n11934, n6052, n11935, n6096, n11915, n5895, n5876, n11930, 
		n6045, n11931, n5862, n5877, n11922, n6051, n11923, n6098, n5942, n10451, 
		n11932, n6050, n11933, n6094, n10452, g4242, n5909, n10620, n10618, n5917, 
		n10616, n5916, n10613, n11791, n5962, n11842, n6063, n11948, n5941, n11947, 
		n5931, n5911, n10612, n5915, n5913, n10609, n10607, n5910, n10605, n5912, 
		g65, n11847, n5949, n5957, n5956, n11779, n11961, n6071, n11906, n5875, 
		n11777, n11872, n5874, n11898, n6073, g4531, n10667, n11967, n11973, n11941, 
		n11790, n5947, n11909, n6054, n6041, n11801, n11769, n11890, n11768, n6043, 
		n11919, n6056, n11844, n6091, n11810, n11879, n11916, n11917, n6038, n10184, 
		n11889, n6059, n11821, n11905, n11760, n5946, n11884, n6061, n11765, n6039, 
		n11831, n6081, n11910, n11802, n6042, n11878, n6057, n11888, n6089, n11766, 
		n6090, n11860, n5878, n11911, n6055, n6040, n5968, n11908, g4578, n11918, 
		n6044, n11881, n6060, n11887, n6099, n11832, n6087, n11798, n5879, n10217, 
		n11880, n6058, n10610, n11787, g4519, g4520, n5967, n5880, n5865, n5870, 
		n10213, n19467, g4480, g4495, g4498, g4501, n19451, n10880, n11896, n6067, 
		n5959, n10448, n11949, n6078, g26959, g4455, n10519, n11882, n5883, n10602, 
		n11965, g4540, g4543, g4567, g4546, n19450, g4570, g4571, n11885, n6083, 
		n5951, n11886, n6086, g4564, n11845, n10231, n11818, n6065, n10429, n11774, 
		n5897, n11838, n5906, n20311, g52, g55, n10232, g46, n11971, n11970, 
		n11835, g47, n11969, g48, g49, g45, g51, g50, n10474, n10475, 
		n10708, n10925, n10876, n10549, n10485, g25689, n10291, g24265, n10363, n10861, 
		n10862, n10860, n10355, n10421, n10713, n10589, n10395, n10540, n10544, n10563, 
		n10871, n10387, n10570, n10542, n10905, n10911, n10569, n10541, n10904, n10386, 
		n10907, n10863, n10827, n10801, n10798, n10813, n10787, n10785, n10786, n10782, 
		n10775, n10811, n10824, n10828, n10772, n10776, n10781, n10783, n10812, n10839, 
		n10837, n10838, n10749, n10746, n10750, n10830, n10833, n10831, n10832, n10808, 
		n10807, n10809, n10806, n10817, n10820, n10765, n10768, n10766, n10767, n10739, 
		n10742, n10818, n10819, n10740, n10741, n10761, n10759, n10760, n10756, n10755, 
		n10757, n10754, n10802, n10791, n10794, n10792, n10793, n10780, n10728, n10726, 
		n10729, n10727, n10730, n10733, n10737, n10731, n10732, n10623, n10626, n10634, 
		n10625, n10627, n10635, n10630, n10638, n10628, n10624, n10632, n10629, n10637, 
		n10891, n10407, n10190, n10935, n10867, n10651, n10641, n10649, n10654, n10645, 
		n10653, n10639, n10647, n10934, n10644, n10868, n10652, n10648, n10650, n10873, 
		n10929, n10933, n10578, n10701, n10709, n10858, n10682, n10162, n10599, n10596, 
		n10427, n10461, g26960, n10598, n10594, n10595, n10869, n10597, n10866, n10317, 
		n10560, n10559, n10384, n10186, n10467, n10359, n10529, n10393, n10712, n10308, 
		n10468, n10829, n10534, n10700, n10714, n10511, n10510, n10512, n10513, n10442, 
		n10734, n10689, n10464, n10230, n10535, n10229, n10573, n10706, n10721, n10723, 
		n10738, n10724, n10725, n10872, n10936, n10710, n10551, n10722, n10720, n10687, 
		n10859, n10895, n10852, n10856, n10853, n10849, n10855, n10850, n10854, n10851, 
		n10473, n10412, n10411, n10707, n10527, n10814, n10788, n10778, n10825, n10834, 
		n10769, n10771, n10747, n10743, n10823, n10745, n10810, n10799, n10795, n10797, 
		n10784, n10711, n10864, n10930, n10658, n10659, n10857, n10389, n10388, n10927, 
		n10926, n10699, n10372, n10550, n10875, n10790, n10672, n10673, n10379, n10374, 
		n10373, n10800, n10789, n10774, n10779, n10835, n10753, n10796, n10844, n10843, 
		n10735, n10846, n10736, n10586, n10848, n10516, n10894, n10591, n10303, n10893, 
		n10661, n10939, n10938, n10580, n10579, n10582, n10581, n10584, n10583, n10585, 
		n10294, n10842, n10816, n10777, n10751, n10764, n10803, n10376, n10815, n10826, 
		n10841, n10748, n10805, n10770, n10744, n10822, n10763, n10847, n10165, n10446, 
		n10445, n10762, n10840, n10773, n10836, n10804, n10821, n10752, n10758, n10436, 
		n10300, n10558, n10212, n10865, n10460, n10919, n10845, n10471, n10470, n10874, 
		n10438, g26885, n10917, n10420, n10419, n10418, n10417, n10415, n10414, n10413, 
		n10937, n10298, n10353, n10918, n10444, n10189, n10668, n10466, n10631, n10636, 
		n10469, n10255, n10715, n10521, n10916, g4467, n10390, n10394, n10400, n10561, 
		n10568, n10567, n10703, n10439, n10396, n10401, n10383, n10410, n10409, n10368, 
		n10433, n10155, n10154, n10157, n10158, n10341, n10425, n10434, n10424, n10435, 
		n10931, n10932, n10587, n10233, n10574, n10215, n10214, n10670, n10577, n10538, 
		n10477, n10482, n10483, n10479, n10480, n10481, n10462, n10296, n10523, n10525, 
		n10377, n10530, n10458, n10375, n10878, n10622, n10280, n10503, n10504, n10702, 
		n10571, n10870, n10912, n10909, n10698, n10633, n10643, n10646, n10640, n10642, 
		n10423, n10422, n10171, n10299, n10173, n10172, n10174, n10301, n10175, n10176, 
		n10476, n10307, n10397, n10562, n10408, n10564, n10539, n10566, n10565, n10381, 
		n10365, n10576, n10575, n10447, n10522, n10524, n10879, n10350, n10351, n10352, 
		n10349, n10218, n10690, n10216, n10557, n10556, n10304, n10329, n10572, n10437, 
		n10180, n10671, n10378, n10518, n10517, n10432, n10472, n10327, n10321, n10322, 
		n10325, n10319, n10324, n10505, n10683, n10928, n10655, n10704, n10716, n10913, 
		n10910, n10906, n10908, n10705, n10278, n10588, n10657, n10181, n10169, n10366, 
		n10367, n10369, n10370, n10590, n10443, n10592, n10695, n10347, n10348, n10305, 
		n10403, n10660, n10364, n10156, n10159, n10164, n10153, n10237, n10356, n10520, 
		n10441, n10440, n10431, n10430, n10688, n10656, n10371, n10416, n10343, n10177, 
		n10297, n10385, n10532, n10553, n10554, n10344, n10398, n10391, n10392, n10345, 
		n10718, n10717, n10924, n10484, n10533, n10920, n10914, n10531, n10478, n10552, 
		n10546, n10548, n10547, n10545, n10287, n10286, n10358, n10674, n10677, n10676, 
		n10678, n10681, n10679, n10675, n10680, n10339, n10306, n10285, n10426, n10258, 
		n10354, n10168, n10279, n10220, n10901, n10526, n10185, n10276, n10281, n10402, 
		n10528, n10399, n10506, n10272, n10271, n10275, n10250, n10251, n10273, n10898, 
		n10902, n10899, n10593, n10555, n10903, n10896, n10897, n10900, n10203, n10207, 
		n10206, n10201, n10208, n10209, n10463, n10465, n10274, n10295, n10270, n10621, 
		n10192, n10193, n10195, n10196, n10915, n10360, n10382, n10265, n10536, n10404, 
		n10266, n10361, n10509, n10267, n10200, n10691, n10693, n10692, n10694, n10697, 
		n10696, n10290, n10183, n10194, n10380, n10405, n10457, n10456, n10238, n10537, 
		n10515, n10282, n10257, n10346, n10245, n10277, n10283, n10922, n10669, n10284, 
		n10256, n10161, n10685, n10340, n10923, n10248, n10204, n10202, n10152, n10320, 
		n10686, n10502, n10684, n10188, n10191, n10178, n10254, n10252, n10249, n10253, 
		n10293, n10182, n10268, n10318, n10323, n10247, n10543, n10719, n10259, n10330, 
		n10219, n10199, n10198, n10151, n10406, n10160, n10362, n10239, n10240, n10243, 
		n10241, n10242, n10921, n10246, n10197, n10338, n10342, n10244, n10328, n10508, 
		n10289, n10514, n10507, n10264, n10262, n10263, n10269, n10302, n10459, n10163, 
		n10331, n10334, n10336, n10332, n10333, n10335, n10292, n10337, n10260, n10261, 
		n10288, n10179, n10326, n10187, n10236, n10235, n6437, n6196, n6197, n6203, 
		n6209, n6208, n6210, n6204, n6207, n6211, n6205, n6206, n6278, n6202, 
		n6198, n6212, n6199, n6201, n6200, n6277, n6301, n6299, n6300, n6225, 
		n6215, n6219, n6213, n6214, n6216, n6217, n6218, n6306, n6298, n6307, 
		n6220, n6295, n6297, n6296, n6230, n6237, n6235, n6227, n6238, n6234, 
		n6228, n6226, n6240, n6233, n6231, n6229, n6232, n6239, n6236, n6309, 
		n6308, n6222, n6224, n6221, n6223, n6294, n6314, n6302, n6291, n6281, 
		n6290, n6283, n6286, n6292, n6285, n6280, n6284, n6279, n6289, n6287, 
		n6282, n6293, n6288, n6313, n6312, n6303, n6305, n6304, n6310, n6311, 
		n6195, n6194, n6193, n6241, n6242, n6247, n6246, n6243, n6245, n6244, 
		n6330, n6341, n6344, n6343, n6342, n6331, n6334, n6336, n6335, n6333, 
		n6332, n6337, n6329, n6345, n6326, n6328, n6324, n6327, n6323, n6321, 
		n6325, n6318, n6315, n6317, n6316, n6322, n6320, n6319, n6338, n6339, 
		n6248, n6340, n6346, n6173, n6174, n6169, n6175, n6171, n6176, n6167, 
		n6172, n6177, n6170, n6166, n6168, n6179, n6178, n6165, n6268, n6185, 
		n6266, n6264, n6265, n6269, n6272, n6271, n6267, n6186, n6262, n6187, 
		n6270, n6184, n6188, n6263, n6180, n6181, n6164, n6189, n6182, n6249, 
		n6252, n6251, n6250, n6259, n6253, n6260, n6258, n6257, n6256, n6254, 
		n6255, n6261, n6183, n6192, n6275, n6274, n6191, n6273, n6190, n6276, 
		n6349, n6348, n6350, n6347, n6368, n6364, n6365, n6366, n6363, n6351, 
		n6367, n6362, n6361, n6352, n6359, n6358, n6357, n6355, n6354, n6356, 
		n6353, n6360, n6369, n6377, n6374, n6376, n6375, n6382, n6383, n6378, 
		n6379, n6380, n6381, n6373, n6371, n6370, n6372, n6387, n6385, n6384, 
		n6386, n5805, n6388, n5804, n6392, n6394, n6393, n5803, n6399, n5802, 
		n6403, n6402, n6401, n5801, n6411, n6413, n6412, n6415, n6418, n6417, 
		n5800, n5799, n6424, n5798, n6428, n6431, n6429, n5797, n6434, n6436, 
		n6433, n5796, n6442, n6444, n6443, n5795, n6449, n6448, n5794, n6450, 
		n5793, n6452, n5792, n6459, n5791, n6463, n6465, n6464, n5790, n6470, 
		n6469, n6474, n6475, n6473, n5789, n6481, n5788, n6487, n5787, n6488, 
		n6490, n6489, n5786, n6494, n5785, n5784, n6498, n6500, n6499, n5783, 
		n5782, n6506, n6507, n5781, n5780, n6513, n6512, n91, n6514, n5779, 
		n5778, n6515, n5777, n6518, n6521, n6519, n5776, n6525, n6527, n5775, 
		n6528, n5774, n6532, n6533, n5773, n5772, n5771, n6539, n6541, n6540, 
		n5770, n5769, n5768, n6549, n6548, n6553, n5767, n5766, n6557, n6560, 
		n6558, n5765, n6563, n5764, n6567, n6569, n6568, n5763, n6574, n6576, 
		n6578, n6572, n6580, n6581, n6575, n5762, n6589, n5761, n6593, n6595, 
		n6594, n5760, n6600, n6601, n6604, n6606, n5759, n6609, n6608, n5758, 
		n6611, n6612, n5757, n6615, n6617, n5756, n6619, n6621, n5755, n6624, 
		n6626, n6625, n5754, n5753, n6634, n6636, n6635, n5752, n6640, n6613, 
		n5751, n6642, n6644, n6643, n5750, n6649, n6651, n5749, n6656, n6655, 
		n5748, n5747, n6661, n5746, n6665, n6667, n6666, n5745, n6671, n6673, 
		n6672, n5744, n6677, n6679, n6678, n5743, n5742, n6688, n5741, n6692, 
		n6693, n6696, n5740, n6698, n6699, n6702, n5739, n6705, n5738, n6712, 
		n6710, n5737, n6717, n6718, n5736, n6722, n6724, n6723, n6726, n5735, 
		n6729, n5734, n6730, n6732, n6731, n5733, n6738, n6740, n6739, n6736, 
		n5732, n5731, n5730, n6755, n6756, n5729, n6762, n5728, n6766, n6768, 
		n6769, n6767, n6770, n5727, n6775, n6777, n6776, n5726, n6781, n6780, 
		n5725, n6786, n6788, n6787, n5724, n6792, n6791, n5723, n6796, n6798, 
		n6797, n6800, n5722, n5721, n6805, n6807, n6806, n5720, n6812, n6814, 
		n6813, n6818, n5719, n6821, n5718, n6824, n6826, n6825, n5717, n6830, 
		n6832, n5716, n6838, n6836, n5715, n6847, n6846, n6845, n6852, n6854, 
		n5714, n6855, n6857, n6856, n5713, n6860, n6862, n5712, n6866, n6867, 
		n5711, n5710, n6874, n6876, n6657, n6875, n5709, n6877, n6878, n5708, 
		n6883, n6884, n5707, n6885, n6887, n6886, n5706, n6683, n5705, n6892, 
		n5704, n6895, n6897, n6896, n5703, n6902, n6904, n6903, n5702, n6909, 
		n6908, n6912, n5701, n5700, n6915, n6914, n57, n6920, n5699, n6921, 
		n6504, n5698, n6923, n6511, n6925, n6614, n6924, n6926, n5697, n6929, 
		n6931, n6928, n5696, n5695, n6939, n6941, n6942, n6940, n6943, n5694, 
		n6945, n6947, n6946, n6670, n5693, n6949, n5692, n6953, n6955, n6954, 
		n6958, n5691, n6962, n6961, n5690, n6967, n6965, n6968, n5689, n5688, 
		n5687, n5686, n6976, n5685, n6980, n5684, n6984, n6985, n5683, n6987, 
		n5682, n6991, n6993, n6992, n5681, n6998, n7000, n6999, n6538, n5680, 
		n7001, n7003, n5679, n7006, n6547, n7008, n7007, n7009, n5678, n7012, 
		n7014, n7013, n5677, n7019, n5676, n7023, n7025, n7024, n5675, n7031, 
		n7032, n7033, n7028, n7037, n7035, n5674, n7042, n5673, n7045, n7047, 
		n6935, n7044, n5672, n7052, n7054, n7053, n7055, n5671, n5670, n7062, 
		n7065, n7063, n5669, n7067, n5668, n7068, n7070, n7069, n5667, n7073, 
		n5666, n5665, n7078, n7080, n7079, n5664, n7085, n7084, n5663, n7092, 
		n7093, n5662, n7099, n5661, n7104, n7106, n7105, n5660, n7112, n5659, 
		n7115, n5658, n7116, n7119, n7117, n5657, n5656, n5655, n5654, n7125, 
		n7127, n7126, n5653, n6447, n6445, n5652, n7135, n5651, n7140, n7139, 
		n7143, n5650, n7145, n7147, n7146, n6571, n5649, n7149, n7151, n7150, 
		n5648, n7155, n7157, n7153, n5647, n7164, n7163, n5646, n5645, n7169, 
		n7171, n7170, n5644, n7175, n7177, n7176, n5643, n7180, n5642, n7183, 
		n7185, n7184, n5641, n5640, n7188, n7190, n7189, n5639, n7193, n7195, 
		n6691, n7194, n7192, n5638, n7204, n5637, n5636, n7209, n7211, n7212, 
		n7210, n5635, n7217, n7216, n5634, n7225, n7227, n7226, n5633, n7232, 
		n7234, n7233, n5632, n7240, n5631, n7244, n6752, n7246, n7245, n7247, 
		n7243, n5630, n7250, n7252, n6542, n7251, n5629, n7256, n7255, n5628, 
		n6827, n7261, n7262, n5627, n5626, n7267, n7269, n7268, n5625, n5624, 
		n7274, n7278, n5623, n7282, n5622, n7284, n7287, n7285, n5621, n7289, 
		n7291, n7290, n6790, n5620, n7292, n7293, n5619, n7297, n5618, n5617, 
		n7301, n7304, n7302, n5616, n7309, n7311, n7295, n7310, n7314, n5615, 
		n7316, n5614, n7318, n7320, n7319, n6660, n5613, n5612, n7323, n7324, 
		n5611, n7328, n7330, n7329, n5610, n7335, n7337, n7336, n5609, n7342, 
		n7294, n5608, n7343, n7346, n7344, n5607, n7350, n7352, n7351, n5606, 
		n7357, n7356, n7355, n7361, n7363, n5605, n7364, n7366, n7365, n5604, 
		n7368, n5603, n7371, n7373, n7074, n7372, n5602, n6495, n5601, n7380, 
		n5600, n7383, n7385, n7384, n5599, n7388, n7389, n5598, n5597, n5596, 
		n7398, n7400, n7399, n5595, n5594, n7406, n7405, n5593, n5592, n5591, 
		n7415, n7417, n5590, n7421, n7423, n7420, n7422, n5589, n7426, n5588, 
		n7431, n5587, n7434, n7435, n7437, n6986, n7436, n6620, n5586, n7441, 
		n7440, n7288, n5585, n7444, n7443, n5584, n7446, n7448, n7447, n5583, 
		n7452, n7454, n7453, n7456, n6964, n5582, n7457, n7459, n7120, n7458, 
		n5581, n5580, n7467, n5579, n7470, n7471, n5578, n5577, n7476, n7478, 
		n7479, n7477, n7480, n5576, n7482, n7484, n7483, n5575, n7488, n5574, 
		n7491, n7492, n7059, n5573, n5572, n7493, n7495, n7494, n5571, n7498, 
		n7500, n7501, n7499, n5570, n7503, n7505, n7504, n5569, n7509, n7511, 
		n7507, n5568, n5567, n7517, n7518, n7516, n7521, n7520, n7519, n7524, 
		n5566, n5565, n7534, n7532, n5564, n7539, n7540, n5563, n5562, n7548, 
		n7547, n5561, n7551, n5560, n7555, n7557, n5559, n6871, n5558, n7559, 
		n7561, n7560, n5557, n7564, n5556, n7567, n7569, n7568, n5555, n5554, 
		n7575, n7577, n7576, n7101, n7574, n5553, n7582, n7580, n7583, n5552, 
		n7585, n5551, n7589, n7591, n7590, n5550, n7597, n7598, n7595, n7594, 
		n5549, n5548, n7603, n5547, n7608, n7610, n7609, n5546, n7613, n7615, 
		n7614, n5545, n7619, n7621, n7620, n5544, n7624, n7623, n7622, n7629, 
		n7631, n6623, n7438, n5543, n7634, n5542, n7637, n7639, n7165, n7638, 
		n5541, n7642, n7643, n7020, n5540, n7647, n7649, n7648, n7652, n5539, 
		n7655, n6893, n7656, n6891, n5538, n7660, n7659, n7658, n7664, n7665, 
		n5537, n7666, n7325, n5536, n5535, n7671, n7046, n7048, n7672, n7205, 
		n7675, n7678, n7677, n7681, n7680, n7679, n7676, n7686, n7685, n7684, 
		n7683, n7674, n7689, n7692, n7695, n7691, n7690, n7688, n7705, n7706, 
		n7704, n7203, n7703, n7673, n5534, n7711, n7712, n5533, n7714, n7715, 
		n5532, n7719, n7721, n7720, n7717, n5531, n5530, n7726, n5529, n7728, 
		n7730, n7729, n6907, n5528, n7733, n7735, n7734, n5527, n5526, n7740, 
		n7741, n5525, n7745, n5524, n7748, n7750, n7749, n5523, n7753, n7754, 
		n7018, n7751, n5522, n5521, n7759, n5520, n7762, n7764, n7763, n7765, 
		n7761, n5519, n7771, n5518, n5517, n7061, n5516, n5515, n7779, n7780, 
		n6493, n5514, n7783, n7784, n7786, n7785, n7789, n6716, n7403, n5513, 
		n7792, n5512, n7797, n7713, n5511, n5510, n7800, n7801, n5509, n7805, 
		n7807, n7806, n5508, n7810, n7812, n7811, n5507, n7816, n7818, n7817, 
		n5506, n7819, n7821, n6782, n7820, n7823, n6783, n5505, n7829, n7831, 
		n7830, n7827, n5504, n7837, n7839, n7838, n5503, n7842, n7844, n7843, 
		n5502, n7847, n7849, n7848, n5501, n5500, n7851, n7853, n7854, n7852, 
		n5499, n7856, n7859, n7858, n7857, n7864, n5498, n7865, n7162, n7641, 
		n7640, n7710, n7636, n5497, n7868, n7867, n64, n7866, n62, n7510, 
		n5496, n7869, n5495, n5494, n7872, n7874, n7873, n5493, n7877, n7879, 
		n7878, n5492, n7882, n5491, n7888, n7889, n7890, n7885, n7894, n7892, 
		n5490, n7897, n5489, n7900, n7902, n7901, n5488, n7906, n7904, n5487, 
		n7910, n5486, n5485, n5484, n7913, n5483, n7915, n5482, n5481, n6658, 
		n5480, n7919, n7920, n5479, n5478, n7925, n7924, n7923, n7927, n7928, 
		n5477, n7929, n7931, n7933, n7932, n7930, n7937, n7936, n7939, n5476, 
		n7942, n7944, n7945, n7943, n5475, n7948, n7950, n7949, n5474, n7951, 
		n5473, n7953, n7952, n5472, n7958, n7960, n7959, n5471, n7962, n7964, 
		n7963, n5470, n7967, n5469, n7970, n7969, n7973, n5468, n7975, n7977, 
		n7978, n7976, n7979, n7755, n7752, n5467, n7778, n5466, n7980, n7982, 
		n7981, n5465, n5464, n7986, n7988, n7987, n5463, n7990, n7992, n7991, 
		n5462, n7994, n7996, n7995, n5461, n8000, n8001, n5460, n8003, n6849, 
		n8004, n7475, n8002, n6848, n7481, n6851, n5459, n8007, n8009, n7077, 
		n8006, n5458, n8011, n8013, n8012, n5457, n8016, n8018, n8017, n7841, 
		n5456, n8021, n8022, n5455, n8026, n8028, n8027, n5454, n8030, n5453, 
		n8034, n5452, n8038, n8040, n8039, n5451, n8044, n8046, n8045, n7231, 
		n5450, n8050, n8052, n8055, n5449, n8057, n8059, n8058, n5448, n8063, 
		n8065, n8064, n5447, n8066, n8068, n8067, n5446, n5445, n8071, n8073, 
		n8072, n5444, n8076, n6918, n5443, n8079, n8081, n8080, n5442, n8086, 
		n8087, n8084, n8091, n8090, n5441, n5440, n8096, n8098, n8097, n5439, 
		n8102, n8100, n8104, n5438, n6784, n5437, n8108, n8109, n7651, n5436, 
		n8112, n5435, n8117, n8115, n8116, n5434, n8119, n8121, n8019, n7428, 
		n8120, n5433, n5432, n8124, n8126, n8122, n5431, n6697, n6510, n5430, 
		n5429, n8132, n8134, n8133, n5428, n8136, n8138, n8137, n5427, n8143, 
		n8141, n5426, n8150, n6551, n8149, n8152, n6555, n5425, n8155, n8157, 
		n8156, n5424, n8159, n8158, n5423, n8163, n8165, n8164, n5422, n8168, 
		n5421, n8172, n7242, n5420, n8176, n8178, n8177, n7538, n5419, n7312, 
		n5418, n5417, n8184, n8183, n5416, n8188, n8190, n8189, n5415, n8192, 
		n5414, n8195, n5413, n8197, n8199, n8198, n7508, n5412, n8202, n6529, 
		n5411, n8205, n5410, n8207, n8206, n5409, n8210, n8212, n8211, n5408, 
		n8214, n8216, n8215, n7698, n5407, n8219, n5406, n8222, n5405, n8227, 
		n8230, n8228, n5404, n5403, n8233, n8235, n7562, n8234, n5402, n6764, 
		n8237, n5401, n8241, n6844, n5400, n8243, n8245, n8244, n5399, n8246, 
		n7845, n5398, n8247, n8249, n8248, n5397, n8254, n8255, n8253, n8252, 
		n5396, n7376, n7644, n7374, n7075, n7375, n5395, n7798, n7315, n5394, 
		n8257, n8258, n8054, n5393, n8263, n8265, n8264, n5392, n8269, n5391, 
		n8271, n6425, n8272, n5390, n8275, n8277, n8276, n5389, n8279, n8281, 
		n8280, n8284, n5388, n8288, n5387, n8291, n8293, n8292, n5386, n8295, 
		n8296, n5385, n5384, n5383, n8305, n8307, n7602, n8306, n5382, n8310, 
		n8312, n8311, n7103, n5381, n8315, n7102, n8314, n5380, n8317, n5379, 
		n8320, n8322, n8321, n5378, n8325, n5377, n8329, n5376, n5375, n8335, 
		n8337, n8336, n5374, n8338, n8340, n8339, n5373, n8344, n7317, n5372, 
		n8346, n8349, n8347, n5371, n8354, n8356, n8174, n8355, n5370, n8359, 
		n8360, n8363, n5369, n8364, n5368, n8368, n8370, n8369, n5367, n5366, 
		n5365, n8374, n8193, n8376, n8375, n8378, n5364, n8379, n5363, n8382, 
		n8381, n5362, n8386, n8387, n5361, n8389, n8390, n8392, n8391, n7907, 
		n7908, n7905, n5360, n8401, n8402, n8377, n7565, n7758, n7757, n5359, 
		n8405, n8407, n8410, n5358, n7308, n7159, n8181, n5357, n8414, n6509, 
		n8413, n8130, n5356, n8415, n8417, n6516, n8416, n5355, n8422, n8421, 
		n5354, n8426, n8428, n8430, n8425, n8432, n8433, n6561, n8427, n5353, 
		n8438, n8439, n8436, n5352, n8442, n8444, n8443, n5351, n8445, n8447, 
		n7645, n8446, n8449, n5350, n8451, n6451, n8450, n5349, n8455, n8457, 
		n8456, n5348, n8461, n7654, n5347, n5346, n8462, n8464, n6522, n6456, 
		n8463, n5345, n8182, n5344, n8468, n8470, n7339, n8466, n5343, n8475, 
		n8477, n8478, n8476, n8479, n8129, n8123, n5342, n8480, n8481, n5341, 
		n5340, n8488, n8487, n5339, n5338, n5337, n8492, n8494, n8496, n8491, 
		n8497, n8498, n8493, n5336, n8504, n6706, n5335, n7828, n8505, n5334, 
		n5333, n5332, n5331, n8511, n8513, n8512, n5330, n8515, n8517, n8516, 
		n5329, n8524, n8522, n5328, n5327, n8531, n8529, n8534, n8533, n8049, 
		n5326, n8538, n5325, n8543, n8545, n8544, n6687, n5324, n8546, n8548, 
		n8547, n5323, n8552, n8554, n8555, n8553, n8556, n7160, n7154, n5322, 
		n8559, n5321, n8562, n8564, n8563, n8566, n8561, n5320, n8569, n8571, 
		n6868, n8570, n8140, n5319, n8575, n8574, n8573, n8576, n8577, n5318, 
		n8578, n5317, n8580, n6531, n8579, n5316, n7429, n8581, n7461, n5315, 
		n8582, n8584, n5314, n5313, n5312, n8589, n8590, n7918, n5311, n5310, 
		n8592, n5309, n8595, n8594, n5308, n8597, n8599, n5307, n8601, n8602, 
		n6689, n5306, n5305, n8605, n8607, n8606, n8459, n5304, n8611, n8613, 
		n8612, n5303, n8617, n8616, n5302, n5301, n8621, n6837, n8620, n8624, 
		n8623, n8358, n5300, n6396, n8629, n5299, n8632, n8633, n8631, n5298, 
		n5297, n8637, n8639, n8640, n8638, n5296, n7581, n8644, n7896, n5295, 
		n8646, n8648, n8647, n5294, n8650, n8651, n8652, n7381, n5293, n8656, 
		n8658, n8657, n8308, n5292, n5291, n8662, n8596, n8618, n5290, n8665, 
		n8666, n5289, n8667, n5288, n8669, n8671, n8670, n7808, n5287, n8672, 
		n6719, n7187, n5286, n8674, n8676, n8675, n8679, n5285, n8681, n8110, 
		n5284, n8682, n8684, n8685, n8683, n8686, n8441, n6759, n8437, n5283, 
		n7870, n5282, n8689, n5281, n8691, n8692, n7514, n5280, n5279, n8696, 
		n8423, n8694, n8697, n6802, n6795, n5278, n8700, n8654, n8701, n8653, 
		n8702, n8704, n8703, n8707, n6816, n8709, n8711, n8713, n8712, n8710, 
		n5277, n8715, n8717, n8716, n8720, n5276, n8724, n8727, n6389, n8725, 
		n8721, n5275, n8728, n8730, n6950, n8729, n6948, n5274, n8733, n5273, 
		n8736, n8737, n5272, n8739, n7051, n8741, n8740, n7058, n5271, n8743, 
		n5270, n8746, n8748, n8747, n5269, n5268, n8750, n8751, n7156, n8077, 
		n5267, n7650, n6622, n5266, n8755, n8757, n8756, n5265, n5264, n5263, 
		n8763, n6605, n8765, n8768, n8767, n8772, n8771, n8770, n8766, n8778, 
		n8777, n8776, n8764, n8780, n8783, n8785, n8782, n8781, n6497, n6675, 
		n8773, n8779, n8792, n7201, n8774, n8793, n8791, n6872, n8790, n6543, 
		n6602, n6603, n7196, n8762, n5262, n8795, n6654, n6471, n6478, n6477, 
		n5261, n8796, n8797, n8798, n8800, n7739, n5260, n6652, n5259, n8805, 
		n7141, n5258, n8806, n8808, n8809, n8810, n8807, n5257, n8814, n8816, 
		n7442, n8819, n7286, n8815, n7439, n5256, n8820, n8822, n8823, n8821, 
		n8035, n5255, n5254, n8827, n8828, n6641, n6793, n8826, n5253, n8834, 
		n8832, n5252, n8837, n7473, n5251, n7646, n8753, n7653, n8434, n5250, 
		n8839, n5249, n8842, n8844, n8845, n8843, n5248, n5247, n8850, n6460, 
		n6462, n8849, n6461, n5246, n8855, n5245, n8856, n6454, n5244, n8857, 
		n8859, n8858, n6997, n5243, n8860, n5242, n8862, n8863, n6535, n8861, 
		n8864, n5241, n7699, n5240, n8865, n8867, n8866, n5239, n8870, n8471, 
		n8719, n5238, n8872, n8874, n8873, n5237, n8878, n8879, n7121, n8876, 
		n8883, n7432, n8882, n5236, n5235, n5234, n8889, n5233, n8892, n5232, 
		n7670, n8161, n5231, n8448, n7530, n7529, n8893, n5230, n8894, n5229, 
		n8898, n8899, n8901, n8404, n8900, n8895, n5228, n8907, n7489, n7486, 
		n5227, n8910, n8911, n7249, n6468, n5226, n8914, n8913, n7738, n5225, 
		n8915, n8917, n7916, n8916, n8465, n5224, n8918, n8920, n6501, n8919, 
		n7191, n5223, n8922, n8924, n8923, n5222, n8500, n5221, n5220, n8927, 
		n8929, n8928, n8083, n5219, n8932, n8934, n8933, n5218, n6863, n5217, 
		n8938, n8940, n8939, n5216, n8943, n8945, n8944, n5215, n8946, n8948, 
		n8947, n5214, n8952, n8954, n7066, n8499, n8953, n5213, n8956, n8957, 
		n7552, n5212, n8961, n5211, n8963, n6432, n7221, n5210, n5209, n8966, 
		n8968, n8967, n5208, n8969, n7390, n7276, n8971, n7391, n8970, n7275, 
		n7393, n7788, n8972, n7392, n7280, n6484, n5207, n5206, n8977, n8979, 
		n7331, n8978, n7326, n5205, n8983, n8984, n8982, n8981, n5204, n5203, 
		n5202, n8988, n8987, n5201, n5200, n8990, n8992, n8991, n5199, n7743, 
		n7770, n5198, n8994, n7781, n6491, n5197, n8997, n8996, n5196, n8999, 
		n8695, n9001, n9000, n9002, n8998, n5195, n9005, n9006, n9004, n9003, 
		n7601, n5194, n5193, n5192, n9011, n9013, n9012, n6676, n5191, n9014, 
		n9015, n6662, n5190, n9018, n9020, n9019, n5189, n9022, n5188, n9025, 
		n9026, n6898, n6972, n7409, n5187, n9029, n9030, n6938, n9028, n6944, 
		n7663, n5186, n9031, n9033, n9032, n9036, n6735, n5185, n9039, n9041, 
		n9040, n9037, n5184, n9045, n6969, n9044, n6970, n5183, n9047, n9049, 
		n9048, n7876, n5182, n9051, n9052, n5181, n5180, n9055, n5179, n9059, 
		n9060, n9062, n6829, n9061, n8835, n8836, n8833, n9058, n5178, n6631, 
		n5177, n9070, n5176, n9073, n9072, n5175, n9078, n9080, n9081, n9079, 
		n9082, n5174, n9088, n9089, n9090, n9085, n9094, n9092, n5173, n9096, 
		n9098, n8659, n8908, n9097, n5172, n9099, n7632, n5171, n9101, n9103, 
		n9102, n8309, n5170, n9106, n9105, n7463, n5169, n7815, n8403, n7813, 
		n5168, n9109, n9111, n9110, n8744, n9112, n5167, n9114, n6590, n9115, 
		n7360, n7137, n6587, n5166, n9118, n6648, n9117, n5165, n9122, n9124, 
		n9123, n5164, n5163, n9126, n9127, n8330, n9131, n9134, n9133, n9138, 
		n9137, n9136, n9132, n9144, n9143, n9142, n9130, n9147, n9150, n9153, 
		n9149, n7382, n9148, n6990, n9146, n9161, n9152, n9162, n9160, n8328, 
		n8075, n7917, n9159, n6682, n9129, n9164, n5162, n5161, n8668, n5160, 
		n7984, n7744, n5159, n9167, n5158, n9168, n9169, n5157, n9171, n9172, 
		n9170, n6834, n5156, n9177, n5155, n9180, n6754, n5154, n8891, n5153, 
		n9183, n9186, n9185, n7411, n9187, n6977, n9184, n9182, n5152, n9188, 
		n5151, n9189, n9191, n9190, n5150, n9193, n7057, n9194, n9192, n8290, 
		n5149, n9196, n9198, n9197, n5148, n9201, n9200, n5147, n9204, n9205, 
		n9207, n6618, n9206, n5146, n9210, n5145, n9215, n9216, n9154, n9214, 
		n5144, n5143, n5142, n9219, n5141, n5140, n9221, n9223, n9222, n5139, 
		n8094, n5138, n9226, n9228, n9227, n9100, n5137, n9231, n8236, n5136, 
		n9232, n9234, n7983, n9233, n7985, n5135, n9236, n9238, n9239, n6779, 
		n6774, n9237, n9240, n6419, n6778, n6421, n5134, n9242, n5133, n9244, 
		n9246, n6963, n9245, n6960, n5132, n5131, n9249, n9251, n9250, n6639, 
		n5130, n9253, n9252, n5129, n9255, n9257, n9256, n5128, n9260, n5127, 
		n7144, n9265, n9267, n9266, n5126, n9269, n6983, n9271, n7523, n9270, 
		n9273, n5125, n7630, n9275, n9274, n5124, n9277, n9278, n5123, n9280, 
		n5122, n9284, n9286, n9285, n5121, n9290, n9289, n5120, n9293, n9295, 
		n7485, n9294, n5119, n9296, n9297, n5118, n9298, n9300, n9299, n7709, 
		n5117, n8557, n5116, n9304, n9305, n9306, n9302, n9309, n7039, n7600, 
		n6453, n9308, n7914, n5115, n9310, n9312, n9311, n7224, n5114, n9313, 
		n7138, n7136, n7536, n5113, n9317, n9319, n9318, n8951, n5112, n9321, 
		n9301, n8527, n8560, n5111, n9324, n9326, n6455, n9325, n6853, n5110, 
		n9327, n9329, n9328, n7322, n5109, n9330, n9331, n9332, n9334, n5108, 
		n9336, n9338, n9337, n8239, n7587, n9335, n5107, n9340, n6597, n5106, 
		n5105, n9341, n9343, n7111, n9342, n5104, n9344, n9346, n9345, n7181, 
		n5103, n9349, n9351, n9353, n9348, n9354, n9355, n7313, n8412, n9350, 
		n5102, n9357, n9359, n9358, n8042, n5101, n9361, n5100, n9364, n9363, 
		n5099, n9367, n7796, n9369, n9368, n9370, n8060, n5098, n9371, n9372, 
		n8362, n5097, n8373, n5096, n9010, n9374, n8526, n8302, n6534, n8962, 
		n8301, n5095, n9376, n6441, n6446, n7133, n5094, n5093, n9379, n9381, 
		n7803, n9380, n9383, n5092, n9384, n7202, n9386, n9385, n6695, n7050, 
		n7200, n7199, n8775, n6694, n5091, n9391, n5090, n9393, n8802, n9395, 
		n9394, n8803, n5089, n9396, n5088, n9397, n5087, n9399, n9401, n9403, 
		n9398, n9404, n9405, n7022, n7528, n9400, n5086, n7206, n5085, n8732, 
		n8603, n8731, n6951, n7946, n5084, n9411, n9412, n9409, n9413, n5083, 
		n9414, n9416, n9415, n8037, n5082, n9418, n9419, n8409, n5081, n6400, 
		n6398, n9422, n8061, n8062, n9423, n6395, n7635, n6638, n8366, n5080, 
		n7348, n9427, n9426, n5079, n9430, n9429, n9433, n5078, n5077, n9436, 
		n9437, n5076, n9439, n9441, n7332, n7410, n9440, n8029, n5075, n5074, 
		n9443, n9445, n6808, n9444, n5073, n9448, n9449, n9447, n5072, n9451, 
		n9453, n9452, n5071, n6646, n6794, n9456, n5070, n7667, n7408, n5069, 
		n9457, n9459, n9458, n5068, n5067, n6869, n5066, n9465, n9464, n9463, 
		n9466, n9467, n7086, n9071, n9247, n6745, n5065, n9469, n9471, n9470, 
		n9472, n8568, n9468, n5064, n9473, n8738, n8909, n8735, n9230, n5063, 
		n9475, n9281, n9476, n5062, n9480, n5061, n9483, n9485, n7731, n9484, 
		n5060, n9487, n9489, n9488, n5059, n9490, n9491, n5058, n5057, n8687, 
		n5056, n9495, n9497, n8023, n9496, n6664, n5055, n9498, n9500, n6789, 
		n6865, n9499, n7782, n5054, n5053, n9503, n8127, n9504, n8125, n9314, 
		n5052, n9505, n9507, n6727, n6416, n7515, n9508, n6773, n6410, n9506, 
		n9509, n8811, n7271, n7273, n7266, n6725, n7265, n8813, n9410, n7272, 
		n6721, n7270, n5051, n9511, n9493, n8660, n8690, n5050, n9514, n5049, 
		n5048, n9516, n5047, n5046, n9518, n9520, n6971, n6899, n7668, n9519, 
		n7846, n5045, n5044, n9521, n9523, n9522, n5043, n9526, n9528, n9530, 
		n7460, n9525, n9531, n9532, n7566, n7756, n9527, n5042, n5041, n9537, 
		n9539, n6570, n9538, n7148, n5040, n9541, n9543, n9542, n5039, n9546, 
		n9547, n5038, n9549, n5037, n9552, n7556, n9554, n5036, n9556, n9555, 
		n5035, n9558, n8935, n9560, n9559, n8936, n5034, n9561, n9563, n9562, 
		n9565, n8759, n5033, n9567, n5032, n5031, n5030, n9572, n9574, n6530, 
		n8203, n9576, n9573, n8959, n5029, n9580, n5028, n9582, n5027, n9583, 
		n5026, n9585, n9434, n5025, n9588, n7370, n7369, n9589, n9587, n5024, 
		n9590, n9592, n7669, n9591, n5023, n5022, n9595, n9597, n8503, n9596, 
		n6708, n7716, n9594, n7661, n6709, n5021, n8550, n8824, n9016, n8549, 
		n8036, n9599, n5020, n9601, n9603, n9602, n9292, n5019, n9604, n9606, 
		n9605, n9609, n9608, n8371, n5018, n9611, n9613, n6627, n9612, n9254, 
		n5017, n9614, n9616, n7026, n9615, n5016, n9619, n9621, n9620, n8942, 
		n5015, n9622, n7397, n9624, n8604, n9623, n9625, n7396, n7395, n5014, 
		n9627, n9629, n9628, n5013, n5012, n9633, n5011, n9635, n9634, n5010, 
		n9636, n7606, n9638, n7005, n9637, n9639, n5009, n9640, n9642, n9641, 
		n5008, n5007, n9646, n9644, n6919, n8460, n5006, n9649, n9113, n9460, 
		n9035, n6733, n9034, n9651, n9650, n9108, n6734, n9652, n9653, n7727, 
		n9461, n5005, n9656, n6439, n7131, n7129, n9050, n7401, n9658, n9657, 
		n7130, n6440, n6438, n9659, n9660, n7791, n6435, n6713, n7790, n7128, 
		n5004, n9662, n8170, n9663, n6859, n5003, n9665, n8530, n9664, n5002, 
		n9666, n9668, n6995, n9024, n9667, n7947, n5001, n5000, n9670, n9502, 
		n9672, n8274, n9671, n9673, n9669, n8273, n8160, n50, n9675, n8799, 
		n9677, n9680, n9679, n9683, n9682, n9681, n9678, n9689, n9688, n9687, 
		n9676, n9691, n9694, n9696, n8535, n9693, n7354, n6900, n9692, n6894, 
		n7349, n9684, n9690, n9703, n8261, n9685, n9704, n8260, n8053, n9702, 
		n7989, n7850, n8801, n9701, n7333, n7804, n9686, n8056, n8051, n9705, 
		n8259, n9707, n9674, n4999, n9709, n9711, n9710, n4998, n9712, n9714, 
		n9713, n8095, n7707, n4997, n9715, n9717, n9716, n7362, n4996, n4995, 
		n9720, n9722, n9721, n4994, n9727, n9647, n9725, n7550, n9643, n4993, 
		n9732, n9733, n7563, n6765, n9731, n6772, n4992, n4991, n4990, n9736, 
		n9738, n9737, n9279, n4989, n6737, n8840, n8474, n6747, n9739, n7088, 
		n6742, n4988, n9743, n9745, n9744, n9746, n9742, n4987, n9747, n4986, 
		n9749, n9751, n9753, n9748, n9754, n9755, n9756, n9750, n4985, n4984, 
		n9758, n9760, n7506, n8980, n9759, n4983, n4982, n8024, n8187, n4981, 
		n9763, n4980, n9764, n9766, n9765, n9768, n4979, n9770, n9772, n9217, 
		n4978, n9774, n6916, n9773, n9179, n4977, n9776, n9777, n9779, n8521, 
		n9778, n7974, n4976, n4975, n4974, n9786, n9788, n9787, n8319, n9724, 
		n4973, n7056, n8287, n8286, n9790, n8742, n4972, n9791, n7094, n9793, 
		n7095, n9792, n4971, n4970, n9767, n9477, n4969, n9794, n8636, n8643, 
		n8642, n9795, n4968, n9796, n8583, n6982, n6981, n7345, n9797, n9798, 
		n9272, n8440, n4967, n9799, n4966, n9801, n8912, n9202, n4965, n9804, 
		n6598, n9803, n6599, n4964, n9806, n9808, n9807, n4963, n9809, n7036, 
		n7030, n7040, n7427, n7347, n7522, n7029, n7472, n8726, n7525, n9812, 
		n7527, n4962, n7173, n7004, n7172, n7168, n8242, n7578, n6890, n4961, 
		n7469, n9814, n9817, n7083, n4960, n9819, n9820, n4959, n9821, n7725, 
		n9564, n8758, n4958, n9823, n9825, n8074, n9021, n7386, n9824, n9163, 
		n4957, n4956, n9827, n7002, n6520, n9828, n6577, n4955, n9833, n6932, 
		n9835, n6930, n9834, n7694, n7682, n6933, n6927, n9832, n6936, n9836, 
		n8985, n4954, n9840, n6650, n9446, n4953, n9841, n8706, n8705, n7769, 
		n9655, n4952, n7283, n4951, n9844, n9846, n9845, n7142, n4950, n9848, 
		n9333, n9850, n9853, n9852, n9856, n9855, n9854, n9851, n9859, n9858, 
		n9857, n9849, n9861, n9864, n9867, n9866, n9863, n7607, n9862, n9860, 
		n9874, n9421, n8904, n9875, n9420, n8905, n9873, n8267, n9872, n9482, 
		n6901, n8906, n8411, n8406, n9847, n4949, n9881, n8256, n9882, n9880, 
		n4948, n9883, n6989, n4947, n4946, n8025, n4945, n9886, n9888, n9887, 
		n9890, n4944, n9891, n4943, n9893, n9895, n7229, n9212, n9894, n8154, 
		n4942, n9896, n4941, n8708, n9632, n4940, n7774, n4939, n7775, n6817, 
		n7746, n6815, n4938, n4937, n4936, n9900, n8118, n9728, n9898, n9729, 
		n7531, n9901, n9899, n8114, n4935, n9904, n7809, n4934, n4933, n9906, 
		n9907, n9909, n9141, n9140, n9908, n9769, n9139, n8145, n8148, n8327, 
		n9771, n8331, n9128, n9912, n8142, n4932, n9915, n9917, n7799, n9916, 
		n9918, n9914, n4931, n9919, n9921, n9920, n8931, n4930, n9922, n9924, 
		n6466, n9923, n4929, n8380, n4928, n9926, n4927, n9929, n9570, n9931, 
		n6720, n9930, n9932, n4926, n9933, n9935, n9934, n4925, n7239, n9938, 
		n7824, n8357, n9937, n9936, n4924, n9382, n9939, n4923, n9941, n4922, 
		n6408, n8101, n7097, n9781, n9946, n7096, n7091, n9945, n4921, n9948, 
		n8841, n8848, n8847, n9949, n9879, n8902, n9950, n9557, n4920, n6956, 
		n9951, n4919, n9953, n9955, n9952, n9954, n4918, n9957, n9942, n9944, 
		n9956, n6537, n9943, n4917, n7110, n7113, n9960, n4916, n9964, n4915, 
		n6839, n9966, n8897, n6841, n8896, n9965, n6843, n9967, n9968, n4914, 
		n9970, n9972, n7760, n9533, n7433, n8880, n8877, n7118, n9973, n9529, 
		n9492, n9535, n9976, n9971, n7462, n4913, n9977, n61, n6485, n7281, 
		n7387, n4912, n9978, n7122, n9980, n9979, n9981, n9225, n9581, n9121, 
		n9120, n9224, n4911, n9984, n4910, n9988, n9987, n4909, n4908, n9989, 
		n4907, n7940, n9991, n4906, n8565, n9993, n9992, n9994, n4905, n9995, 
		n9997, n8266, n9209, n7611, n9996, n9486, n4904, n4903, n9038, n8958, 
		n8955, n9998, n4902, n9999, n10001, n6492, n10000, n8610, n4901, n10002, 
		n4900, n4899, n10003, n6861, n9617, n4898, n4897, n10005, n10007, n7880, 
		n6858, n10006, n4896, n4895, n10010, n10012, n10011, n4894, n7718, n10016, 
		n4893, n10017, n10019, n10018, n7451, n4892, n10021, n10023, n10022, n7899, 
		n7700, n4891, n4890, n10025, n10026, n9263, n10029, n10032, n10031, n10035, 
		n10034, n10033, n10030, n10038, n10037, n10036, n10028, n10040, n10043, n10046, 
		n10042, n10041, n8078, n10039, n10054, n10045, n8395, n10055, n10053, n9259, 
		n6629, n10052, n9258, n7881, n10027, n10056, n7213, n4889, n6801, n10058, 
		n9432, n10057, n8722, n8567, n10059, n8698, n4888, n10004, n8699, n7922, 
		n8424, n4887, n4886, n10062, n7662, n10061, n7487, n9377, n7307, n4885, 
		n10064, n10066, n10065, n4884, n7263, n4883, n4882, n10071, n10073, n8082, 
		n10072, n9283, n4881, n10074, n10076, n10075, n9631, n4880, n10079, n9023, 
		n6680, n10080, n9158, n6809, n4879, n10082, n4878, n10083, n8818, n10085, 
		n10084, n9982, n8318, n6645, n6647, n8232, n7207, n8831, n4877, n10087, 
		n10089, n6744, n6588, n10088, n7794, n6591, n10086, n7358, n7795, n7954, 
		n6746, n4876, n10092, n10094, n7903, n6668, n9056, n10093, n9494, n4875, 
		n10095, n10097, n10096, n8294, n4874, n10099, n6758, n6757, n6753, n7836, 
		n8506, n4873, n9347, n10101, n10100, n7182, n7502, n6704, n4872, n4871, 
		n10104, n4870, n10107, n10108, n10111, n9262, n9261, n8388, n8398, n4869, 
		n10113, n10115, n10114, n10116, n7767, n10112, n4868, n10118, n9735, n10117, 
		n9734, n4867, n6632, n7776, n6630, n10119, n10120, n10122, n7545, n6811, 
		n4866, n10123, n10125, n6502, n9802, n10124, n6503, n4865, n10127, n9963, 
		n9816, n6405, n88, n4864, n10129, n10130, n10128, n9544, n9545, n4863, 
		n4862, n4861, n4860, n10137, n4859, n8673, n6476, n8383, n8384, n4858, 
		n9515, n4857, n6479, n4856, n10138, n9610, n8608, n8458, n10140, n10139, 
		n8609, n4855, n10142, n10143, n10110, n9175, n10144, n8397, n10047, n8394, 
		n4854, n10146, n10148, n9784, n8587, n10147, n7123, n4853, n10149, n7616, 
		n10150, n6564, n7617, n4852, n8282, n10892, n10940, n8283, n9199, n4851, 
		n10942, n7860, n10944, n7862, n7861, n10943, n7863, n10946, n10949, n7060, 
		n10948, n10947, n7855, n10941, n4850, n8591, n7893, n10950, n9235, n4849, 
		n10952, n10954, n10953, n4848, n8761, n4847, n10956, n10958, n10957, n4846, 
		n10961, n10963, n10962, n4845, n6628, n8887, n4844, n10965, n8752, n7657, 
		n10966, n6973, n7158, n8551, n7161, n7220, n4843, n10967, n10969, n7015, 
		n9986, n10968, n8645, n4842, n10970, n10972, n8139, n10971, n4841, n10069, 
		n8107, n4840, n7571, n7573, n7572, n6554, n6550, n4839, n8655, n4838, 
		n10976, n10979, n10978, n10977, n10982, n4837, n8010, n10984, n10983, n85, 
		n8300, n8008, n4836, n10985, n9211, n6905, n10986, n9892, n7027, n4835, 
		n10987, n10989, n10988, n10070, n7497, n4834, n10990, n10992, n6681, n8558, 
		n10991, n8162, n6996, n4833, n10994, n10993, n4832, n10995, n8454, n10997, 
		n10996, n10998, n10141, n7997, n8278, n7592, n10067, n7107, n8313, n9104, 
		n9229, n8678, n8677, n7998, n4831, n11002, n11003, n10999, n7108, n11000, 
		n11001, n4830, n8641, n6546, n6545, n7258, n4829, n11007, n9057, n11008, 
		n7702, n4828, n11009, n8754, n11011, n11010, n8486, n11012, n9822, n10959, 
		n8634, n11013, n7043, n10134, n11014, n10135, n8485, n11016, n11015, n7935, 
		n7367, n10960, n4827, n11017, n11019, n11018, n4826, n4825, n11022, n11021, 
		n4824, n8144, n11025, n8146, n11027, n11024, n11023, n7197, n8147, n11026, 
		n4823, n8005, n7605, n7604, n6584, n6579, n6582, n9303, n11030, n6585, 
		n9829, n11031, n6583, n4822, n4821, n11033, n11035, n11034, n4820, n9959, 
		n11038, n9958, n9940, n4819, n11039, n11041, n7965, n6480, n7321, n11040, 
		n4818, n11042, n11044, n11043, n4817, n11045, n9540, n11047, n8520, n11046, 
		n10132, n11048, n9435, n10131, n8518, n9438, n11049, n7424, n11050, n9783, 
		n7971, n9782, n4816, n4815, n11053, n9462, n11052, n8993, n7558, n9762, 
		n4814, n7544, n7513, n7512, n4813, n11054, n11055, n6711, n4812, n11056, 
		n11058, n9320, n9961, n7883, n11057, n4811, n4810, n8467, n8472, n11059, 
		n8871, n9568, n6565, n4809, n11062, n8221, n8350, n8218, n8352, n11063, 
		n9455, n4808, n11065, n11067, n8015, n9474, n8431, n9007, n11068, n11069, 
		n8723, n8734, n6559, n11070, n8429, n8435, n11071, n11066, n4807, n11072, 
		n11074, n8191, n8888, n7496, n8171, n11073, n8930, n4806, n11075, n6831, 
		n9173, n6835, n9063, n11077, n9388, n9706, n11078, n11076, n9178, n11081, 
		n11084, n11083, n11087, n11086, n11085, n11082, n11090, n11089, n11088, n11080, 
		n11092, n11095, n11098, n11097, n11094, n8937, n7747, n11093, n7017, n8649, 
		n11091, n11106, n11099, n9065, n11107, n9174, n9066, n11105, n9176, n9761, 
		n7961, n11104, n8749, n9067, n11079, n11110, n7466, n4805, n11111, n11113, 
		n11112, n6423, n4804, n7254, n6467, n8482, n9203, n9027, n4803, n10050, 
		n4802, n11114, n11116, n8208, n11115, n7215, n7909, n7208, n7214, n8393, 
		n11118, n11117, n4801, n11120, n11122, n8250, n8186, n6669, n8020, n11121, 
		n7708, n4800, n11123, n11125, n11124, n11037, n4799, n11128, n4798, n11130, 
		n7418, n11129, n7416, n8194, n11131, n7419, n9575, n9579, n9577, n9375, 
		n4797, n11133, n7626, n11134, n8680, n9077, n11132, n7625, n9083, n7633, 
		n9084, n7628, n4796, n11135, n11137, n8251, n8099, n11136, n11006, n4795, 
		n11139, n11138, n8854, n8853, n4794, n11140, n8180, n11141, n8572, n6616, 
		n9208, n7222, n7723, n4793, n11143, n11145, n9087, n7450, n9800, n11144, 
		n4792, n11146, n7166, n4791, n4790, n11150, n8240, n6771, n11149, n7586, 
		n11148, n11151, n11152, n7840, n7921, n7814, n9107, n9075, n9741, n7584, 
		n4789, n8484, n8830, n4788, n11153, n7132, n11154, n6957, n9884, n6952, 
		n6988, n6959, n4787, n11155, n11157, n7306, n7490, n7742, n7596, n7303, 
		n11158, n9752, n9757, n11159, n6910, n11156, n9095, n4786, n4785, n9889, 
		n7465, n7464, n4784, n11161, n11163, n11162, n10013, n4783, n11166, n7072, 
		n8941, n9885, n6483, n9983, n9323, n4782, n11169, n11171, n11173, n8453, 
		n6881, n11177, n11176, n11179, n11178, n11175, n11181, n8469, n11180, n8718, 
		n11172, n11170, n11182, n11184, n11185, n11186, n11183, n4781, n7912, n4780, 
		n11189, n11190, n7468, n11188, n11187, n4779, n11192, n7546, n8285, n6810, 
		n8289, n4778, n9877, n4777, n11193, n10106, n11194, n8048, n7237, n8268, 
		n11195, n8868, n7235, n7236, n8047, n8213, n8514, n11126, n11036, n10078, 
		n9630, n9626, n11164, n10015, n10014, n8270, n9654, n11196, n11198, n11197, 
		n8886, n9069, n7941, n11200, n10121, n10103, n10105, n9826, n10077, n8869, 
		n4776, n11201, n10964, n8131, n8167, n9322, n9512, n8166, n4775, n11202, 
		n9985, n11203, n7011, n8950, n4774, n11204, n9093, n8885, n7956, n9241, 
		n9243, n4773, n11205, n11207, n6906, n8688, n11206, n8334, n7230, n4772, 
		n11208, n11210, n10020, n9406, n9086, n6407, n6911, n9407, n7021, n11212, 
		n9402, n11211, n11213, n8093, n8151, n11209, n4771, n4770, n8846, n6751, 
		n6750, n7445, n4769, n11215, n11217, n7178, n8995, n6870, n11216, n4768, 
		n11218, n11220, n8949, n7016, n11165, n11219, n10951, n7966, n4767, n9181, 
		n7772, n8890, n7768, n11199, n7114, n4766, n11221, n11223, n8483, n7253, 
		n6426, n7257, n7259, n11222, n4765, n11004, n4764, n8420, n8585, n8418, 
		n6517, n8419, n7833, n9813, n11225, n7834, n4763, n11226, n7802, n8926, 
		n8925, n7064, n11227, n8495, n9975, n7526, n9974, n8501, n7884, n8088, 
		n8085, n7279, n8974, n6486, n9810, n11228, n6610, n8502, n9811, n11231, 
		n11229, n8128, n4762, n11232, n11234, n8593, n8964, n7886, n9356, n7887, 
		n6430, n11236, n9352, n9831, n9830, n9593, n11235, n11032, n11238, n11237, 
		n9378, n6966, n11233, n7218, n4761, n11240, n7535, n11239, n7134, n6917, 
		n9648, n9902, n9424, n9316, n6637, n11241, n4760, n9548, n4759, n11243, 
		n11244, n11242, n4758, n11246, n11248, n7938, n7934, n4757, n11252, n11255, 
		n7152, n11254, n11253, n4756, n11005, n11256, n8600, n6975, n4755, n4754, 
		n11259, n6703, n11261, n11264, n11263, n11267, n11266, n11265, n11262, n11273, 
		n11272, n11271, n11260, n11275, n11278, n11280, n8626, n11277, n7957, n7174, 
		n11276, n9501, n8615, n11268, n11274, n11287, n8628, n11269, n11288, n8625, 
		n8361, n11286, n8875, n9785, n11285, n8135, n6785, n11270, n6700, n6701, 
		n11258, n4753, n4752, n11291, n11290, n8196, n10945, n11292, n8523, n9578, 
		n6819, n9195, n6524, n6526, n6523, n7379, n4751, n8784, n4750, n4749, 
		n11096, n4748, n9151, n4747, n4746, n4745, n4744, n4743, n4742, n10044, 
		n4741, n4740, n4739, n4738, n7693, n4737, n9695, n4736, n4735, n4734, 
		n4733, n4732, n4731, n11279, n4730, n9865, n4729, n4728, n4727, n4726, 
		n4725, n4724, n4723, n4722, n4721, n4720, n4719, n4718, n4717, n11306, 
		n11224, n11307, n11309, n11300, n11298, n11297, n11308, n6536, n11302, n11305, 
		n4716, n11312, n4715, n4714, n9046, n4713, n4712, n4711, n4710, n7327, 
		n4709, n8745, n4708, n4707, n11245, n4706, n9618, n4705, n4704, n4703, 
		n4702, n4701, n4700, n47, n4699, n6566, n4698, n4697, n9600, n4696, 
		n9805, n4695, n4694, n4693, n6978, n8598, n11127, n6979, n4692, n11317, 
		n11316, n4691, n11319, n11321, n6879, n11322, n11320, n9569, n8714, n4690, 
		n4689, n11326, n11325, n4688, n11310, n4687, n11329, n11328, n11103, n11109, 
		n4686, n11333, n11332, n9700, n9408, n4685, n11337, n11336, n11295, n9157, 
		n4684, n11341, n11340, n8789, n8794, n4683, n8921, n4682, n11345, n11344, 
		n11293, n10051, n4681, n11313, n6508, n11348, n7871, n7999, n11349, n4680, 
		n9510, n4679, n4678, n11351, n11350, n11284, n11289, n4677, n11355, n11354, 
		n11294, n7701, n4676, n11359, n11358, n9871, n9878, n4675, n11362, n11363, 
		n7425, n9947, n9553, n7554, n7737, n7736, n4674, n4673, n4672, n11365, 
		n11366, n6828, n9524, n6823, n6715, n8973, n4671, n4670, n4669, n7696, 
		n4668, n9868, n4667, n10048, n4666, n9697, n4665, n9155, n4664, n11281, 
		n4663, n11100, n4662, n8786, n4661, n11369, n11370, n8032, n8031, n11368, 
		n4660, n11371, n9584, n9220, n4659, n4658, n4657, n11373, n8326, n7773, 
		n11372, n4656, n11374, n6544, n4655, n11343, n4654, n11342, n4653, n11334, 
		n4652, n11335, n4651, n11352, n4650, n11339, n4649, n11361, n4648, n11353, 
		n4647, n11346, n4646, n11356, n4645, n11330, n4644, n11338, n4643, n11347, 
		n4642, n11360, n4641, n11357, n4640, n11331, n4639, n11375, n7260, n4638, 
		n4637, n7553, n4636, n4635, n4634, n4633, n4632, n4631, n4630, n4629, 
		n4628, n11191, n4627, n7697, n4626, n9698, n4625, n11282, n4624, n8787, 
		n4623, n11101, n4622, n9156, n4621, n9869, n4620, n10049, n4619, n11377, 
		n11378, n9815, n9818, n11327, n7972, n8519, n9780, n11051, n11379, n10126, 
		n4618, n4617, n4616, n8304, n11382, n11383, n11384, n8303, n10091, n11381, 
		n11380, n4615, n4614, n4613, n11388, n4612, n11389, n6760, n11251, n4611, 
		n11386, n11392, n11393, n4610, n11323, n11395, n11174, n7618, n9566, n4609, 
		n4608, n10133, n4607, n4606, n11397, n4605, n11399, n9513, n4604, n11400, 
		n6889, n4603, n11401, n6686, n4602, n11402, n11391, n11250, n11376, n4601, 
		n11403, n6763, n6761, n11398, n11247, n11249, n4600, n46, n11404, n11405, 
		n6409, n7766, n7098, n9962, n4599, n4598, n11406, n11407, n7898, n11318, 
		n6714, n7402, n7787, n9661, n11408, n8975, n4597, n11314, n4596, n11409, 
		n4595, n11410, n4594, n11412, n11414, n11413, n11301, n11415, n11417, n11304, 
		n11296, n11299, n11416, n11160, n11303, n11324, n11411, n4593, n8298, n11419, 
		n8297, n8299, n10098, n8324, n9789, n9723, n7081, n7082, n8323, n4592, 
		n7542, n11420, n7541, n7543, n8179, n9360, n8041, n9417, n8201, n8200, 
		n8175, n4591, n11421, n4590, n11422, n4589, n11423, n4588, n11424, n4587, 
		n11425, n4586, n11427, n11428, n11426, n8452, n4585, n11432, n75, n9534, 
		n11431, n11433, n10024, n4584, n11315, n9990, n4583, n11435, n95, n6586, 
		n11434, n11436, n8508, n4582, n9009, n4581, n11311, n4580, n11418, n4579, 
		n11438, n4578, n11439, n11437, n4577, n11441, n8804, n9264, n11442, n8825, 
		n9536, n4576, n11443, n7412, n4575, n4574, n11444, n7968, n11445, n11440, 
		n9291, n7413, n9288, n11446, n8976, n7911, n4573, n9054, n11449, n11450, 
		n11451, n9053, n7533, n11448, n9425, n8630, n8223, n11447, n11385, n11452, 
		n8224, n11142, n8225, n4572, n11430, n11454, n11453, n4571, n9268, n4570, 
		n11458, n11457, n11459, n6685, n11390, n11456, n11455, n4569, n4568, n4567, 
		n11460, n8769, n9925, n8788, n4566, n11461, n7167, n11147, n11102, n4565, 
		n11463, n9135, n9586, n11462, n4564, n11464, n6505, n6922, n11283, n4563, 
		n11466, n7377, n7378, n11465, n4562, n11467, n9165, n9166, n9870, n4561, 
		n11469, n9842, n9843, n11468, n4560, n11470, n7474, n8838, n9699, n4559, 
		n11471, n11473, n8473, n11472, n11060, n11061, n7340, n8341, n6882, n6458, 
		n7334, n39, n11474, n11476, n11477, n11478, n8105, n11479, n8353, n11481, 
		n11482, n7241, n11484, n9911, n8231, n11483, n11486, n11487, n11028, n11480, 
		n11475, n10068, n10973, n37, n11488, n11490, n11491, n11492, n8507, n11493, 
		n9366, n11495, n11496, n8220, n11498, n8351, n8399, n11497, n11500, n11501, 
		n10009, n9839, n11494, n11489, n11503, n10955, n8760, n36, n8852, n8851, 
		n7341, n8342, n11429, n6684, n9390, n9969, n22, n21, n6414, n6390, 
		n6457, n8812, n6420, n11505, n9450, n11507, n11509, n11511, n11510, n11508, 
		n11513, n11512, n11506, n8509, n11516, n11519, n8111, n11515, n11525, n6820, 
		n6804, n11524, n11531, n11533, n11530, n11529, n11528, n7124, n11546, n11547, 
		n6728, n11545, n11551, n6974, n10136, n11549, n11555, n11554, n11257, n11553, 
		n11552, n9571, n11558, n11560, n11559, n7076, n8070, n11518, n11557, n10008, 
		n11556, n11563, n11567, n11566, n11565, n11564, n9905, n11562, n9125, n11572, 
		n11575, n9248, n8588, n11571, n11570, n11576, n11580, n11568, n11579, n11540, 
		n11578, n11541, n11577, n11542, n11544, n11387, n11587, n11589, n8332, n11590, 
		n11592, n11593, n11536, n6659, n8539, n11591, n11595, n11539, n11537, n11543, 
		n7109, n8367, n11586, n11599, n9431, n11020, n11561, n11396, n11605, n11606, 
		n8333, n7264, n11604, n11588, n11603, n11608, n11612, n8537, n8986, n11611, 
		n8510, n11610, n8372, n7588, n11609, n9218, n11616, n11617, n11521, n11618, 
		n7777, n11548, n11550, n11615, n11622, n11623, n11626, n7993, n11625, n11581, 
		n8043, n11597, n11214, n11535, n11624, n11634, n11532, n11614, n11534, n11538, 
		n8586, n11633, n6803, n11621, n8965, n11638, n11639, n11522, n11517, n11600, 
		n11602, n7394, n11569, n8693, n11637, n8619, n11643, n11647, n9607, n7593, 
		n11646, n11596, n11598, n11628, n11649, n11645, n7296, n11582, n9897, n11583, 
		n11644, n8209, n11594, n7041, n11642, n11573, n11527, n11620, n7455, n11636, 
		n11601, n11574, n11520, n11641, n6799, n10102, n11526, n11619, n11607, n11523, 
		n11514, n11654, n11653, n11613, n11629, n11635, n11584, n11585, n11650, n11630, 
		n11627, n11632, n11640, n11648, n11652, n11631, n11651, n11168, n8489, n11656, 
		n11657, n8829, n8635, n6880, n11660, n11661, n8536, n11662, n7687, n6607, 
		n7198, n11659, n11664, n11665, n9145, n9910, n9213, n9389, n8396, n10145, 
		n10109, n7049, n9373, n8903, n8408, n9876, n8262, n11663, n7338, n9064, 
		n6833, n11108, n7300, n11673, n11677, n7895, n11676, n6573, n11675, n7449, 
		n11674, n7038, n11672, n7599, n6562, n8014, n9008, n11671, n7089, n8089, 
		n11670, n7430, n8881, n11668, n8884, n7891, n11679, n9091, n11667, n9307, 
		n7034, n8092, n11680, n11678, n11655, n11681, n7414, n11682, n8960, n8525, 
		n11658, n11683, n11064, n8490, n11684, n11685, n10974, n7825, n8106, n7549, 
		n7822, n7826, n8528, n8532, n11485, n9068, n8173, n6840, n6842, n8400, 
		n9454, n11499, n11666, n7612, n11686, n11688, n11687, n9365, n8989, n6596, 
		n9517, n11694, n7090, n7087, n6741, n9076, n9074, n8238, n11693, n9276, 
		n7627, n9042, n9428, n7926, n7832, n11692, n7955, n7359, n7793, n10063, 
		n11691, n8316, n6850, n7100, n7223, n7219, n7722, n11690, n7579, n9339, 
		n7724, n9043, n11689, n9598, n10090, n9315, n6743, n11696, n6397, n7835, 
		n11695, n11697, n11699, n11698, n6391, n6422, n11700, n11701, n9913, n9708, 
		n8229, n8226, n9387, n7238, n11394, n11669, n9718, n11703, n6690, n7353, 
		n7407, n8385, n6674, n7186, n11704, n9017, n6663, n6482, n7071, n6653, 
		n7010, n7875, n6994, n11702, n8817, n6427, n6888, n8185, n9119, n11705, 
		n9116, n6864, n7248, n8069, n7228, n9478, n9282, n8169, n9287, n11167, 
		n9719, n11707, n11706, n11504, n11708, n11230, n9442, n11709, n11710, n11119, 
		n9837, n8217, n8348, n8345, n11711, n9645, n11712, n9726, n9903, n9730, 
		n6633, n9740, n7537, n6913, n9775, n8365, n7570, n8614, n11716, n6556, 
		n6496, n9479, n11715, n8661, n7404, n11714, n10081, n8343, n6748, n11713, 
		n8204, n6749, n10975, n6937, n6707, n7305, n11718, n11720, n11719, n11722, 
		n11725, n11717, n8540, n8541, n6472, n10980, n8542, n11721, n11724, n11723, 
		n8622, n11726, n9838, n11727, n6592, n11502, n9481, n9362, n6822, n8153, 
		n11364, n8103, n8113, n10060, n11367, n7277, n11728, n11729, n11733, n11737, 
		n11738, n11735, n11734, n9928, n6873, n9927, n11731, n11736, n11745, n9392, 
		n11746, n8033, n11732, n7179, n11730, n11743, n11740, n11742, n11741, n6934, 
		n11747, n11739, n11744, n11748, n11029, n11749, n7732, n6404, n6552, n6406, 
		n8663, n11751, n11750, n8664, n11752, n11754, n11753, n7298, n11756, n11755, 
		n7299, n11758, n11757, n9550, n9551, n10981, n11759, n8627, troj0_0_counter_0_, troj0_0_counter_1_, 
		troj0_0_counter_2_, troj0_0_n1, troj0_0_n2, troj0_0_n3, troj0_0_n4, troj0_0_n5, troj0_0_N7, troj0_0_N5, troj0_0_N4, troj0_0_n6, 
		troj0_0_N3, troj0_0_N2, Trojan_out_0_0, Trigger_en_0_0, tempn5237;

	dfxbp_1 DFF_1088_Q_reg( .D(n5549), .CLK(CLK), .Q(n11944) );
	dfxtp_1 DFF_1067_Q_reg( .D(n5536), .CLK(CLK), .Q(n10166) );
	dfxtp_1 DFF_657_Q_reg( .D(n5236), .CLK(CLK), .Q(n10890) );
	dfxtp_1 DFF_507_Q_reg( .D(n5139), .CLK(CLK), .Q(n10167) );
	dfxtp_1 DFF_498_Q_reg( .D(n5132), .CLK(CLK), .Q(n10886) );
	dfxtp_1 DFF_196_Q_reg( .D(n4909), .CLK(CLK), .Q(n10884) );
	dfxtp_1 DFF_190_Q_reg( .D(n4904), .CLK(CLK), .Q(n10885) );
	dfxtp_1 DFF_144_Q_reg( .D(n4872), .CLK(CLK), .Q(n10888) );
	dfxtp_1 DFF_80_Q_reg( .D(n4826), .CLK(CLK), .Q(n10883) );
	dfxtp_1 DFF_75_Q_reg( .D(n4822), .CLK(CLK), .Q(n10889) );
	dfxbp_1 DFF_1387_Q_reg( .D(n5772), .CLK(CLK), .Q(n11781), .Q_N(n6079) );
	dfxtp_1 DFF_64_Q_reg( .D(n4811), .CLK(CLK), .Q(n10887) );
	dfxbp_1 DFF_753_Q_reg( .D(n5306), .CLK(CLK), .Q_N(n5958) );
	dfxbp_1 DFF_685_Q_reg( .D(n5254), .CLK(CLK), .Q(n11974), .Q_N(n6068) );
	dfxbp_1 DFF_1187_Q_reg( .D(n5622), .CLK(CLK), .Q_N(n6031) );
	dfxbp_1 DFF_1083_Q_reg( .D(n5545), .CLK(CLK), .Q_N(n5952) );
	dfxbp_1 DFF_116_Q_reg( .D(n4854), .CLK(CLK), .Q(n11895), .Q_N(n5960) );
	dfxbp_1 DFF_282_Q_reg( .D(n4976), .CLK(CLK), .Q(n11876) );
	dfxbp_1 DFF_1230_Q_reg( .D(n5657), .CLK(CLK), .Q(n11945), .Q_N(n5953) );
	dfxbp_1 DFF_689_Q_reg( .D(n5257), .CLK(CLK), .Q_N(n6032) );
	dfxbp_1 DFF_428_Q_reg( .D(n5081), .CLK(CLK), .Q(n11963), .Q_N(n5882) );
	dfxtp_1 DFF_1191_Q_reg( .D(n5625), .CLK(CLK), .Q(n10601) );
	dfxtp_1 DFF_1176_Q_reg( .D(n5613), .CLK(CLK), .Q(n10600) );
	dfxtp_1 DFF_532_Q_reg( .D(n5153), .CLK(CLK), .Q(n10210) );
	dfxbp_1 DFF_1014_Q_reg( .D(n5495), .CLK(CLK), .Q(n11799) );
	dfxtp_1 DFF_294_Q_reg( .D(n4987), .CLK(CLK), .Q(n10603) );
	dfxtp_1 DFF_654_Q_reg( .D(n4759), .CLK(CLK), .Q(g20763) );
	dfxbp_1 DFF_96_Q_reg( .D(n4839), .CLK(CLK), .Q(n11955) );
	dfxbp_1 DFF_509_Q_reg( .D(n5141), .CLK(CLK), .Q(n11892) );
	dfxbp_1 DFF_349_Q_reg( .D(n5027), .CLK(CLK), .Q(n11859) );
	dfxbp_1 DFF_1245_Q_reg( .D(n5669), .CLK(CLK), .Q(n11775), .Q_N(n5955) );
	dfxbp_1 DFF_1125_Q_reg( .D(n5573), .CLK(CLK), .Q_N(n5872) );
	dfxbp_1 DFF_1178_Q_reg( .D(n5615), .CLK(CLK), .Q(n11936), .Q_N(n6066) );
	dfxtp_1 DFF_1301_Q_reg( .D(n4760), .CLK(CLK), .Q(g20652) );
	dfxbp_1 DFF_958_Q_reg( .D(n5456), .CLK(CLK), .Q(n11907), .Q_N(n5899) );
	dfxtp_1 DFF_1396_Q_reg( .D(n5779), .CLK(CLK), .Q(n10611) );
	dfxbp_1 DFF_1304_Q_reg( .D(n5712), .CLK(CLK), .Q(n11943), .Q_N(n5903) );
	dfxtp_1 DFF_458_Q_reg( .D(n5106), .CLK(CLK), .Q(n10614) );
	dfxbp_1 DFF_723_Q_reg( .D(n5282), .CLK(CLK), .Q(n11956), .Q_N(n5902) );
	dfxtp_1 DFF_235_Q_reg( .D(n4937), .CLK(CLK), .Q(n10608) );
	dfxbp_1 DFF_653_Q_reg( .D(n5234), .CLK(CLK), .Q(n11972), .Q_N(n5900) );
	dfxtp_1 DFF_377_Q_reg( .D(n5045), .CLK(CLK), .Q(n10606) );
	dfxbp_1 DFF_304_Q_reg( .D(n4996), .CLK(CLK), .Q(n11839) );
	dfxtp_1 DFF_166_Q_reg( .D(n4887), .CLK(CLK), .Q(n10619) );
	dfxbp_1 DFF_584_Q_reg( .D(n5188), .CLK(CLK), .Q(n11942), .Q_N(n5898) );
	dfxtp_1 DFF_603_Q_reg( .D(n5201), .CLK(CLK), .Q(n10604) );
	dfxbp_1 DFF_776_Q_reg( .D(n5322), .CLK(CLK), .Q(n11968), .Q_N(n5901) );
	dfxtp_1 DFF_299_Q_reg( .D(n4991), .CLK(CLK), .Q(n10615) );
	dfxbp_1 DFF_27_Q_reg( .D(n4783), .CLK(CLK), .Q(n11960), .Q_N(n5904) );
	dfxtp_1 DFF_810_Q_reg( .D(n5347), .CLK(CLK), .Q(n10617) );
	dfxtp_1 DFF_1352_Q_reg( .D(n4750), .CLK(CLK), .Q(g13049) );
	dfxtp_1 DFF_695_Q_reg( .D(n4735), .CLK(CLK), .Q(g17813) );
	dfxtp_1 DFF_783_Q_reg( .D(n4738), .CLK(CLK), .Q(g17678) );
	dfxtp_1 DFF_666_Q_reg( .D(n5241), .CLK(CLK), .Q(n10224) );
	dfxtp_1 DFF_163_Q_reg( .D(n4729), .CLK(CLK), .Q(g13099) );
	dfxtp_1 DFF_971_Q_reg( .D(n4744), .CLK(CLK), .Q(g17871) );
	dfxtp_1 DFF_780_Q_reg( .D(n4737), .CLK(CLK), .Q(g17764) );
	dfxtp_1 DFF_1023_Q_reg( .D(n5501), .CLK(CLK), .Q(n10221) );
	dfxtp_1 DFF_616_Q_reg( .D(n4733), .CLK(CLK), .Q(g13039) );
	dfxtp_1 DFF_765_Q_reg( .D(n4736), .CLK(CLK), .Q(g17787) );
	dfxtp_1 DFF_360_Q_reg( .D(n4731), .CLK(CLK), .Q(g17639) );
	dfxtp_1 DFF_281_Q_reg( .D(n4975), .CLK(CLK), .Q(n10225) );
	dfxtp_1 DFF_1155_Q_reg( .D(n4747), .CLK(CLK), .Q(g14421) );
	dfxtp_1 DFF_856_Q_reg( .D(n4740), .CLK(CLK), .Q(g16874) );
	dfxtp_1 DFF_1359_Q_reg( .D(n4751), .CLK(CLK), .Q(g16686) );
	dfxtp_1 DFF_1303_Q_reg( .D(n5711), .CLK(CLK), .Q(n10228) );
	dfxtp_1 DFF_34_Q_reg( .D(n4728), .CLK(CLK), .Q(g14451) );
	dfxtp_1 DFF_873_Q_reg( .D(n4741), .CLK(CLK), .Q(g16924) );
	dfxtp_1 DFF_1300_Q_reg( .D(n4749), .CLK(CLK), .Q(g16722) );
	dfxtp_1 DFF_290_Q_reg( .D(n4983), .CLK(CLK), .Q(n10227) );
	dfxtp_1 DFF_642_Q_reg( .D(n4734), .CLK(CLK), .Q(g14518) );
	dfxtp_1 DFF_367_Q_reg( .D(n4732), .CLK(CLK), .Q(g16955) );
	dfxtp_1 DFF_1219_Q_reg( .D(n4748), .CLK(CLK), .Q(g16748) );
	dfxtp_1 DFF_995_Q_reg( .D(n5482), .CLK(CLK), .Q(n10226) );
	dfxtp_1 DFF_1087_Q_reg( .D(n4745), .CLK(CLK), .Q(g13068) );
	dfxtp_1 DFF_848_Q_reg( .D(n4739), .CLK(CLK), .Q(g17819) );
	dfxtp_1 DFF_279_Q_reg( .D(n4730), .CLK(CLK), .Q(g17715) );
	dfxtp_1 DFF_22_Q_reg( .D(n4778), .CLK(CLK), .Q(n10223) );
	dfxtp_1 DFF_1119_Q_reg( .D(n4746), .CLK(CLK), .Q(g13085) );
	dfxtp_1 DFF_970_Q_reg( .D(n4743), .CLK(CLK), .Q(g17845) );
	dfxtp_1 DFF_898_Q_reg( .D(n4742), .CLK(CLK), .Q(g17743) );
	dfxtp_1 DFF_53_Q_reg( .D(n4803), .CLK(CLK), .Q(n10222) );
	dfxtp_1 DFF_709_Q_reg( .D(n4597), .CLK(CLK), .Q(g341) );
	dfxbp_1 DFF_1003_Q_reg( .D(n5486), .CLK(CLK), .Q(n11937), .Q_N(n6092) );
	dfxtp_1 DFF_652_Q_reg( .D(n5233), .CLK(CLK), .Q(n10881) );
	dfxbp_1 DFF_10_Q_reg( .D(n4767), .CLK(CLK), .Q_N(n5919) );
	dfxbp_1 DFF_525_Q_reg( .D(n5150), .CLK(CLK), .Q(n11913), .Q_N(n5905) );
	dfxbp_1 DFF_278_Q_reg( .D(n4973), .CLK(CLK), .Q(n11912), .Q_N(n5887) );
	dfxbp_1 DFF_113_Q_reg( .D(n4852), .CLK(CLK), .Q(n11940), .Q_N(n5948) );
	dfxtp_1 DFF_292_Q_reg( .D(n4985), .CLK(CLK), .Q(n10170) );
	dfxtp_1 DFF_1042_Q_reg( .D(n5517), .CLK(CLK), .Q(n10449) );
	dfxtp_1 DFF_238_Q_reg( .D(n4940), .CLK(CLK), .Q(n10205) );
	dfxbp_1 DFF_1126_Q_reg( .D(n5574), .CLK(CLK), .Q(n11789), .Q_N(n5950) );
	dfxbp_1 DFF_1365_Q_reg( .D(n5754), .CLK(CLK), .Q(n11966), .Q_N(n5954) );
	dfxbp_1 DFF_900_Q_reg( .D(n5412), .CLK(CLK), .Q(n11938), .Q_N(n6072) );
	dfxtp_1 DFF_866_Q_reg( .D(n5385), .CLK(CLK), .Q(n10501) );
	dfxbp_1 DFF_252_Q_reg( .D(n4953), .CLK(CLK), .Q(n11843), .Q_N(n6080) );
	dfxtp_1 DFF_988_Q_reg( .D(n5477), .CLK(CLK), .Q(n10877) );
	dfxtp_1 DFF_902_Q_reg( .D(n5414), .CLK(CLK), .Q(n10357) );
	dfxbp_1 DFF_510_Q_reg( .D(n5142), .CLK(CLK), .Q(n11761), .Q_N(n6085) );
	dfxtp_1 DFF_544_Q_reg( .D(n5162), .CLK(CLK), .Q(n10428) );
	dfxbp_1 DFF_324_Q_reg( .D(n5012), .CLK(CLK), .Q(n11763), .Q_N(n6084) );
	dfxtp_1 DFF_972_Q_reg( .D(n5465), .CLK(CLK), .Q(n10882) );
	dfxtp_1 DFF_357_Q_reg( .D(n4758), .CLK(CLK), .Q(g20901) );
	dfxtp_1 DFF_143_Q_reg( .D(n4602), .CLK(CLK), .Q(g496) );
	dfxtp_1 DFF_752_Q_reg( .D(n47), .CLK(CLK), .Q(g12368) );
	dfxtp_1 DFF_7_Q_reg( .D(n4765), .CLK(CLK), .Q(n10662) );
	dfxbp_1 DFF_88_Q_reg( .D(n4831), .CLK(CLK), .Q(n11857), .Q_N(n5888) );
	dfxtp_1 DFF_515_Q_reg( .D(n4584), .CLK(CLK), .Q(g12184) );
	dfxtp_1 DFF_256_Q_reg( .D(n4957), .CLK(CLK), .Q(n10664) );
	dfxbp_1 DFF_876_Q_reg( .D(n5392), .CLK(CLK), .Q(n11858), .Q_N(n6082) );
	dfxbp_1 DFF_745_Q_reg( .D(n5299), .CLK(CLK), .Q(n11819), .Q_N(n6053) );
	dfxbp_1 DFF_1060_Q_reg( .D(n5530), .CLK(CLK), .Q(n11954), .Q_N(n6088) );
	dfxbp_1 DFF_555_Q_reg( .D(n5168), .CLK(CLK), .Q_N(n5914) );
	dfxtp_1 DFF_258_Q_reg( .D(n4959), .CLK(CLK), .Q(n10663) );
	dfxtp_1 DFF_612_Q_reg( .D(n4582), .CLK(CLK), .Q(g8291) );
	dfxbp_1 DFF_842_Q_reg( .D(n5366), .CLK(CLK), .Q_N(n5920) );
	dfxbp_1 DFF_597_Q_reg( .D(n5197), .CLK(CLK), .Q(n11826), .Q_N(n6070) );
	dfxtp_1 DFF_715_Q_reg( .D(n5274), .CLK(CLK), .Q(n10234) );
	dfxtp_1 DFF_1308_Q_reg( .D(n88), .CLK(CLK), .Q(g8416) );
	dfxbp_1 DFF_421_Q_reg( .D(n5077), .CLK(CLK), .Q(n11834), .Q_N(n5970) );
	dfxbp_1 DFF_131_Q_reg( .D(n4864), .CLK(CLK), .Q(n11914), .Q_N(n5907) );
	dfxbp_1 DFF_1144_Q_reg( .D(n5590), .CLK(CLK), .Q(n11939), .Q_N(n6062) );
	dfxtp_1 DFF_880_Q_reg( .D(n85), .CLK(CLK), .Q(n10450) );
	dfxtp_1 DFF_185_Q_reg( .D(n4583), .CLK(CLK), .Q(g10500) );
	dfxbp_1 DFF_791_Q_reg( .D(n5333), .CLK(CLK), .Q_N(n5944) );
	dfxbp_1 DFF_24_Q_reg( .D(n4780), .CLK(CLK), .Q_N(n19679) );
	dfxbp_1 DFF_936_Q_reg( .D(n5439), .CLK(CLK), .Q(n11807), .Q_N(n6069) );
	dfxtp_1 DFF_758_Q_reg( .D(n4593), .CLK(CLK), .Q(g933) );
	dfxbp_1 DFF_563_Q_reg( .D(n5802), .CLK(CLK), .Q(n11957), .Q_N(n5884) );
	dfxbp_1 DFF_580_Q_reg( .D(n5184), .CLK(CLK), .Q(n11828), .Q_N(n5932) );
	dfxtp_1 DFF_127_Q_reg( .D(n4860), .CLK(CLK), .Q(n10455) );
	dfxtp_1 DFF_334_Q_reg( .D(n61), .CLK(CLK), .Q(g8475) );
	dfxtp_1 DFF_1072_Q_reg( .D(n4585), .CLK(CLK), .Q(g10527) );
	dfxbp_1 DFF_171_Q_reg( .D(n4891), .CLK(CLK), .Q_N(n5945) );
	dfxbp_1 DFF_577_Q_reg( .D(n5182), .CLK(CLK), .Q(n11829), .Q_N(n5934) );
	dfxbp_1 DFF_1419_Q_reg( .D(n5797), .CLK(CLK), .Q(n11959), .Q_N(n5908) );
	dfxbp_1 DFF_211_Q_reg( .D(n4919), .CLK(CLK), .Q(n11891), .Q_N(n6033) );
	dfxbp_1 DFF_740_Q_reg( .D(n5296), .CLK(CLK), .Q(n11861) );
	dfxbp_1 DFF_1092_Q_reg( .D(n5553), .CLK(CLK), .Q_N(n19677) );
	dfxbp_1 DFF_1189_Q_reg( .D(n5624), .CLK(CLK), .Q(n11788), .Q_N(n5961) );
	dfxtp_1 DFF_754_Q_reg( .D(n4592), .CLK(CLK), .Q(g1277) );
	dfxtp_1 DFF_323_Q_reg( .D(n5011), .CLK(CLK), .Q(n10454) );
	dfxbp_1 DFF_822_Q_reg( .D(n5355), .CLK(CLK), .Q(n11816), .Q_N(n5933) );
	dfxbp_1 DFF_594_Q_reg( .D(n5195), .CLK(CLK), .Q(n11862), .Q_N(n5881) );
	dfxbp_1 DFF_1089_Q_reg( .D(n5550), .CLK(CLK), .Q(n11866), .Q_N(n6074) );
	dfxbp_1 DFF_943_Q_reg( .D(n5442), .CLK(CLK), .Q(n11864), .Q_N(n5866) );
	dfxbp_1 DFF_658_Q_reg( .D(n5237), .CLK(CLK), .Q(n11865), .Q_N(n5969) );
	dfxbp_1 DFF_567_Q_reg( .D(n5174), .CLK(CLK), .Q(n11867), .Q_N(n6076) );
	dfxbp_1 DFF_472_Q_reg( .D(n5116), .CLK(CLK), .Q(n11869), .Q_N(n6077) );
	dfxbp_1 DFF_1254_Q_reg( .D(n5675), .CLK(CLK), .Q(n11863), .Q_N(n5871) );
	dfxbp_1 DFF_1009_Q_reg( .D(n5491), .CLK(CLK), .Q(n11868), .Q_N(n6075) );
	dfxtp_1 DFF_739_Q_reg( .D(n4575), .CLK(CLK), .Q(g10122) );
	dfxtp_1 DFF_325_Q_reg( .D(n5013), .CLK(CLK), .Q(n10665) );
	dfxtp_1 DFF_1417_Q_reg( .D(n5795), .CLK(CLK), .Q(n10453) );
	dfxbp_1 DFF_320_Q_reg( .D(n5008), .CLK(CLK), .Q(n11897), .Q_N(n6064) );
	dfxtp_1 DFF_1384_Q_reg( .D(n5770), .CLK(CLK), .Q(n10666) );
	dfxbp_1 DFF_1043_Q_reg( .D(n5518), .CLK(CLK), .Q(n11964) );
	dfxtp_1 DFF_858_Q_reg( .D(n5378), .CLK(CLK), .Q(n10211) );
	dfxtp_1 DFF_1049_Q_reg( .D(n4581), .CLK(CLK), .Q(g8788) );
	dfxbp_1 DFF_773_Q_reg( .D(n5320), .CLK(CLK), .Q_N(n5940) );
	dfxbp_1 DFF_51_Q_reg( .D(n4801), .CLK(CLK), .Q_N(n5938) );
	dfxbp_1 DFF_476_Q_reg( .D(n5118), .CLK(CLK), .Q(n11952), .Q_N(n6014) );
	dfxbp_1 DFF_71_Q_reg( .D(n4818), .CLK(CLK), .Q(n11951), .Q_N(n6016) );
	dfxbp_1 DFF_257_Q_reg( .D(n4958), .CLK(CLK), .Q_N(n5923) );
	dfxbp_1 DFF_633_Q_reg( .D(n5219), .CLK(CLK), .Q_N(n5930) );
	dfxbp_1 DFF_192_Q_reg( .D(n4905), .CLK(CLK), .Q_N(n5926) );
	dfxbp_1 DFF_1355_Q_reg( .D(n5746), .CLK(CLK), .Q_N(n5925) );
	dfxbp_1 DFF_370_Q_reg( .D(n5041), .CLK(CLK), .Q_N(n5935) );
	dfxbp_1 DFF_419_Q_reg( .D(n5076), .CLK(CLK), .Q_N(n5936) );
	dfxbp_1 DFF_1166_Q_reg( .D(n5605), .CLK(CLK), .Q(n11900), .Q_N(n6006) );
	dfxbp_1 DFF_225_Q_reg( .D(n4930), .CLK(CLK), .Q(n11899), .Q_N(n5987) );
	dfxbp_1 DFF_134_Q_reg( .D(n4866), .CLK(CLK), .Q_N(n5937) );
	dfxbp_1 DFF_640_Q_reg( .D(n5224), .CLK(CLK), .Q(n11823), .Q_N(n6018) );
	dfxbp_1 DFF_9_Q_reg( .D(n4766), .CLK(CLK), .Q(n11856), .Q_N(n6019) );
	dfxtp_1 DFF_1210_Q_reg( .D(n5642), .CLK(CLK), .Q(n10500) );
	dfxbp_1 DFF_1128_Q_reg( .D(n5576), .CLK(CLK), .Q(n11874), .Q_N(n5976) );
	dfxbp_1 DFF_868_Q_reg( .D(n5387), .CLK(CLK), .Q(n11873), .Q_N(n5977) );
	dfxbp_1 DFF_1160_Q_reg( .D(n5600), .CLK(CLK), .Q_N(n5921) );
	dfxbp_1 DFF_917_Q_reg( .D(n5423), .CLK(CLK), .Q(n11811), .Q_N(n5973) );
	dfxbp_1 DFF_108_Q_reg( .D(n4849), .CLK(CLK), .Q(n11875), .Q_N(n6010) );
	dfxbp_1 DFF_105_Q_reg( .D(n4846), .CLK(CLK), .Q(n11850), .Q_N(n6011) );
	dfxbp_1 DFF_1058_Q_reg( .D(n5529), .CLK(CLK), .Q(n11883), .Q_N(n5979) );
	dfxbp_1 DFF_815_Q_reg( .D(n5352), .CLK(CLK), .Q(n11817), .Q_N(n5980) );
	dfxbp_1 DFF_1085_Q_reg( .D(n5547), .CLK(CLK), .Q_N(n5924) );
	dfxbp_1 DFF_854_Q_reg( .D(n5375), .CLK(CLK), .Q(n11815), .Q_N(n5978) );
	dfxbp_1 DFF_949_Q_reg( .D(n5447), .CLK(CLK), .Q(n11806), .Q_N(n5986) );
	dfxtp_1 DFF_336_Q_reg( .D(n5017), .CLK(CLK), .Q(n10495) );
	dfxbp_1 DFF_1052_Q_reg( .D(n5524), .CLK(CLK), .Q_N(n5929) );
	dfxbp_1 DFF_730_Q_reg( .D(n5288), .CLK(CLK), .Q(n11871), .Q_N(n6002) );
	dfxbp_1 DFF_345_Q_reg( .D(n5024), .CLK(CLK), .Q(n11870), .Q_N(n6003) );
	dfxbp_1 DFF_1120_Q_reg( .D(n5570), .CLK(CLK), .Q_N(n5922) );
	dfxbp_1 DFF_628_Q_reg( .D(n5217), .CLK(CLK), .Q(n11824), .Q_N(n5982) );
	dfxbp_1 DFF_1244_Q_reg( .D(n5668), .CLK(CLK), .Q(n11785), .Q_N(n5971) );
	dfxtp_1 DFF_1177_Q_reg( .D(n5614), .CLK(CLK), .Q(n10499) );
	dfxbp_1 DFF_588_Q_reg( .D(n5190), .CLK(CLK), .Q(n11827), .Q_N(n6004) );
	dfxbp_1 DFF_291_Q_reg( .D(n4984), .CLK(CLK), .Q(n11841), .Q_N(n6005) );
	dfxtp_1 DFF_779_Q_reg( .D(n5325), .CLK(CLK), .Q(n10493) );
	dfxbp_1 DFF_1013_Q_reg( .D(n5494), .CLK(CLK), .Q(n11800), .Q_N(n5985) );
	dfxtp_1 DFF_414_Q_reg( .D(n5074), .CLK(CLK), .Q(n10498) );
	dfxbp_1 DFF_397_Q_reg( .D(n5060), .CLK(CLK), .Q_N(n5927) );
	dfxbp_1 DFF_179_Q_reg( .D(n4897), .CLK(CLK), .Q(n11894), .Q_N(n6008) );
	dfxbp_1 DFF_904_Q_reg( .D(n5416), .CLK(CLK), .Q(n11893), .Q_N(n5974) );
	dfxbp_1 DFF_59_Q_reg( .D(n4807), .CLK(CLK), .Q_N(n5928) );
	dfxbp_1 DFF_483_Q_reg( .D(n5122), .CLK(CLK), .Q(n11833), .Q_N(n6012) );
	dfxbp_1 DFF_82_Q_reg( .D(n4827), .CLK(CLK), .Q(n11851), .Q_N(n6013) );
	dfxtp_1 DFF_298_Q_reg( .D(n4990), .CLK(CLK), .Q(n10494) );
	dfxbp_1 DFF_1186_Q_reg( .D(n5621), .CLK(CLK), .Q(n11903), .Q_N(n5993) );
	dfxbp_1 DFF_950_Q_reg( .D(n5448), .CLK(CLK), .Q(n11902), .Q_N(n5972) );
	dfxbp_1 DFF_1212_Q_reg( .D(n5644), .CLK(CLK), .Q_N(n5939) );
	dfxbp_1 DFF_983_Q_reg( .D(n5472), .CLK(CLK), .Q(n11803), .Q_N(n5992) );
	dfxbp_1 DFF_1095_Q_reg( .D(n5556), .CLK(CLK), .Q(n11793), .Q_N(n5999) );
	dfxtp_1 DFF_497_Q_reg( .D(n5131), .CLK(CLK), .Q(n10497) );
	dfxbp_1 DFF_895_Q_reg( .D(n5408), .CLK(CLK), .Q(n11812), .Q_N(n5994) );
	dfxbp_1 DFF_1297_Q_reg( .D(n5707), .CLK(CLK), .Q(n11783), .Q_N(n6015) );
	dfxtp_1 DFF_55_Q_reg( .D(n4805), .CLK(CLK), .Q(n10496) );
	dfxtp_1 DFF_651_Q_reg( .D(n5232), .CLK(CLK), .Q(n10312) );
	dfxtp_1 DFF_124_Q_reg( .D(n4859), .CLK(CLK), .Q(n10316) );
	dfxtp_1 DFF_926_Q_reg( .D(n5431), .CLK(CLK), .Q(n10313) );
	dfxtp_1 DFF_1055_Q_reg( .D(n5527), .CLK(CLK), .Q(n10309) );
	dfxtp_1 DFF_1134_Q_reg( .D(n5581), .CLK(CLK), .Q(n10315) );
	dfxtp_1 DFF_300_Q_reg( .D(n4992), .CLK(CLK), .Q(n10310) );
	dfxtp_1 DFF_87_Q_reg( .D(n4830), .CLK(CLK), .Q(n10314) );
	dfxtp_1 DFF_14_Q_reg( .D(n4770), .CLK(CLK), .Q(n10311) );
	dfxbp_1 DFF_4_Q_reg( .D(n4763), .CLK(CLK), .Q(n11762), .Q_N(n6030) );
	dfxbp_1 DFF_65_Q_reg( .D(n4812), .CLK(CLK), .Q(n11852), .Q_N(n6025) );
	dfxbp_1 DFF_1247_Q_reg( .D(n5670), .CLK(CLK), .Q(n11784), .Q_N(n5984) );
	dfxbp_1 DFF_625_Q_reg( .D(n5214), .CLK(CLK), .Q(n11825), .Q_N(n6001) );
	dfxtp_1 DFF_457_Q_reg( .D(n5105), .CLK(CLK), .Q(n10488) );
	dfxbp_1 DFF_727_Q_reg( .D(n5285), .CLK(CLK), .Q(n11773), .Q_N(n6027) );
	dfxbp_1 DFF_61_Q_reg( .D(n4808), .CLK(CLK), .Q(n11853), .Q_N(n6026) );
	dfxbp_1 DFF_1097_Q_reg( .D(n5558), .CLK(CLK), .Q(n11792), .Q_N(n5989) );
	dfxbp_1 DFF_1380_Q_reg( .D(n5766), .CLK(CLK), .Q(n11782), .Q_N(n6024) );
	dfxbp_1 DFF_890_Q_reg( .D(n5403), .CLK(CLK), .Q(n11813), .Q_N(n5995) );
	dfxtp_1 DFF_960_Q_reg( .D(n5458), .CLK(CLK), .Q(n10486) );
	dfxbp_1 DFF_1096_Q_reg( .D(n5557), .CLK(CLK), .Q(n11772), .Q_N(n6036) );
	dfxbp_1 DFF_1231_Q_reg( .D(n5658), .CLK(CLK), .Q(n11786), .Q_N(n6021) );
	dfxbp_1 DFF_1030_Q_reg( .D(n5507), .CLK(CLK), .Q(n11796), .Q_N(n5990) );
	dfxbp_1 DFF_204_Q_reg( .D(n4914), .CLK(CLK), .Q(n11846), .Q_N(n6007) );
	dfxtp_1 DFF_1026_Q_reg( .D(n5504), .CLK(CLK), .Q(n10489) );
	dfxbp_1 DFF_273_Q_reg( .D(n4968), .CLK(CLK), .Q(n11764), .Q_N(n6029) );
	dfxbp_1 DFF_930_Q_reg( .D(n5434), .CLK(CLK), .Q(n11808), .Q_N(n5996) );
	dfxbp_1 DFF_887_Q_reg( .D(n5400), .CLK(CLK), .Q(n11814), .Q_N(n5975) );
	dfxbp_1 DFF_1025_Q_reg( .D(n5503), .CLK(CLK), .Q(n11797), .Q_N(n5991) );
	dfxtp_1 DFF_1171_Q_reg( .D(n5608), .CLK(CLK), .Q(n10487) );
	dfxbp_1 DFF_255_Q_reg( .D(n4956), .CLK(CLK), .Q(n11767), .Q_N(n6037) );
	dfxbp_1 DFF_1394_Q_reg( .D(n5777), .CLK(CLK), .Q(n11780), .Q_N(n6023) );
	dfxbp_1 DFF_924_Q_reg( .D(n5429), .CLK(CLK), .Q(n11809), .Q_N(n5981) );
	dfxbp_1 DFF_641_Q_reg( .D(n5225), .CLK(CLK), .Q(n11822), .Q_N(n6000) );
	dfxtp_1 DFF_465_Q_reg( .D(n5111), .CLK(CLK), .Q(n10490) );
	dfxbp_1 DFF_246_Q_reg( .D(n4948), .CLK(CLK), .Q(n11776), .Q_N(n6028) );
	dfxbp_1 DFF_564_Q_reg( .D(n5173), .CLK(CLK), .Q(n11830), .Q_N(n5983) );
	dfxbp_1 DFF_735_Q_reg( .D(n5293), .CLK(CLK), .Q(n11820), .Q_N(n5997) );
	dfxbp_1 DFF_1172_Q_reg( .D(n5609), .CLK(CLK), .Q(n11770), .Q_N(n6034) );
	dfxbp_1 DFF_973_Q_reg( .D(n5466), .CLK(CLK), .Q(n11804), .Q_N(n6022) );
	dfxbp_1 DFF_1422_Q_reg( .D(n5798), .CLK(CLK), .Q(n11778), .Q_N(n5998) );
	dfxbp_1 DFF_968_Q_reg( .D(n5464), .CLK(CLK), .Q(n11805), .Q_N(n6020) );
	dfxtp_1 DFF_2_Q_reg( .D(n4762), .CLK(CLK), .Q(n10491) );
	dfxbp_1 DFF_1258_Q_reg( .D(n5677), .CLK(CLK), .Q(n11771), .Q_N(n6035) );
	dfxbp_1 DFF_41_Q_reg( .D(n4793), .CLK(CLK), .Q(n11854), .Q_N(n6017) );
	dfxbp_1 DFF_16_Q_reg( .D(n4772), .CLK(CLK), .Q(n11855), .Q_N(n5988) );
	dfxbp_1 DFF_173_Q_reg( .D(n4893), .CLK(CLK), .Q(n11848), .Q_N(n6009) );
	dfxtp_1 DFF_306_Q_reg( .D(n4997), .CLK(CLK), .Q(n10492) );
	dfxtp_1 DFF_1033_Q_reg( .D(n4616), .CLK(CLK), .Q(g20654) );
	dfxbp_1 DFF_302_Q_reg( .D(n4994), .CLK(CLK), .Q(n11840), .Q_N(n5886) );
	dfxbp_1 DFF_1331_Q_reg( .D(n5730), .CLK(CLK), .Q(n11901), .Q_N(n5896) );
	dfxbp_1 DFF_379_Q_reg( .D(n5047), .CLK(CLK), .Q(n11962) );
	dfxbp_1 DFF_581_Q_reg( .D(n5185), .CLK(CLK), .Q_N(n5867) );
	dfxtp_1 DFF_1220_Q_reg( .D(n4618), .CLK(CLK), .Q(g111) );
	dfxbp_1 DFF_623_Q_reg( .D(n5213), .CLK(CLK), .Q(n11946), .Q_N(n5894) );
	dfxbp_1 DFF_45_Q_reg( .D(n4797), .CLK(CLK), .Q_N(n5869) );
	dfxbp_1 DFF_1071_Q_reg( .D(n5540), .CLK(CLK), .Q(n11920), .Q_N(n6048) );
	dfxbp_1 DFF_1140_Q_reg( .D(n5587), .CLK(CLK), .Q(n11921) );
	dfxbp_1 DFF_462_Q_reg( .D(n5108), .CLK(CLK), .Q_N(n5873) );
	dfxbp_1 DFF_993_Q_reg( .D(n5480), .CLK(CLK), .Q(n11904), .Q_N(n5890) );
	dfxbp_1 DFF_301_Q_reg( .D(n4993), .CLK(CLK), .Q_N(n5864) );
	dfxbp_1 DFF_841_Q_reg( .D(n5365), .CLK(CLK), .Q(n11926), .Q_N(n6049) );
	dfxbp_1 DFF_1031_Q_reg( .D(n5508), .CLK(CLK), .Q(n11927), .Q_N(n6097) );
	dfxbp_1 DFF_1337_Q_reg( .D(n5733), .CLK(CLK), .Q_N(n5918) );
	dfxbp_1 DFF_387_Q_reg( .D(n5053), .CLK(CLK), .Q(n11877), .Q_N(n5892) );
	dfxbp_1 DFF_928_Q_reg( .D(n5432), .CLK(CLK), .Q_N(n5943) );
	dfxbp_1 DFF_444_Q_reg( .D(n5093), .CLK(CLK), .Q(n11924), .Q_N(n6046) );
	dfxbp_1 DFF_499_Q_reg( .D(n5133), .CLK(CLK), .Q(n11925), .Q_N(n6095) );
	dfxbp_1 DFF_1063_Q_reg( .D(n5532), .CLK(CLK), .Q(n11795), .Q_N(n5965) );
	dfxbp_1 DFF_319_Q_reg( .D(n5007), .CLK(CLK), .Q(n11837), .Q_N(n5885) );
	dfxtp_1 DFF_1111_Q_reg( .D(n4617), .CLK(CLK), .Q(g85) );
	dfxbp_1 DFF_1070_Q_reg( .D(n5539), .CLK(CLK), .Q(n11950), .Q_N(n5893) );
	dfxbp_1 DFF_1093_Q_reg( .D(n5554), .CLK(CLK), .Q(n11794), .Q_N(n5963) );
	dfxbp_1 DFF_964_Q_reg( .D(n5460), .CLK(CLK), .Q_N(n5868) );
	dfxbp_1 DFF_322_Q_reg( .D(n5010), .CLK(CLK), .Q(n11928), .Q_N(n6047) );
	dfxbp_1 DFF_1213_Q_reg( .D(n5645), .CLK(CLK), .Q(n11929), .Q_N(n6093) );
	dfxbp_1 DFF_1064_Q_reg( .D(n5533), .CLK(CLK), .Q(n11953), .Q_N(n5891) );
	dfxbp_1 DFF_342_Q_reg( .D(n5022), .CLK(CLK), .Q(n11836), .Q_N(n5964) );
	dfxbp_1 DFF_552_Q_reg( .D(n5167), .CLK(CLK), .Q(n11958), .Q_N(n5889) );
	dfxbp_1 DFF_153_Q_reg( .D(n4877), .CLK(CLK), .Q(n11849), .Q_N(n5966) );
	dfxbp_1 DFF_583_Q_reg( .D(n5187), .CLK(CLK), .Q_N(n5863) );
	dfxbp_1 DFF_1277_Q_reg( .D(n5692), .CLK(CLK), .Q(n11934), .Q_N(n6052) );
	dfxbp_1 DFF_1418_Q_reg( .D(n5796), .CLK(CLK), .Q(n11935), .Q_N(n6096) );
	dfxbp_1 DFF_865_Q_reg( .D(n5384), .CLK(CLK), .Q_N(g23759) );
	dfxbp_1 DFF_705_Q_reg( .D(n5268), .CLK(CLK), .Q(n11915), .Q_N(n5895) );
	dfxbp_1 DFF_1216_Q_reg( .D(n5648), .CLK(CLK), .Q_N(n5876) );
	dfxbp_1 DFF_1179_Q_reg( .D(n5616), .CLK(CLK), .Q(n11930), .Q_N(n6045) );
	dfxbp_1 DFF_520_Q_reg( .D(n5147), .CLK(CLK), .Q(n11931) );
	dfxbp_1 DFF_1028_Q_reg( .D(n5505), .CLK(CLK), .Q_N(n5862) );
	dfxbp_1 DFF_576_Q_reg( .D(n5181), .CLK(CLK), .Q_N(g23652) );
	dfxbp_1 DFF_818_Q_reg( .D(n5353), .CLK(CLK), .Q_N(n5877) );
	dfxbp_1 DFF_488_Q_reg( .D(n5126), .CLK(CLK), .Q(n11922), .Q_N(n6051) );
	dfxbp_1 DFF_825_Q_reg( .D(n5356), .CLK(CLK), .Q(n11923), .Q_N(n6098) );
	dfxbp_1 DFF_1051_Q_reg( .D(n5523), .CLK(CLK), .Q_N(n5942) );
	dfxtp_1 DFF_364_Q_reg( .D(n5038), .CLK(CLK), .Q(n10451) );
	dfxbp_1 DFF_814_Q_reg( .D(n5351), .CLK(CLK), .Q(n11932), .Q_N(n6050) );
	dfxbp_1 DFF_1163_Q_reg( .D(n5603), .CLK(CLK), .Q(n11933), .Q_N(n6094) );
	dfxtp_1 DFF_1182_Q_reg( .D(n5619), .CLK(CLK), .Q(n10452) );
	dfxtp_1 DFF_944_Q_reg( .D(n4580), .CLK(CLK), .Q(g8919) );
	dfxtp_1 DFF_919_Q_reg( .D(n4594), .CLK(CLK), .Q(g4242) );
	dfxtp_1 DFF_125_Q_reg( .D(n4573), .CLK(CLK), .Q(g21270) );
	dfxbp_1 DFF_224_Q_reg( .D(n4929), .CLK(CLK), .Q_N(n5909) );
	dfxtp_1 DFF_1256_Q_reg( .D(n4595), .CLK(CLK), .Q(g8277) );
	dfxtp_1 DFF_259_Q_reg( .D(n4960), .CLK(CLK), .Q(n10620) );
	dfxtp_1 DFF_1414_Q_reg( .D(n4596), .CLK(CLK), .Q(g8342) );
	dfxtp_1 DFF_1298_Q_reg( .D(n5708), .CLK(CLK), .Q(n10618) );
	dfxbp_1 DFF_1214_Q_reg( .D(n5646), .CLK(CLK), .Q_N(n5917) );
	dfxtp_1 DFF_460_Q_reg( .D(n4590), .CLK(CLK), .Q(g8398) );
	dfxtp_1 DFF_478_Q_reg( .D(n5119), .CLK(CLK), .Q(n10616) );
	dfxbp_1 DFF_423_Q_reg( .D(n5078), .CLK(CLK), .Q_N(n5916) );
	dfxtp_1 DFF_1228_Q_reg( .D(n5655), .CLK(CLK), .Q(n10613) );
	dfxbp_1 DFF_1116_Q_reg( .D(n5568), .CLK(CLK), .Q(n11791), .Q_N(n5962) );
	dfxbp_1 DFF_288_Q_reg( .D(n4981), .CLK(CLK), .Q(n11842), .Q_N(n6063) );
	dfxbp_1 DFF_248_Q_reg( .D(n4949), .CLK(CLK), .Q(n11948), .Q_N(n5941) );
	dfxbp_1 DFF_1217_Q_reg( .D(n5649), .CLK(CLK), .Q(n11947), .Q_N(n5931) );
	dfxbp_1 DFF_1400_Q_reg( .D(n5783), .CLK(CLK), .Q_N(n5911) );
	dfxtp_1 DFF_503_Q_reg( .D(n4591), .CLK(CLK), .Q(g9615) );
	dfxtp_1 DFF_539_Q_reg( .D(n5158), .CLK(CLK), .Q(n10612) );
	dfxbp_1 DFF_1162_Q_reg( .D(n5602), .CLK(CLK), .Q_N(n5915) );
	dfxbp_1 DFF_543_Q_reg( .D(n5161), .CLK(CLK), .Q_N(n5913) );
	dfxtp_1 DFF_376_Q_reg( .D(n4589), .CLK(CLK), .Q(g9680) );
	dfxtp_1 DFF_396_Q_reg( .D(n5059), .CLK(CLK), .Q(n10609) );
	dfxtp_1 DFF_86_Q_reg( .D(n4587), .CLK(CLK), .Q(g9741) );
	dfxtp_1 DFF_838_Q_reg( .D(n5362), .CLK(CLK), .Q(n10607) );
	dfxbp_1 DFF_251_Q_reg( .D(n4952), .CLK(CLK), .Q_N(n5910) );
	dfxtp_1 DFF_371_Q_reg( .D(n4588), .CLK(CLK), .Q(g9817) );
	dfxtp_1 DFF_732_Q_reg( .D(n5290), .CLK(CLK), .Q(n10605) );
	dfxbp_1 DFF_1130_Q_reg( .D(n5578), .CLK(CLK), .Q_N(n5912) );
	dfxtp_1 DFF_961_Q_reg( .D(n4600), .CLK(CLK), .Q(g65) );
	dfxbp_1 DFF_186_Q_reg( .D(n4901), .CLK(CLK), .Q(n11847), .Q_N(n5949) );
	dfxbp_1 DFF_184_Q_reg( .D(n4900), .CLK(CLK), .Q_N(n5957) );
	dfxbp_1 DFF_436_Q_reg( .D(n5088), .CLK(CLK), .Q_N(n5956) );
	dfxbp_1 DFF_1399_Q_reg( .D(n5782), .CLK(CLK), .Q(n11779) );
	dfxbp_1 DFF_1107_Q_reg( .D(n5562), .CLK(CLK), .Q(n11961), .Q_N(n6071) );
	dfxbp_1 DFF_935_Q_reg( .D(n5438), .CLK(CLK), .Q(n11906), .Q_N(n5875) );
	dfxbp_1 DFF_796_Q_reg( .D(n5338), .CLK(CLK), .Q(n11777) );
	dfxbp_1 DFF_699_Q_reg( .D(n5265), .CLK(CLK), .Q(n11872), .Q_N(n5874) );
	dfxbp_1 DFF_604_Q_reg( .D(n5202), .CLK(CLK), .Q(n11898), .Q_N(n6073) );
	dfxtp_1 DFF_607_Q_reg( .D(n4610), .CLK(CLK), .Q(g4531) );
	dfxtp_1 DFF_1299_Q_reg( .D(n5709), .CLK(CLK), .Q(n10667) );
	dfxbp_1 DFF_609_Q_reg( .D(n5205), .CLK(CLK), .Q(n11967) );
	dfxbp_1 DFF_417_Q_reg( .D(n5075), .CLK(CLK), .Q(n11973) );
	dfxbp_1 DFF_1311_Q_reg( .D(n5716), .CLK(CLK), .Q(n11941) );
	dfxbp_1 DFF_1121_Q_reg( .D(n5571), .CLK(CLK), .Q(n11790), .Q_N(n5947) );
	dfxbp_1 DFF_1211_Q_reg( .D(n5643), .CLK(CLK), .Q(n11909), .Q_N(n6054) );
	dfxbp_1 DFF_1284_Q_reg( .D(n5698), .CLK(CLK), .Q_N(n6041) );
	dfxbp_1 DFF_1006_Q_reg( .D(n5488), .CLK(CLK), .Q(n11801) );
	dfxbp_1 DFF_743_Q_reg( .D(n5298), .CLK(CLK), .Q(n11769) );
	dfxbp_1 DFF_207_Q_reg( .D(n4915), .CLK(CLK), .Q(n11890) );
	dfxbp_1 DFF_679_Q_reg( .D(n5249), .CLK(CLK), .Q(n11768), .Q_N(n6043) );
	dfxbp_1 DFF_213_Q_reg( .D(n4921), .CLK(CLK), .Q(n11919), .Q_N(n6056) );
	dfxbp_1 DFF_249_Q_reg( .D(n4950), .CLK(CLK), .Q(n11844), .Q_N(n6091) );
	dfxbp_1 DFF_922_Q_reg( .D(n5427), .CLK(CLK), .Q(n11810) );
	dfxbp_1 DFF_1424_Q_reg( .D(n5800), .CLK(CLK), .Q(n11879) );
	dfxbp_1 DFF_78_Q_reg( .D(n4824), .CLK(CLK), .Q(n11916) );
	dfxbp_1 DFF_443_Q_reg( .D(n5092), .CLK(CLK), .Q(n11917) );
	dfxbp_1 DFF_1409_Q_reg( .D(n5790), .CLK(CLK), .Q_N(n6038) );
	dfxtp_1 DFF_1302_Q_reg( .D(n5710), .CLK(CLK), .Q(n10184) );
	dfxbp_1 DFF_696_Q_reg( .D(n5262), .CLK(CLK), .Q(n11889), .Q_N(n6059) );
	dfxbp_1 DFF_697_Q_reg( .D(n5263), .CLK(CLK), .Q(n11821) );
	dfxbp_1 DFF_684_Q_reg( .D(n5253), .CLK(CLK), .Q(n11905) );
	dfxbp_1 DFF_688_Q_reg( .D(n5256), .CLK(CLK), .Q(n11760), .Q_N(n5946) );
	dfxbp_1 DFF_955_Q_reg( .D(n5453), .CLK(CLK), .Q(n11884), .Q_N(n6061) );
	dfxbp_1 DFF_243_Q_reg( .D(n4945), .CLK(CLK), .Q(n11765), .Q_N(n6039) );
	dfxbp_1 DFF_535_Q_reg( .D(n5156), .CLK(CLK), .Q(n11831), .Q_N(n6081) );
	dfxbp_1 DFF_313_Q_reg( .D(n5003), .CLK(CLK), .Q(n11910) );
	dfxbp_1 DFF_987_Q_reg( .D(n5476), .CLK(CLK), .Q(n11802), .Q_N(n6042) );
	dfxbp_1 DFF_1278_Q_reg( .D(n5693), .CLK(CLK), .Q(n11878), .Q_N(n6057) );
	dfxbp_1 DFF_332_Q_reg( .D(n5015), .CLK(CLK), .Q(n11888), .Q_N(n6089) );
	dfxbp_1 DFF_714_Q_reg( .D(n50), .CLK(CLK), .Q(n11766), .Q_N(n6090) );
	dfxbp_1 DFF_742_Q_reg( .D(n5297), .CLK(CLK), .Q(n11860), .Q_N(n5878) );
	dfxbp_1 DFF_274_Q_reg( .D(n4969), .CLK(CLK), .Q(n11911), .Q_N(n6055) );
	dfxbp_1 DFF_1260_Q_reg( .D(n5679), .CLK(CLK), .Q_N(n6040) );
	dfxbp_1 DFF_857_Q_reg( .D(n5377), .CLK(CLK), .Q_N(n5968) );
	dfxbp_1 DFF_221_Q_reg( .D(n39), .CLK(CLK), .Q(n11908) );
	dfxtp_1 DFF_439_Q_reg( .D(n4606), .CLK(CLK), .Q(g4578) );
	dfxbp_1 DFF_1203_Q_reg( .D(n5636), .CLK(CLK), .Q(n11918), .Q_N(n6044) );
	dfxbp_1 DFF_1004_Q_reg( .D(n5487), .CLK(CLK), .Q(n11881), .Q_N(n6060) );
	dfxbp_1 DFF_287_Q_reg( .D(n4980), .CLK(CLK), .Q(n11887), .Q_N(n6099) );
	dfxbp_1 DFF_493_Q_reg( .D(n5128), .CLK(CLK), .Q(n11832), .Q_N(n6087) );
	dfxbp_1 DFF_1021_Q_reg( .D(n5500), .CLK(CLK), .Q(n11798), .Q_N(n5879) );
	dfxtp_1 DFF_1079_Q_reg( .D(n5542), .CLK(CLK), .Q(n10217) );
	dfxbp_1 DFF_1018_Q_reg( .D(n5498), .CLK(CLK), .Q(n11880), .Q_N(n6058) );
	dfxtp_1 DFF_310_Q_reg( .D(n5000), .CLK(CLK), .Q(n10610) );
	dfxbp_1 DFF_1205_Q_reg( .D(n5638), .CLK(CLK), .Q(n11787) );
	dfxtp_1 DFF_1345_Q_reg( .D(n4572), .CLK(CLK), .Q(g4519) );
	dfxtp_1 DFF_991_Q_reg( .D(n4569), .CLK(CLK), .Q(g4520) );
	dfxbp_1 DFF_1209_Q_reg( .D(n5641), .CLK(CLK), .Q_N(n5967) );
	dfxbp_1 DFF_383_Q_reg( .D(n5049), .CLK(CLK), .Q_N(n5880) );
	dfxbp_1 DFF_911_Q_reg( .D(n5418), .CLK(CLK), .Q_N(n5865) );
	dfxbp_1 DFF_129_Q_reg( .D(n4862), .CLK(CLK), .Q_N(n5870) );
	dfxtp_1 DFF_1415_Q_reg( .D(n5794), .CLK(CLK), .Q(n10213) );
	dfxbp_1 DFF_26_Q_reg( .D(n4782), .CLK(CLK), .Q_N(n19467) );
	dfxtp_1 DFF_624_Q_reg( .D(n4611), .CLK(CLK), .Q(g4480) );
	dfxtp_1 DFF_268_Q_reg( .D(n4604), .CLK(CLK), .Q(g4495) );
	dfxtp_1 DFF_352_Q_reg( .D(n4605), .CLK(CLK), .Q(g4498) );
	dfxtp_1 DFF_744_Q_reg( .D(n4612), .CLK(CLK), .Q(g4501) );
	dfxbp_1 DFF_384_Q_reg( .D(n5050), .CLK(CLK), .Q_N(n19451) );
	dfxtp_1 DFF_1296_Q_reg( .D(n5706), .CLK(CLK), .Q(n10880) );
	dfxbp_1 DFF_813_Q_reg( .D(n5350), .CLK(CLK), .Q(n11896), .Q_N(n6067) );
	dfxtp_1 DFF_1265_Q_reg( .D(n4586), .CLK(CLK), .Q(g10306) );
	dfxbp_1 DFF_663_Q_reg( .D(n91), .CLK(CLK), .Q_N(n5959) );
	dfxtp_1 DFF_234_Q_reg( .D(n4578), .CLK(CLK), .Q(g7257) );
	dfxtp_1 DFF_613_Q_reg( .D(n5207), .CLK(CLK), .Q(n10448) );
	dfxtp_1 DFF_1073_Q_reg( .D(n4576), .CLK(CLK), .Q(g7243) );
	dfxbp_1 DFF_1002_Q_reg( .D(n5485), .CLK(CLK), .Q(n11949), .Q_N(n6078) );
	dfxtp_1 DFF_1305_Q_reg( .D(n4571), .CLK(CLK), .Q(g26959) );
	dfxtp_1 DFF_530_Q_reg( .D(n4609), .CLK(CLK), .Q(g4455) );
	dfxtp_1 DFF_1146_Q_reg( .D(n5592), .CLK(CLK), .Q(n10519) );
	dfxbp_1 DFF_250_Q_reg( .D(n4951), .CLK(CLK), .Q(n11882), .Q_N(n5883) );
	dfxtp_1 DFF_348_Q_reg( .D(n4579), .CLK(CLK), .Q(g7260) );
	dfxtp_1 DFF_1225_Q_reg( .D(n4577), .CLK(CLK), .Q(g7245) );
	dfxtp_1 DFF_1272_Q_reg( .D(n5688), .CLK(CLK), .Q(n10602) );
	dfxtp_1 DFF_1411_Q_reg( .D(n4574), .CLK(CLK), .Q(g12832) );
	dfxbp_1 DFF_350_Q_reg( .D(n5028), .CLK(CLK), .Q(n11965) );
	dfxtp_1 DFF_1022_Q_reg( .D(n4615), .CLK(CLK), .Q(g4540) );
	dfxtp_1 DFF_226_Q_reg( .D(n4603), .CLK(CLK), .Q(g4543) );
	dfxtp_1 DFF_56_Q_reg( .D(n4601), .CLK(CLK), .Q(g4567) );
	dfxtp_1 DFF_816_Q_reg( .D(n4613), .CLK(CLK), .Q(g4546) );
	dfxbp_1 DFF_1330_Q_reg( .D(n5729), .CLK(CLK), .Q_N(n19450) );
	dfxtp_1 DFF_1362_Q_reg( .D(n4570), .CLK(CLK), .Q(g4570) );
	dfxtp_1 DFF_528_Q_reg( .D(n4568), .CLK(CLK), .Q(g4571) );
	dfxbp_1 DFF_38_Q_reg( .D(n4791), .CLK(CLK), .Q(n11885), .Q_N(n6083) );
	dfxbp_1 DFF_121_Q_reg( .D(n4858), .CLK(CLK), .Q_N(n5951) );
	dfxbp_1 DFF_808_Q_reg( .D(n5345), .CLK(CLK), .Q(n11886), .Q_N(n6086) );
	dfxtp_1 DFF_491_Q_reg( .D(n4608), .CLK(CLK), .Q(g4564) );
	dfxbp_1 DFF_228_Q_reg( .D(n4932), .CLK(CLK), .Q(n11845) );
	dfxtp_1 DFF_1397_Q_reg( .D(n5780), .CLK(CLK), .Q(n10231) );
	dfxbp_1 DFF_749_Q_reg( .D(n5303), .CLK(CLK), .Q(n11818), .Q_N(n6065) );
	dfxtp_1 DFF_413_Q_reg( .D(n5073), .CLK(CLK), .Q(n10429) );
	dfxbp_1 DFF_1289_Q_reg( .D(n5701), .CLK(CLK), .Q(n11774), .Q_N(n5897) );
	dfxbp_1 DFF_311_Q_reg( .D(n5001), .CLK(CLK), .Q(n11838), .Q_N(n5906) );
	dfxbp_1 DFF_1381_Q_reg( .D(n5767), .CLK(CLK), .Q_N(n20311) );
	dfxtp_1 DFF_206_Q_reg( .D(n5144), .CLK(CLK), .Q(g52) );
	dfxtp_1 DFF_621_Q_reg( .D(n4599), .CLK(CLK), .Q(g55) );
	dfxtp_1 DFF_1074_Q_reg( .D(n4599), .CLK(CLK), .Q(n10232) );
	dfxtp_1 DFF_477_Q_reg( .D(n4607), .CLK(CLK), .Q(g46) );
	dfxbp_1 DFF_1222_Q_reg( .D(n4607), .CLK(CLK), .Q(n11971) );
	dfxbp_1 DFF_619_Q_reg( .D(n5210), .CLK(CLK), .Q(n11970) );
	dfxbp_1 DFF_355_Q_reg( .D(n5031), .CLK(CLK), .Q(n11835) );
	dfxtp_1 DFF_829_Q_reg( .D(n4614), .CLK(CLK), .Q(g47) );
	dfxbp_1 DFF_761_Q_reg( .D(n4614), .CLK(CLK), .Q(n11969) );
	dfxtp_1 DFF_150_Q_reg( .D(n5164), .CLK(CLK), .Q(g48) );
	dfxtp_1 DFF_1322_Q_reg( .D(n5031), .CLK(CLK), .Q(g49) );
	dfxtp_1 DFF_514_Q_reg( .D(n5210), .CLK(CLK), .Q(g45) );
	dfxtp_1 DFF_420_Q_reg( .D(n5332), .CLK(CLK), .Q(g51) );
	dfxtp_1 DFF_1012_Q_reg( .D(n5656), .CLK(CLK), .Q(g50) );
	dfxtp_1 DFF_1157_Q_reg( .D(n5598), .CLK(CLK), .Q(n10474) );
	dfxtp_1 DFF_276_Q_reg( .D(n4971), .CLK(CLK), .Q(n10475) );
	dfxtp_1 DFF_766_Q_reg( .D(n5313), .CLK(CLK), .Q(n10708) );
	dfxtp_1 DFF_215_Q_reg( .D(n4923), .CLK(CLK), .Q(n10925) );
	dfxtp_1 DFF_210_Q_reg( .D(n4918), .CLK(CLK), .Q(n10876) );
	dfxtp_1 DFF_756_Q_reg( .D(n5308), .CLK(CLK), .Q(n10549) );
	dfxtp_1 DFF_1269_Q_reg( .D(n5686), .CLK(CLK), .Q(n10485) );
	dfxtp_1 DFF_527_Q_reg( .D(n4702), .CLK(CLK), .Q(g25689) );
	dfxtp_1 DFF_434_Q_reg( .D(n5086), .CLK(CLK), .Q(n10291) );
	dfxtp_1 DFF_126_Q_reg( .D(n4702), .CLK(CLK), .Q(g24265) );
	dfxtp_1 DFF_893_Q_reg( .D(n5406), .CLK(CLK), .Q(n10363) );
	dfxtp_1 DFF_69_Q_reg( .D(n4816), .CLK(CLK), .Q(n10861) );
	dfxtp_1 DFF_236_Q_reg( .D(n4938), .CLK(CLK), .Q(n10862) );
	dfxtp_1 DFF_608_Q_reg( .D(n5204), .CLK(CLK), .Q(n10860) );
	dfxtp_1 DFF_1262_Q_reg( .D(n4669), .CLK(CLK), .Q(g14635) );
	dfxtp_1 DFF_836_Q_reg( .D(n4666), .CLK(CLK), .Q(g14749) );
	dfxtp_1 DFF_537_Q_reg( .D(n4664), .CLK(CLK), .Q(g14597) );
	dfxtp_1 DFF_76_Q_reg( .D(n4662), .CLK(CLK), .Q(g13865) );
	dfxtp_1 DFF_369_Q_reg( .D(n4663), .CLK(CLK), .Q(g13881) );
	dfxtp_1 DFF_662_Q_reg( .D(n4665), .CLK(CLK), .Q(g13906) );
	dfxtp_1 DFF_1102_Q_reg( .D(n4668), .CLK(CLK), .Q(g14673) );
	dfxtp_1 DFF_905_Q_reg( .D(n4667), .CLK(CLK), .Q(g14705) );
	dfxtp_1 DFF_601_Q_reg( .D(n5199), .CLK(CLK), .Q(n10355) );
	dfxtp_1 DFF_1315_Q_reg( .D(n5720), .CLK(CLK), .Q(n10421) );
	dfxtp_1 DFF_194_Q_reg( .D(n4907), .CLK(CLK), .Q(n10713) );
	dfxtp_1 DFF_338_Q_reg( .D(n5019), .CLK(CLK), .Q(n10589) );
	dfxtp_1 DFF_789_Q_reg( .D(n5331), .CLK(CLK), .Q(n10395) );
	dfxtp_1 DFF_83_Q_reg( .D(n4828), .CLK(CLK), .Q(n10540) );
	dfxtp_1 DFF_359_Q_reg( .D(n5034), .CLK(CLK), .Q(n10544) );
	dfxtp_1 DFF_582_Q_reg( .D(n5186), .CLK(CLK), .Q(n10563) );
	dfxtp_1 DFF_593_Q_reg( .D(n5194), .CLK(CLK), .Q(n10871) );
	dfxtp_1 DFF_788_Q_reg( .D(n5330), .CLK(CLK), .Q(n10387) );
	dfxtp_1 DFF_1241_Q_reg( .D(n5665), .CLK(CLK), .Q(n10570) );
	dfxtp_1 DFF_859_Q_reg( .D(n5379), .CLK(CLK), .Q(n10542) );
	dfxtp_1 DFF_867_Q_reg( .D(n5386), .CLK(CLK), .Q(n10905) );
	dfxtp_1 DFF_1274_Q_reg( .D(n5690), .CLK(CLK), .Q(n10911) );
	dfxtp_1 DFF_901_Q_reg( .D(n5413), .CLK(CLK), .Q(n10569) );
	dfxtp_1 DFF_454_Q_reg( .D(n5102), .CLK(CLK), .Q(n10541) );
	dfxtp_1 DFF_1109_Q_reg( .D(n5564), .CLK(CLK), .Q(n10904) );
	dfxtp_1 DFF_1153_Q_reg( .D(n5596), .CLK(CLK), .Q(n10386) );
	dfxtp_1 DFF_720_Q_reg( .D(n5279), .CLK(CLK), .Q(n10907) );
	dfxtp_1 DFF_1041_Q_reg( .D(n5516), .CLK(CLK), .Q(n10863) );
	dfxtp_1 DFF_1234_Q_reg( .D(n4717), .CLK(CLK), .Q(g11447) );
	dfxtp_1 DFF_480_Q_reg( .D(n4722), .CLK(CLK), .Q(g8783) );
	dfxtp_1 DFF_909_Q_reg( .D(n4726), .CLK(CLK), .Q(g8784) );
	dfxtp_1 DFF_565_Q_reg( .D(n4724), .CLK(CLK), .Q(g8785) );
	dfxtp_1 DFF_1224_Q_reg( .D(n4688), .CLK(CLK), .Q(g8786) );
	dfxtp_1 DFF_1416_Q_reg( .D(n4720), .CLK(CLK), .Q(g8787) );
	dfxtp_1 DFF_704_Q_reg( .D(n4716), .CLK(CLK), .Q(g8789) );
	dfxtp_1 DFF_707_Q_reg( .D(n5270), .CLK(CLK), .Q(n10827) );
	dfxtp_1 DFF_638_Q_reg( .D(n5223), .CLK(CLK), .Q(n10801) );
	dfxtp_1 DFF_659_Q_reg( .D(n5238), .CLK(CLK), .Q(n10798) );
	dfxtp_1 DFF_479_Q_reg( .D(n5120), .CLK(CLK), .Q(n10813) );
	dfxtp_1 DFF_627_Q_reg( .D(n5216), .CLK(CLK), .Q(n10787) );
	dfxtp_1 DFF_884_Q_reg( .D(n5398), .CLK(CLK), .Q(n10785) );
	dfxtp_1 DFF_938_Q_reg( .D(n5440), .CLK(CLK), .Q(n10786) );
	dfxtp_1 DFF_84_Q_reg( .D(n4829), .CLK(CLK), .Q(n10782) );
	dfxtp_1 DFF_267_Q_reg( .D(n4964), .CLK(CLK), .Q(n10775) );
	dfxtp_1 DFF_947_Q_reg( .D(n5445), .CLK(CLK), .Q(n10811) );
	dfxtp_1 DFF_72_Q_reg( .D(n4819), .CLK(CLK), .Q(n10824) );
	dfxtp_1 DFF_982_Q_reg( .D(n5471), .CLK(CLK), .Q(n10828) );
	dfxtp_1 DFF_877_Q_reg( .D(n5393), .CLK(CLK), .Q(n10772) );
	dfxtp_1 DFF_526_Q_reg( .D(n5151), .CLK(CLK), .Q(n10776) );
	dfxtp_1 DFF_392_Q_reg( .D(n5056), .CLK(CLK), .Q(n10781) );
	dfxtp_1 DFF_219_Q_reg( .D(n4926), .CLK(CLK), .Q(n10783) );
	dfxtp_1 DFF_1350_Q_reg( .D(n5744), .CLK(CLK), .Q(n10812) );
	dfxtp_1 DFF_1218_Q_reg( .D(n5650), .CLK(CLK), .Q(n10839) );
	dfxtp_1 DFF_670_Q_reg( .D(n5244), .CLK(CLK), .Q(n10837) );
	dfxtp_1 DFF_1386_Q_reg( .D(n5771), .CLK(CLK), .Q(n10838) );
	dfxtp_1 DFF_1174_Q_reg( .D(n5611), .CLK(CLK), .Q(n10749) );
	dfxtp_1 DFF_617_Q_reg( .D(n5209), .CLK(CLK), .Q(n10746) );
	dfxtp_1 DFF_967_Q_reg( .D(n5463), .CLK(CLK), .Q(n10750) );
	dfxtp_1 DFF_1197_Q_reg( .D(n5630), .CLK(CLK), .Q(n10830) );
	dfxtp_1 DFF_1401_Q_reg( .D(n5784), .CLK(CLK), .Q(n10833) );
	dfxtp_1 DFF_1351_Q_reg( .D(n5745), .CLK(CLK), .Q(n10831) );
	dfxtp_1 DFF_1208_Q_reg( .D(n5640), .CLK(CLK), .Q(n10832) );
	dfxtp_1 DFF_156_Q_reg( .D(n4880), .CLK(CLK), .Q(n10808) );
	dfxtp_1 DFF_986_Q_reg( .D(n5475), .CLK(CLK), .Q(n10807) );
	dfxtp_1 DFF_550_Q_reg( .D(n5165), .CLK(CLK), .Q(n10809) );
	dfxtp_1 DFF_91_Q_reg( .D(n4834), .CLK(CLK), .Q(n10806) );
	dfxtp_1 DFF_1259_Q_reg( .D(n5678), .CLK(CLK), .Q(n10817) );
	dfxtp_1 DFF_321_Q_reg( .D(n5009), .CLK(CLK), .Q(n10820) );
	dfxtp_1 DFF_241_Q_reg( .D(n4943), .CLK(CLK), .Q(n10765) );
	dfxtp_1 DFF_920_Q_reg( .D(n5425), .CLK(CLK), .Q(n10768) );
	dfxtp_1 DFF_1201_Q_reg( .D(n5634), .CLK(CLK), .Q(n10766) );
	dfxtp_1 DFF_17_Q_reg( .D(n4773), .CLK(CLK), .Q(n10767) );
	dfxtp_1 DFF_610_Q_reg( .D(n5206), .CLK(CLK), .Q(n10739) );
	dfxtp_1 DFF_1294_Q_reg( .D(n5704), .CLK(CLK), .Q(n10742) );
	dfxtp_1 DFF_738_Q_reg( .D(n5295), .CLK(CLK), .Q(n10818) );
	dfxtp_1 DFF_309_Q_reg( .D(n4999), .CLK(CLK), .Q(n10819) );
	dfxtp_1 DFF_1024_Q_reg( .D(n5502), .CLK(CLK), .Q(n10740) );
	dfxtp_1 DFF_1169_Q_reg( .D(n5607), .CLK(CLK), .Q(n10741) );
	dfxtp_1 DFF_1011_Q_reg( .D(n5493), .CLK(CLK), .Q(n10761) );
	dfxtp_1 DFF_1366_Q_reg( .D(n5755), .CLK(CLK), .Q(n10759) );
	dfxtp_1 DFF_494_Q_reg( .D(n5129), .CLK(CLK), .Q(n10760) );
	dfxtp_1 DFF_314_Q_reg( .D(n5004), .CLK(CLK), .Q(n10756) );
	dfxtp_1 DFF_634_Q_reg( .D(n5220), .CLK(CLK), .Q(n10755) );
	dfxtp_1 DFF_1123_Q_reg( .D(n5572), .CLK(CLK), .Q(n10757) );
	dfxtp_1 DFF_158_Q_reg( .D(n4882), .CLK(CLK), .Q(n10754) );
	dfxtp_1 DFF_100_Q_reg( .D(n4842), .CLK(CLK), .Q(n10802) );
	dfxtp_1 DFF_390_Q_reg( .D(n5055), .CLK(CLK), .Q(n10791) );
	dfxtp_1 DFF_13_Q_reg( .D(n4769), .CLK(CLK), .Q(n10794) );
	dfxtp_1 DFF_750_Q_reg( .D(n5304), .CLK(CLK), .Q(n10792) );
	dfxtp_1 DFF_602_Q_reg( .D(n5200), .CLK(CLK), .Q(n10793) );
	dfxtp_1 DFF_1007_Q_reg( .D(n5489), .CLK(CLK), .Q(n10780) );
	dfxtp_1 DFF_637_Q_reg( .D(n5222), .CLK(CLK), .Q(n10728) );
	dfxtp_1 DFF_682_Q_reg( .D(n5251), .CLK(CLK), .Q(n10726) );
	dfxtp_1 DFF_1050_Q_reg( .D(n5522), .CLK(CLK), .Q(n10729) );
	dfxtp_1 DFF_442_Q_reg( .D(n5091), .CLK(CLK), .Q(n10727) );
	dfxtp_1 DFF_77_Q_reg( .D(n4823), .CLK(CLK), .Q(n10730) );
	dfxtp_1 DFF_1266_Q_reg( .D(n5683), .CLK(CLK), .Q(n10733) );
	dfxtp_1 DFF_1180_Q_reg( .D(n5617), .CLK(CLK), .Q(n10737) );
	dfxtp_1 DFF_832_Q_reg( .D(n5358), .CLK(CLK), .Q(n10731) );
	dfxtp_1 DFF_1114_Q_reg( .D(n5566), .CLK(CLK), .Q(n10732) );
	dfxtp_1 DFF_702_Q_reg( .D(n5267), .CLK(CLK), .Q(n10623) );
	dfxtp_1 DFF_903_Q_reg( .D(n5415), .CLK(CLK), .Q(n10626) );
	dfxtp_1 DFF_558_Q_reg( .D(n5169), .CLK(CLK), .Q(n10634) );
	dfxtp_1 DFF_216_Q_reg( .D(n4924), .CLK(CLK), .Q(n10625) );
	dfxtp_1 DFF_1086_Q_reg( .D(n5548), .CLK(CLK), .Q(n10627) );
	dfxtp_1 DFF_264_Q_reg( .D(n4962), .CLK(CLK), .Q(n10635) );
	dfxtp_1 DFF_212_Q_reg( .D(n4920), .CLK(CLK), .Q(n10630) );
	dfxtp_1 DFF_1226_Q_reg( .D(n5653), .CLK(CLK), .Q(n10638) );
	dfxtp_1 DFF_912_Q_reg( .D(n5419), .CLK(CLK), .Q(n10628) );
	dfxtp_1 DFF_1268_Q_reg( .D(n5685), .CLK(CLK), .Q(n10624) );
	dfxtp_1 DFF_6_Q_reg( .D(n4764), .CLK(CLK), .Q(n10632) );
	dfxtp_1 DFF_649_Q_reg( .D(n5231), .CLK(CLK), .Q(n10629) );
	dfxtp_1 DFF_882_Q_reg( .D(n5396), .CLK(CLK), .Q(n10637) );
	dfxtp_1 DFF_389_Q_reg( .D(n4721), .CLK(CLK), .Q(g11770) );
	dfxtp_1 DFF_1286_Q_reg( .D(n4718), .CLK(CLK), .Q(g8915) );
	dfxtp_1 DFF_485_Q_reg( .D(n4723), .CLK(CLK), .Q(g8916) );
	dfxtp_1 DFF_992_Q_reg( .D(n4727), .CLK(CLK), .Q(g8917) );
	dfxtp_1 DFF_418_Q_reg( .D(n4715), .CLK(CLK), .Q(g8918) );
	dfxtp_1 DFF_1338_Q_reg( .D(n4719), .CLK(CLK), .Q(g8920) );
	dfxtp_1 DFF_31_Q_reg( .D(n4786), .CLK(CLK), .Q(n10891) );
	dfxtp_1 DFF_674_Q_reg( .D(n5247), .CLK(CLK), .Q(n10407) );
	dfxtp_1 DFF_1029_Q_reg( .D(n5506), .CLK(CLK), .Q(n10190) );
	dfxtp_1 DFF_747_Q_reg( .D(n5301), .CLK(CLK), .Q(n10935) );
	dfxtp_1 DFF_456_Q_reg( .D(n5104), .CLK(CLK), .Q(n10867) );
	dfxtp_1 DFF_1398_Q_reg( .D(n5781), .CLK(CLK), .Q(n10651) );
	dfxtp_1 DFF_632_Q_reg( .D(n5218), .CLK(CLK), .Q(n10641) );
	dfxtp_1 DFF_1332_Q_reg( .D(n5731), .CLK(CLK), .Q(n10649) );
	dfxtp_1 DFF_356_Q_reg( .D(n5032), .CLK(CLK), .Q(n10654) );
	dfxtp_1 DFF_341_Q_reg( .D(n5021), .CLK(CLK), .Q(n10645) );
	dfxtp_1 DFF_29_Q_reg( .D(n4785), .CLK(CLK), .Q(n10653) );
	dfxtp_1 DFF_433_Q_reg( .D(n5085), .CLK(CLK), .Q(n10639) );
	dfxtp_1 DFF_1154_Q_reg( .D(n5597), .CLK(CLK), .Q(n10647) );
	dfxtp_1 DFF_782_Q_reg( .D(n5327), .CLK(CLK), .Q(n10934) );
	dfxtp_1 DFF_693_Q_reg( .D(n5260), .CLK(CLK), .Q(n10644) );
	dfxtp_1 DFF_441_Q_reg( .D(n5090), .CLK(CLK), .Q(n10868) );
	dfxtp_1 DFF_1383_Q_reg( .D(n5769), .CLK(CLK), .Q(n10652) );
	dfxtp_1 DFF_275_Q_reg( .D(n4970), .CLK(CLK), .Q(n10648) );
	dfxtp_1 DFF_388_Q_reg( .D(n5054), .CLK(CLK), .Q(n10650) );
	dfxtp_1 DFF_687_Q_reg( .D(n5255), .CLK(CLK), .Q(n10873) );
	dfxtp_1 DFF_490_Q_reg( .D(n5127), .CLK(CLK), .Q(n10929) );
	dfxtp_1 DFF_692_Q_reg( .D(n5259), .CLK(CLK), .Q(n10933) );
	dfxtp_1 DFF_781_Q_reg( .D(n5326), .CLK(CLK), .Q(n10578) );
	dfxtp_1 DFF_15_Q_reg( .D(n4771), .CLK(CLK), .Q(n10701) );
	dfxtp_1 DFF_1336_Q_reg( .D(n5732), .CLK(CLK), .Q(n10709) );
	dfxtp_1 DFF_1139_Q_reg( .D(n5586), .CLK(CLK), .Q(n10858) );
	dfxtp_1 DFF_0_Q_reg( .D(n5801), .CLK(CLK), .Q(n10682) );
	dfxtp_1 DFF_154_Q_reg( .D(n4878), .CLK(CLK), .Q(n10162) );
	dfxtp_1 DFF_997_Q_reg( .D(n4712), .CLK(CLK), .Q(g8235) );
	dfxtp_1 DFF_686_Q_reg( .D(n4707), .CLK(CLK), .Q(g7540) );
	dfxtp_1 DFF_254_Q_reg( .D(n4955), .CLK(CLK), .Q(n10599) );
	dfxtp_1 DFF_1206_Q_reg( .D(n5639), .CLK(CLK), .Q(n10596) );
	dfxtp_1 DFF_710_Q_reg( .D(n5272), .CLK(CLK), .Q(n10427) );
	dfxtp_1 DFF_270_Q_reg( .D(n4965), .CLK(CLK), .Q(n10461) );
	dfxtp_1 DFF_630_Q_reg( .D(n4706), .CLK(CLK), .Q(g9555) );
	dfxtp_1 DFF_85_Q_reg( .D(n4696), .CLK(CLK), .Q(g9617) );
	dfxtp_1 DFF_1316_Q_reg( .D(n4714), .CLK(CLK), .Q(g9682) );
	dfxtp_1 DFF_317_Q_reg( .D(n4699), .CLK(CLK), .Q(g8215) );
	dfxtp_1 DFF_861_Q_reg( .D(n4710), .CLK(CLK), .Q(g9743) );
	dfxtp_1 DFF_147_Q_reg( .D(n4697), .CLK(CLK), .Q(g8344) );
	dfxtp_1 DFF_830_Q_reg( .D(n4709), .CLK(CLK), .Q(g8279) );
	dfxtp_1 DFF_1118_Q_reg( .D(n4695), .CLK(CLK), .Q(g8353) );
	dfxtp_1 DFF_1100_Q_reg( .D(n4694), .CLK(CLK), .Q(g8403) );
	dfxtp_1 DFF_981_Q_reg( .D(n4711), .CLK(CLK), .Q(g8283) );
	dfxtp_1 DFF_615_Q_reg( .D(n4705), .CLK(CLK), .Q(g26960) );
	dfxtp_1 DFF_585_Q_reg( .D(n4704), .CLK(CLK), .Q(g14189) );
	dfxtp_1 DFF_561_Q_reg( .D(n4703), .CLK(CLK), .Q(g14201) );
	dfxtp_1 DFF_1106_Q_reg( .D(n4713), .CLK(CLK), .Q(g14217) );
	dfxtp_1 DFF_152_Q_reg( .D(n4698), .CLK(CLK), .Q(g14096) );
	dfxtp_1 DFF_404_Q_reg( .D(n4701), .CLK(CLK), .Q(g14125) );
	dfxtp_1 DFF_380_Q_reg( .D(n4700), .CLK(CLK), .Q(g14147) );
	dfxtp_1 DFF_764_Q_reg( .D(n4708), .CLK(CLK), .Q(g14167) );
	dfxtp_1 DFF_647_Q_reg( .D(n5229), .CLK(CLK), .Q(n10598) );
	dfxtp_1 DFF_229_Q_reg( .D(n4933), .CLK(CLK), .Q(n10594) );
	dfxtp_1 DFF_574_Q_reg( .D(n5179), .CLK(CLK), .Q(n10595) );
	dfxtp_1 DFF_778_Q_reg( .D(n5324), .CLK(CLK), .Q(n10869) );
	dfxtp_1 DFF_837_Q_reg( .D(n5361), .CLK(CLK), .Q(n10597) );
	dfxtp_1 DFF_52_Q_reg( .D(n4802), .CLK(CLK), .Q(n10866) );
	dfxtp_1 DFF_73_Q_reg( .D(n4820), .CLK(CLK), .Q(n10317) );
	dfxtp_1 DFF_70_Q_reg( .D(n4817), .CLK(CLK), .Q(n10560) );
	dfxtp_1 DFF_1227_Q_reg( .D(n5654), .CLK(CLK), .Q(n10559) );
	dfxtp_1 DFF_672_Q_reg( .D(n4725), .CLK(CLK), .Q(g8178) );
	dfxtp_1 DFF_178_Q_reg( .D(n4725), .CLK(CLK), .Q(g8132) );
	dfxtp_1 DFF_1059_Q_reg( .D(n4756), .CLK(CLK), .Q(g21176) );
	dfxtp_1 DFF_934_Q_reg( .D(n4691), .CLK(CLK), .Q(g18881) );
	dfxtp_1 DFF_1200_Q_reg( .D(n5633), .CLK(CLK), .Q(n10384) );
	dfxtp_1 DFF_416_Q_reg( .D(n46), .CLK(CLK), .Q(n10186) );
	dfxtp_1 DFF_1131_Q_reg( .D(n5579), .CLK(CLK), .Q(n10467) );
	dfxtp_1 DFF_502_Q_reg( .D(n5135), .CLK(CLK), .Q(n10359) );
	dfxtp_1 DFF_28_Q_reg( .D(n4784), .CLK(CLK), .Q(n10529) );
	dfxtp_1 DFF_157_Q_reg( .D(n4881), .CLK(CLK), .Q(n10393) );
	dfxtp_1 DFF_1151_Q_reg( .D(n5595), .CLK(CLK), .Q(n10712) );
	dfxtp_1 DFF_123_Q_reg( .D(n4643), .CLK(CLK), .Q(g17685) );
	dfxtp_1 DFF_23_Q_reg( .D(n4779), .CLK(CLK), .Q(n10308) );
	dfxtp_1 DFF_1407_Q_reg( .D(n5788), .CLK(CLK), .Q(n10468) );
	dfxtp_1 DFF_626_Q_reg( .D(n5215), .CLK(CLK), .Q(n10829) );
	dfxtp_1 DFF_728_Q_reg( .D(n5286), .CLK(CLK), .Q(n10534) );
	dfxtp_1 DFF_1282_Q_reg( .D(n5696), .CLK(CLK), .Q(n10700) );
	dfxtp_1 DFF_448_Q_reg( .D(n5097), .CLK(CLK), .Q(n10714) );
	dfxtp_1 DFF_519_Q_reg( .D(n5146), .CLK(CLK), .Q(n10511) );
	dfxtp_1 DFF_916_Q_reg( .D(n5422), .CLK(CLK), .Q(n10510) );
	dfxtp_1 DFF_587_Q_reg( .D(n5189), .CLK(CLK), .Q(n10512) );
	dfxtp_1 DFF_199_Q_reg( .D(n4911), .CLK(CLK), .Q(n10513) );
	dfxtp_1 DFF_1108_Q_reg( .D(n5563), .CLK(CLK), .Q(n10442) );
	dfxtp_1 DFF_542_Q_reg( .D(n5160), .CLK(CLK), .Q(n10734) );
	dfxtp_1 DFF_109_Q_reg( .D(n4670), .CLK(CLK), .Q(g9048) );
	dfxtp_1 DFF_343_Q_reg( .D(n5023), .CLK(CLK), .Q(n10689) );
	dfxtp_1 DFF_1124_Q_reg( .D(n21), .CLK(CLK), .Q(n10464) );
	dfxtp_1 DFF_130_Q_reg( .D(n4863), .CLK(CLK), .Q(n10230) );
	dfxtp_1 DFF_160_Q_reg( .D(n4883), .CLK(CLK), .Q(n10535) );
	dfxtp_1 DFF_107_Q_reg( .D(n4848), .CLK(CLK), .Q(n10229) );
	dfxtp_1 DFF_792_Q_reg( .D(n5334), .CLK(CLK), .Q(n10573) );
	dfxtp_1 DFF_855_Q_reg( .D(n5376), .CLK(CLK), .Q(n10706) );
	dfxtp_1 DFF_469_Q_reg( .D(n5113), .CLK(CLK), .Q(n10721) );
	dfxtp_1 DFF_809_Q_reg( .D(n5346), .CLK(CLK), .Q(n10723) );
	dfxtp_1 DFF_32_Q_reg( .D(n4787), .CLK(CLK), .Q(n10738) );
	dfxtp_1 DFF_504_Q_reg( .D(n5136), .CLK(CLK), .Q(n10724) );
	dfxtp_1 DFF_1137_Q_reg( .D(n5584), .CLK(CLK), .Q(n10725) );
	dfxtp_1 DFF_25_Q_reg( .D(n4781), .CLK(CLK), .Q(n10872) );
	dfxtp_1 DFF_1061_Q_reg( .D(n5531), .CLK(CLK), .Q(n10936) );
	dfxtp_1 DFF_677_Q_reg( .D(n5248), .CLK(CLK), .Q(n10710) );
	dfxtp_1 DFF_21_Q_reg( .D(n4777), .CLK(CLK), .Q(n10551) );
	dfxtp_1 DFF_1135_Q_reg( .D(n5582), .CLK(CLK), .Q(n10722) );
	dfxtp_1 DFF_959_Q_reg( .D(n5457), .CLK(CLK), .Q(n10720) );
	dfxtp_1 DFF_1081_Q_reg( .D(n4671), .CLK(CLK), .Q(g11678) );
	dfxtp_1 DFF_1412_Q_reg( .D(n5792), .CLK(CLK), .Q(n10687) );
	dfxtp_1 DFF_239_Q_reg( .D(n4941), .CLK(CLK), .Q(n10859) );
	dfxtp_1 DFF_128_Q_reg( .D(n4861), .CLK(CLK), .Q(n10895) );
	dfxtp_1 DFF_918_Q_reg( .D(n5424), .CLK(CLK), .Q(n10852) );
	dfxtp_1 DFF_839_Q_reg( .D(n5363), .CLK(CLK), .Q(n10856) );
	dfxtp_1 DFF_826_Q_reg( .D(n5357), .CLK(CLK), .Q(n10853) );
	dfxtp_1 DFF_644_Q_reg( .D(n5226), .CLK(CLK), .Q(n10849) );
	dfxtp_1 DFF_559_Q_reg( .D(n5170), .CLK(CLK), .Q(n10855) );
	dfxtp_1 DFF_136_Q_reg( .D(n4868), .CLK(CLK), .Q(n10850) );
	dfxtp_1 DFF_1195_Q_reg( .D(n5629), .CLK(CLK), .Q(n10854) );
	dfxtp_1 DFF_1138_Q_reg( .D(n5585), .CLK(CLK), .Q(n10851) );
	dfxtp_1 DFF_482_Q_reg( .D(n5121), .CLK(CLK), .Q(n10473) );
	dfxtp_1 DFF_1237_Q_reg( .D(n5663), .CLK(CLK), .Q(n10412) );
	dfxtp_1 DFF_1159_Q_reg( .D(n5599), .CLK(CLK), .Q(n10411) );
	dfxtp_1 DFF_161_Q_reg( .D(n4884), .CLK(CLK), .Q(n10707) );
	dfxtp_1 DFF_89_Q_reg( .D(n4832), .CLK(CLK), .Q(n10527) );
	dfxtp_1 DFF_340_Q_reg( .D(n5020), .CLK(CLK), .Q(n10814) );
	dfxtp_1 DFF_333_Q_reg( .D(n5016), .CLK(CLK), .Q(n10788) );
	dfxtp_1 DFF_151_Q_reg( .D(n4876), .CLK(CLK), .Q(n10778) );
	dfxtp_1 DFF_12_Q_reg( .D(n4768), .CLK(CLK), .Q(n10825) );
	dfxtp_1 DFF_645_Q_reg( .D(n5227), .CLK(CLK), .Q(n10834) );
	dfxtp_1 DFF_93_Q_reg( .D(n4836), .CLK(CLK), .Q(n10769) );
	dfxtp_1 DFF_183_Q_reg( .D(n4899), .CLK(CLK), .Q(n10771) );
	dfxtp_1 DFF_1032_Q_reg( .D(n5509), .CLK(CLK), .Q(n10747) );
	dfxtp_1 DFF_1175_Q_reg( .D(n5612), .CLK(CLK), .Q(n10743) );
	dfxtp_1 DFF_1356_Q_reg( .D(n5747), .CLK(CLK), .Q(n10823) );
	dfxtp_1 DFF_1348_Q_reg( .D(n5742), .CLK(CLK), .Q(n10745) );
	dfxtp_1 DFF_253_Q_reg( .D(n4954), .CLK(CLK), .Q(n10810) );
	dfxtp_1 DFF_1325_Q_reg( .D(n5725), .CLK(CLK), .Q(n10799) );
	dfxtp_1 DFF_1040_Q_reg( .D(n5515), .CLK(CLK), .Q(n10795) );
	dfxtp_1 DFF_1363_Q_reg( .D(n5752), .CLK(CLK), .Q(n10797) );
	dfxtp_1 DFF_1423_Q_reg( .D(n5799), .CLK(CLK), .Q(n10784) );
	dfxtp_1 DFF_721_Q_reg( .D(n5280), .CLK(CLK), .Q(n10711) );
	dfxtp_1 DFF_974_Q_reg( .D(n5467), .CLK(CLK), .Q(n10864) );
	dfxtp_1 DFF_864_Q_reg( .D(n5383), .CLK(CLK), .Q(n10930) );
	dfxtp_1 DFF_231_Q_reg( .D(n4934), .CLK(CLK), .Q(n10658) );
	dfxtp_1 DFF_177_Q_reg( .D(n4896), .CLK(CLK), .Q(n10659) );
	dfxtp_1 DFF_1250_Q_reg( .D(n5671), .CLK(CLK), .Q(n10857) );
	dfxtp_1 DFF_94_Q_reg( .D(n4837), .CLK(CLK), .Q(n10389) );
	dfxtp_1 DFF_1017_Q_reg( .D(n5497), .CLK(CLK), .Q(n10388) );
	dfxtp_1 DFF_1357_Q_reg( .D(n5748), .CLK(CLK), .Q(n10927) );
	dfxtp_1 DFF_142_Q_reg( .D(n4871), .CLK(CLK), .Q(n10926) );
	dfxtp_1 DFF_1403_Q_reg( .D(n5785), .CLK(CLK), .Q(n10699) );
	dfxtp_1 DFF_101_Q_reg( .D(n4641), .CLK(CLK), .Q(g17604) );
	dfxtp_1 DFF_524_Q_reg( .D(n5149), .CLK(CLK), .Q(n10372) );
	dfxtp_1 DFF_786_Q_reg( .D(n5329), .CLK(CLK), .Q(n10550) );
	dfxtp_1 DFF_208_Q_reg( .D(n4916), .CLK(CLK), .Q(n10875) );
	dfxtp_1 DFF_44_Q_reg( .D(n4796), .CLK(CLK), .Q(n10790) );
	dfxtp_1 DFF_233_Q_reg( .D(n4936), .CLK(CLK), .Q(n10672) );
	dfxtp_1 DFF_931_Q_reg( .D(n5435), .CLK(CLK), .Q(n10673) );
	dfxtp_1 DFF_538_Q_reg( .D(n4567), .CLK(CLK), .Q(n10379) );
	dfxtp_1 DFF_1005_Q_reg( .D(n4561), .CLK(CLK), .Q(n10374) );
	dfxtp_1 DFF_198_Q_reg( .D(n4560), .CLK(CLK), .Q(n10373) );
	dfxtp_1 DFF_923_Q_reg( .D(n5428), .CLK(CLK), .Q(n10800) );
	dfxtp_1 DFF_307_Q_reg( .D(n4998), .CLK(CLK), .Q(n10789) );
	dfxtp_1 DFF_398_Q_reg( .D(n5061), .CLK(CLK), .Q(n10774) );
	dfxtp_1 DFF_172_Q_reg( .D(n4892), .CLK(CLK), .Q(n10779) );
	dfxtp_1 DFF_1280_Q_reg( .D(n5694), .CLK(CLK), .Q(n10835) );
	dfxtp_1 DFF_92_Q_reg( .D(n4835), .CLK(CLK), .Q(n10753) );
	dfxtp_1 DFF_187_Q_reg( .D(n4902), .CLK(CLK), .Q(n10796) );
	dfxtp_1 DFF_470_Q_reg( .D(n5114), .CLK(CLK), .Q(n10844) );
	dfxtp_1 DFF_534_Q_reg( .D(n5155), .CLK(CLK), .Q(n10843) );
	dfxtp_1 DFF_1104_Q_reg( .D(n5561), .CLK(CLK), .Q(n10735) );
	dfxtp_1 DFF_946_Q_reg( .D(n5444), .CLK(CLK), .Q(n10846) );
	dfxtp_1 DFF_811_Q_reg( .D(n5348), .CLK(CLK), .Q(n10736) );
	dfxtp_1 DFF_164_Q_reg( .D(n4886), .CLK(CLK), .Q(n10586) );
	dfxtp_1 DFF_1036_Q_reg( .D(n5512), .CLK(CLK), .Q(n10848) );
	dfxtp_1 DFF_770_Q_reg( .D(n5317), .CLK(CLK), .Q(n10516) );
	dfxtp_1 DFF_277_Q_reg( .D(n4972), .CLK(CLK), .Q(n10894) );
	dfxtp_1 DFF_453_Q_reg( .D(n5101), .CLK(CLK), .Q(n10591) );
	dfxtp_1 DFF_316_Q_reg( .D(n5005), .CLK(CLK), .Q(n10303) );
	dfxtp_1 DFF_614_Q_reg( .D(n5208), .CLK(CLK), .Q(n10893) );
	dfxtp_1 DFF_1198_Q_reg( .D(n5631), .CLK(CLK), .Q(n10661) );
	dfxtp_1 DFF_1314_Q_reg( .D(n5719), .CLK(CLK), .Q(n10939) );
	dfxtp_1 DFF_932_Q_reg( .D(n5436), .CLK(CLK), .Q(n10938) );
	dfxtp_1 DFF_425_Q_reg( .D(n5080), .CLK(CLK), .Q(n10580) );
	dfxtp_1 DFF_487_Q_reg( .D(n5125), .CLK(CLK), .Q(n10579) );
	dfxtp_1 DFF_570_Q_reg( .D(n5176), .CLK(CLK), .Q(n10582) );
	dfxtp_1 DFF_1240_Q_reg( .D(n5664), .CLK(CLK), .Q(n10581) );
	dfxtp_1 DFF_1202_Q_reg( .D(n5635), .CLK(CLK), .Q(n10584) );
	dfxtp_1 DFF_862_Q_reg( .D(n5381), .CLK(CLK), .Q(n10583) );
	dfxtp_1 DFF_984_Q_reg( .D(n5473), .CLK(CLK), .Q(n10585) );
	dfxtp_1 DFF_1393_Q_reg( .D(n5776), .CLK(CLK), .Q(n10294) );
	dfxtp_1 DFF_1410_Q_reg( .D(n5791), .CLK(CLK), .Q(n10842) );
	dfxtp_1 DFF_1317_Q_reg( .D(n5721), .CLK(CLK), .Q(n10816) );
	dfxtp_1 DFF_1255_Q_reg( .D(n5676), .CLK(CLK), .Q(n10777) );
	dfxtp_1 DFF_464_Q_reg( .D(n5110), .CLK(CLK), .Q(n10751) );
	dfxtp_1 DFF_1307_Q_reg( .D(n5714), .CLK(CLK), .Q(n10764) );
	dfxtp_1 DFF_1406_Q_reg( .D(n5787), .CLK(CLK), .Q(n10803) );
	dfxtp_1 DFF_599_Q_reg( .D(n4563), .CLK(CLK), .Q(n10376) );
	dfxtp_1 DFF_590_Q_reg( .D(n5192), .CLK(CLK), .Q(n10815) );
	dfxtp_1 DFF_227_Q_reg( .D(n4931), .CLK(CLK), .Q(n10826) );
	dfxtp_1 DFF_1263_Q_reg( .D(n5681), .CLK(CLK), .Q(n10841) );
	dfxtp_1 DFF_957_Q_reg( .D(n5455), .CLK(CLK), .Q(n10748) );
	dfxtp_1 DFF_1264_Q_reg( .D(n5682), .CLK(CLK), .Q(n10805) );
	dfxtp_1 DFF_471_Q_reg( .D(n5115), .CLK(CLK), .Q(n10770) );
	dfxtp_1 DFF_378_Q_reg( .D(n5046), .CLK(CLK), .Q(n10744) );
	dfxtp_1 DFF_102_Q_reg( .D(n4843), .CLK(CLK), .Q(n10822) );
	dfxtp_1 DFF_337_Q_reg( .D(n5018), .CLK(CLK), .Q(n10763) );
	dfxtp_1 DFF_1223_Q_reg( .D(n5652), .CLK(CLK), .Q(n10847) );
	dfxtp_1 DFF_1181_Q_reg( .D(n5618), .CLK(CLK), .Q(n10165) );
	dfxtp_1 DFF_600_Q_reg( .D(n4628), .CLK(CLK), .Q(g13259) );
	dfxtp_1 DFF_363_Q_reg( .D(n5037), .CLK(CLK), .Q(n10446) );
	dfxtp_1 DFF_327_Q_reg( .D(n4638), .CLK(CLK), .Q(g13272) );
	dfxtp_1 DFF_1313_Q_reg( .D(n5718), .CLK(CLK), .Q(n10445) );
	dfxtp_1 DFF_579_Q_reg( .D(n5183), .CLK(CLK), .Q(n10762) );
	dfxtp_1 DFF_1378_Q_reg( .D(n5764), .CLK(CLK), .Q(n10840) );
	dfxtp_1 DFF_1291_Q_reg( .D(n5703), .CLK(CLK), .Q(n10773) );
	dfxtp_1 DFF_729_Q_reg( .D(n5287), .CLK(CLK), .Q(n10836) );
	dfxtp_1 DFF_312_Q_reg( .D(n5002), .CLK(CLK), .Q(n10804) );
	dfxtp_1 DFF_19_Q_reg( .D(n4775), .CLK(CLK), .Q(n10821) );
	dfxtp_1 DFF_945_Q_reg( .D(n5443), .CLK(CLK), .Q(n10752) );
	dfxtp_1 DFF_484_Q_reg( .D(n5123), .CLK(CLK), .Q(n10758) );
	dfxtp_1 DFF_937_Q_reg( .D(n4692), .CLK(CLK), .Q(g19357) );
	dfxtp_1 DFF_1190_Q_reg( .D(n22), .CLK(CLK), .Q(n10436) );
	dfxtp_1 DFF_447_Q_reg( .D(n5096), .CLK(CLK), .Q(n10300) );
	dfxtp_1 DFF_1207_Q_reg( .D(n4689), .CLK(CLK), .Q(g19334) );
	dfxtp_1 DFF_1192_Q_reg( .D(n5626), .CLK(CLK), .Q(n10558) );
	dfxtp_1 DFF_361_Q_reg( .D(n5035), .CLK(CLK), .Q(n10212) );
	dfxtp_1 DFF_716_Q_reg( .D(n5275), .CLK(CLK), .Q(n10865) );
	dfxtp_1 DFF_980_Q_reg( .D(n5470), .CLK(CLK), .Q(n10460) );
	dfxtp_1 DFF_373_Q_reg( .D(n5042), .CLK(CLK), .Q(n10919) );
	dfxtp_1 DFF_763_Q_reg( .D(n5312), .CLK(CLK), .Q(n10845) );
	dfxtp_1 DFF_1057_Q_reg( .D(n5528), .CLK(CLK), .Q(n10471) );
	dfxtp_1 DFF_375_Q_reg( .D(n5044), .CLK(CLK), .Q(n10470) );
	dfxtp_1 DFF_202_Q_reg( .D(n4913), .CLK(CLK), .Q(n10874) );
	dfxtp_1 DFF_899_Q_reg( .D(n5411), .CLK(CLK), .Q(n10438) );
	dfxtp_1 DFF_1329_Q_reg( .D(n4693), .CLK(CLK), .Q(g26885) );
	dfxtp_1 DFF_843_Q_reg( .D(n5367), .CLK(CLK), .Q(n10917) );
	dfxtp_1 DFF_840_Q_reg( .D(n5364), .CLK(CLK), .Q(n10420) );
	dfxtp_1 DFF_39_Q_reg( .D(n4792), .CLK(CLK), .Q(n10419) );
	dfxtp_1 DFF_347_Q_reg( .D(n5026), .CLK(CLK), .Q(n10418) );
	dfxtp_1 DFF_1285_Q_reg( .D(n5699), .CLK(CLK), .Q(n10417) );
	dfxtp_1 DFF_731_Q_reg( .D(n5289), .CLK(CLK), .Q(n10415) );
	dfxtp_1 DFF_1188_Q_reg( .D(n5623), .CLK(CLK), .Q(n10414) );
	dfxtp_1 DFF_683_Q_reg( .D(n5252), .CLK(CLK), .Q(n10413) );
	dfxtp_1 DFF_1349_Q_reg( .D(n5743), .CLK(CLK), .Q(n10937) );
	dfxtp_1 DFF_1341_Q_reg( .D(n5736), .CLK(CLK), .Q(n10298) );
	dfxtp_1 DFF_718_Q_reg( .D(n5277), .CLK(CLK), .Q(n10353) );
	dfxtp_1 DFF_722_Q_reg( .D(n5281), .CLK(CLK), .Q(n10918) );
	dfxtp_1 DFF_531_Q_reg( .D(n5152), .CLK(CLK), .Q(n10444) );
	dfxtp_1 DFF_1373_Q_reg( .D(n5761), .CLK(CLK), .Q(n10189) );
	dfxtp_1 DFF_43_Q_reg( .D(n4795), .CLK(CLK), .Q(n10668) );
	dfxtp_1 DFF_711_Q_reg( .D(n4675), .CLK(CLK), .Q(g17291) );
	dfxtp_1 DFF_422_Q_reg( .D(n4672), .CLK(CLK), .Q(g17320) );
	dfxtp_1 DFF_1340_Q_reg( .D(n5735), .CLK(CLK), .Q(n10466) );
	dfxtp_1 DFF_643_Q_reg( .D(n4673), .CLK(CLK), .Q(g17316) );
	dfxtp_1 DFF_146_Q_reg( .D(n4674), .CLK(CLK), .Q(g17404) );
	dfxtp_1 DFF_1267_Q_reg( .D(n5684), .CLK(CLK), .Q(n10631) );
	dfxtp_1 DFF_1369_Q_reg( .D(n5757), .CLK(CLK), .Q(n10636) );
	dfxtp_1 DFF_481_Q_reg( .D(n64), .CLK(CLK), .Q(n10469) );
	dfxtp_1 DFF_1374_Q_reg( .D(n4559), .CLK(CLK), .Q(n10255) );
	dfxtp_1 DFF_261_Q_reg( .D(n4961), .CLK(CLK), .Q(n10715) );
	dfxtp_1 DFF_870_Q_reg( .D(n5388), .CLK(CLK), .Q(n10521) );
	dfxtp_1 DFF_1078_Q_reg( .D(n4757), .CLK(CLK), .Q(g20557) );
	dfxtp_1 DFF_1251_Q_reg( .D(n5672), .CLK(CLK), .Q(n10916) );
	dfxtp_1 DFF_549_Q_reg( .D(n4681), .CLK(CLK), .Q(g4467) );
	dfxtp_1 DFF_1235_Q_reg( .D(n5661), .CLK(CLK), .Q(n10390) );
	dfxtp_1 DFF_1090_Q_reg( .D(n5551), .CLK(CLK), .Q(n10394) );
	dfxtp_1 DFF_896_Q_reg( .D(n5409), .CLK(CLK), .Q(n10400) );
	dfxtp_1 DFF_409_Q_reg( .D(n5069), .CLK(CLK), .Q(n10561) );
	dfxtp_1 DFF_303_Q_reg( .D(n4995), .CLK(CLK), .Q(n10568) );
	dfxtp_1 DFF_431_Q_reg( .D(n5083), .CLK(CLK), .Q(n10567) );
	dfxtp_1 DFF_1008_Q_reg( .D(n5490), .CLK(CLK), .Q(n10703) );
	dfxtp_1 DFF_885_Q_reg( .D(n4690), .CLK(CLK), .Q(g8870) );
	dfxtp_1 DFF_112_Q_reg( .D(n4851), .CLK(CLK), .Q(n10439) );
	dfxtp_1 DFF_162_Q_reg( .D(n4885), .CLK(CLK), .Q(n10396) );
	dfxtp_1 DFF_874_Q_reg( .D(n5390), .CLK(CLK), .Q(n10401) );
	dfxtp_1 DFF_119_Q_reg( .D(n4856), .CLK(CLK), .Q(n10383) );
	dfxtp_1 DFF_149_Q_reg( .D(n4875), .CLK(CLK), .Q(n10410) );
	dfxtp_1 DFF_913_Q_reg( .D(n5420), .CLK(CLK), .Q(n10409) );
	dfxtp_1 DFF_1252_Q_reg( .D(n5673), .CLK(CLK), .Q(n10368) );
	dfxtp_1 DFF_533_Q_reg( .D(n5154), .CLK(CLK), .Q(n10433) );
	dfxtp_1 DFF_393_Q_reg( .D(n5057), .CLK(CLK), .Q(n10155) );
	dfxtp_1 DFF_104_Q_reg( .D(n4845), .CLK(CLK), .Q(n10154) );
	dfxtp_1 DFF_473_Q_reg( .D(n5117), .CLK(CLK), .Q(n10157) );
	dfxtp_1 DFF_245_Q_reg( .D(n4947), .CLK(CLK), .Q(n10158) );
	dfxtp_1 DFF_1122_Q_reg( .D(n4659), .CLK(CLK), .Q(g17400) );
	dfxtp_1 DFF_1110_Q_reg( .D(n4658), .CLK(CLK), .Q(g17423) );
	dfxtp_1 DFF_678_Q_reg( .D(n4683), .CLK(CLK), .Q(g9497) );
	dfxtp_1 DFF_545_Q_reg( .D(n4680), .CLK(CLK), .Q(g9553) );
	dfxtp_1 DFF_489_Q_reg( .D(n4755), .CLK(CLK), .Q(g21292) );
	dfxtp_1 DFF_203_Q_reg( .D(n4660), .CLK(CLK), .Q(g9251) );
	dfxtp_1 DFF_1027_Q_reg( .D(n4657), .CLK(CLK), .Q(g9019) );
	dfxtp_1 DFF_1044_Q_reg( .D(n4752), .CLK(CLK), .Q(g20899) );
	dfxtp_1 DFF_132_Q_reg( .D(n4754), .CLK(CLK), .Q(g21245) );
	dfxtp_1 DFF_358_Q_reg( .D(n5033), .CLK(CLK), .Q(n10341) );
	dfxtp_1 DFF_141_Q_reg( .D(n4564), .CLK(CLK), .Q(g25219) );
	dfxtp_1 DFF_508_Q_reg( .D(n5140), .CLK(CLK), .Q(n10425) );
	dfxtp_1 DFF_201_Q_reg( .D(n4912), .CLK(CLK), .Q(n10434) );
	dfxtp_1 DFF_951_Q_reg( .D(n5449), .CLK(CLK), .Q(n10424) );
	dfxtp_1 DFF_451_Q_reg( .D(n5099), .CLK(CLK), .Q(n10435) );
	dfxtp_1 DFF_985_Q_reg( .D(n5474), .CLK(CLK), .Q(n10931) );
	dfxtp_1 DFF_461_Q_reg( .D(n5107), .CLK(CLK), .Q(n10932) );
	dfxtp_1 DFF_1253_Q_reg( .D(n5674), .CLK(CLK), .Q(n10587) );
	dfxtp_1 DFF_1391_Q_reg( .D(n5775), .CLK(CLK), .Q(n10233) );
	dfxtp_1 DFF_803_Q_reg( .D(n5342), .CLK(CLK), .Q(n10574) );
	dfxtp_1 DFF_90_Q_reg( .D(n4833), .CLK(CLK), .Q(n10215) );
	dfxtp_1 DFF_1371_Q_reg( .D(n5759), .CLK(CLK), .Q(n10214) );
	dfxtp_1 DFF_1389_Q_reg( .D(n5773), .CLK(CLK), .Q(n10670) );
	dfxtp_1 DFF_223_Q_reg( .D(n4928), .CLK(CLK), .Q(n10577) );
	dfxtp_1 DFF_95_Q_reg( .D(n4838), .CLK(CLK), .Q(n10538) );
	dfxtp_1 DFF_820_Q_reg( .D(n5354), .CLK(CLK), .Q(n10477) );
	dfxtp_1 DFF_455_Q_reg( .D(n5103), .CLK(CLK), .Q(n10482) );
	dfxtp_1 DFF_435_Q_reg( .D(n5087), .CLK(CLK), .Q(n10483) );
	dfxtp_1 DFF_795_Q_reg( .D(n5337), .CLK(CLK), .Q(n10479) );
	dfxtp_1 DFF_374_Q_reg( .D(n5043), .CLK(CLK), .Q(n10480) );
	dfxtp_1 DFF_1376_Q_reg( .D(n5763), .CLK(CLK), .Q(n10481) );
	dfxtp_1 DFF_1326_Q_reg( .D(n5726), .CLK(CLK), .Q(n10462) );
	dfxtp_1 DFF_1364_Q_reg( .D(n5753), .CLK(CLK), .Q(n10296) );
	dfxtp_1 DFF_284_Q_reg( .D(n4978), .CLK(CLK), .Q(n10523) );
	dfxtp_1 DFF_1288_Q_reg( .D(n5700), .CLK(CLK), .Q(n10525) );
	dfxtp_1 DFF_5_Q_reg( .D(n4565), .CLK(CLK), .Q(n10377) );
	dfxtp_1 DFF_175_Q_reg( .D(n4895), .CLK(CLK), .Q(n10530) );
	dfxtp_1 DFF_382_Q_reg( .D(n5048), .CLK(CLK), .Q(n10458) );
	dfxtp_1 DFF_1320_Q_reg( .D(n4562), .CLK(CLK), .Q(n10375) );
	dfxtp_1 DFF_1000_Q_reg( .D(n5484), .CLK(CLK), .Q(n10878) );
	dfxtp_1 DFF_757_Q_reg( .D(n5309), .CLK(CLK), .Q(n10622) );
	dfxtp_1 DFF_1270_Q_reg( .D(n5687), .CLK(CLK), .Q(n10280) );
	dfxtp_1 DFF_1306_Q_reg( .D(n5713), .CLK(CLK), .Q(n10503) );
	dfxtp_1 DFF_1360_Q_reg( .D(n5750), .CLK(CLK), .Q(n10504) );
	dfxtp_1 DFF_1035_Q_reg( .D(n5511), .CLK(CLK), .Q(n10702) );
	dfxtp_1 DFF_1117_Q_reg( .D(n5569), .CLK(CLK), .Q(n10571) );
	dfxtp_1 DFF_719_Q_reg( .D(n5278), .CLK(CLK), .Q(n10870) );
	dfxtp_1 DFF_921_Q_reg( .D(n5426), .CLK(CLK), .Q(n10912) );
	dfxtp_1 DFF_169_Q_reg( .D(n4889), .CLK(CLK), .Q(n10909) );
	dfxtp_1 DFF_767_Q_reg( .D(n5314), .CLK(CLK), .Q(n10698) );
	dfxtp_1 DFF_1276_Q_reg( .D(n5691), .CLK(CLK), .Q(n10633) );
	dfxtp_1 DFF_145_Q_reg( .D(n4873), .CLK(CLK), .Q(n10643) );
	dfxtp_1 DFF_1358_Q_reg( .D(n5749), .CLK(CLK), .Q(n10646) );
	dfxtp_1 DFF_897_Q_reg( .D(n5410), .CLK(CLK), .Q(n10640) );
	dfxtp_1 DFF_1215_Q_reg( .D(n5647), .CLK(CLK), .Q(n10642) );
	dfxtp_1 DFF_486_Q_reg( .D(n5124), .CLK(CLK), .Q(n10423) );
	dfxtp_1 DFF_66_Q_reg( .D(n4813), .CLK(CLK), .Q(n10422) );
	dfxtp_1 DFF_793_Q_reg( .D(n5335), .CLK(CLK), .Q(n10171) );
	dfxtp_1 DFF_189_Q_reg( .D(n4903), .CLK(CLK), .Q(n10299) );
	dfxtp_1 DFF_889_Q_reg( .D(n5402), .CLK(CLK), .Q(n10173) );
	dfxtp_1 DFF_297_Q_reg( .D(n4989), .CLK(CLK), .Q(n10172) );
	dfxtp_1 DFF_1236_Q_reg( .D(n5662), .CLK(CLK), .Q(n10174) );
	dfxtp_1 DFF_1344_Q_reg( .D(n5739), .CLK(CLK), .Q(n10301) );
	dfxtp_1 DFF_174_Q_reg( .D(n4894), .CLK(CLK), .Q(n10175) );
	dfxtp_1 DFF_1037_Q_reg( .D(n5513), .CLK(CLK), .Q(n10176) );
	dfxtp_1 DFF_881_Q_reg( .D(n5395), .CLK(CLK), .Q(n10476) );
	dfxtp_1 DFF_844_Q_reg( .D(n5368), .CLK(CLK), .Q(n10307) );
	dfxtp_1 DFF_50_Q_reg( .D(n4800), .CLK(CLK), .Q(n10397) );
	dfxtp_1 DFF_106_Q_reg( .D(n4847), .CLK(CLK), .Q(n10562) );
	dfxtp_1 DFF_700_Q_reg( .D(n5266), .CLK(CLK), .Q(n10408) );
	dfxtp_1 DFF_1339_Q_reg( .D(n5734), .CLK(CLK), .Q(n10564) );
	dfxtp_1 DFF_318_Q_reg( .D(n5006), .CLK(CLK), .Q(n10539) );
	dfxtp_1 DFF_280_Q_reg( .D(n4974), .CLK(CLK), .Q(n10566) );
	dfxtp_1 DFF_954_Q_reg( .D(n5452), .CLK(CLK), .Q(n10565) );
	dfxtp_1 DFF_846_Q_reg( .D(n5370), .CLK(CLK), .Q(n10381) );
	dfxtp_1 DFF_952_Q_reg( .D(n5450), .CLK(CLK), .Q(n10365) );
	dfxtp_1 DFF_242_Q_reg( .D(n4944), .CLK(CLK), .Q(n10576) );
	dfxtp_1 DFF_197_Q_reg( .D(n4910), .CLK(CLK), .Q(n10575) );
	dfxtp_1 DFF_1185_Q_reg( .D(n4652), .CLK(CLK), .Q(g17722) );
	dfxtp_1 DFF_1354_Q_reg( .D(n4655), .CLK(CLK), .Q(g16624) );
	dfxtp_1 DFF_956_Q_reg( .D(n5454), .CLK(CLK), .Q(n10447) );
	dfxtp_1 DFF_1112_Q_reg( .D(n5565), .CLK(CLK), .Q(n10522) );
	dfxtp_1 DFF_1_Q_reg( .D(n4761), .CLK(CLK), .Q(n10524) );
	dfxtp_1 DFF_1149_Q_reg( .D(n5593), .CLK(CLK), .Q(n10879) );
	dfxtp_1 DFF_575_Q_reg( .D(n5180), .CLK(CLK), .Q(n10350) );
	dfxtp_1 DFF_598_Q_reg( .D(n5198), .CLK(CLK), .Q(n10351) );
	dfxtp_1 DFF_271_Q_reg( .D(n4966), .CLK(CLK), .Q(n10352) );
	dfxtp_1 DFF_1068_Q_reg( .D(n5537), .CLK(CLK), .Q(n10349) );
	dfxtp_1 DFF_362_Q_reg( .D(n5036), .CLK(CLK), .Q(n10218) );
	dfxtp_1 DFF_1368_Q_reg( .D(n5756), .CLK(CLK), .Q(n10690) );
	dfxtp_1 DFF_399_Q_reg( .D(n5062), .CLK(CLK), .Q(n10216) );
	dfxtp_1 DFF_283_Q_reg( .D(n4977), .CLK(CLK), .Q(n10557) );
	dfxtp_1 DFF_1039_Q_reg( .D(n5514), .CLK(CLK), .Q(n10556) );
	dfxtp_1 DFF_368_Q_reg( .D(n5040), .CLK(CLK), .Q(n10304) );
	dfxtp_1 DFF_1164_Q_reg( .D(n5604), .CLK(CLK), .Q(n10329) );
	dfxtp_1 DFF_963_Q_reg( .D(n5459), .CLK(CLK), .Q(n10572) );
	dfxtp_1 DFF_852_Q_reg( .D(n5373), .CLK(CLK), .Q(n10437) );
	dfxtp_1 DFF_872_Q_reg( .D(n5389), .CLK(CLK), .Q(n10180) );
	dfxtp_1 DFF_736_Q_reg( .D(n5294), .CLK(CLK), .Q(n10671) );
	dfxtp_1 DFF_664_Q_reg( .D(n4566), .CLK(CLK), .Q(n10378) );
	dfxtp_1 DFF_785_Q_reg( .D(n4650), .CLK(CLK), .Q(g16693) );
	dfxtp_1 DFF_979_Q_reg( .D(n5469), .CLK(CLK), .Q(n10518) );
	dfxtp_1 DFF_1343_Q_reg( .D(n5738), .CLK(CLK), .Q(n10517) );
	dfxtp_1 DFF_1319_Q_reg( .D(n5722), .CLK(CLK), .Q(n10432) );
	dfxtp_1 DFF_133_Q_reg( .D(n4865), .CLK(CLK), .Q(n10472) );
	dfxtp_1 DFF_1347_Q_reg( .D(n5741), .CLK(CLK), .Q(n10327) );
	dfxtp_1 DFF_835_Q_reg( .D(n5360), .CLK(CLK), .Q(n10321) );
	dfxtp_1 DFF_1261_Q_reg( .D(n5680), .CLK(CLK), .Q(n10322) );
	dfxtp_1 DFF_33_Q_reg( .D(n4788), .CLK(CLK), .Q(n10325) );
	dfxtp_1 DFF_768_Q_reg( .D(n5315), .CLK(CLK), .Q(n10319) );
	dfxtp_1 DFF_1075_Q_reg( .D(n5541), .CLK(CLK), .Q(n10324) );
	dfxtp_1 DFF_589_Q_reg( .D(n5191), .CLK(CLK), .Q(n10505) );
	dfxtp_1 DFF_755_Q_reg( .D(n5307), .CLK(CLK), .Q(n10683) );
	dfxtp_1 DFF_929_Q_reg( .D(n5433), .CLK(CLK), .Q(n10928) );
	dfxtp_1 DFF_708_Q_reg( .D(n5271), .CLK(CLK), .Q(n10655) );
	dfxtp_1 DFF_994_Q_reg( .D(n5481), .CLK(CLK), .Q(n10704) );
	dfxtp_1 DFF_733_Q_reg( .D(n5291), .CLK(CLK), .Q(n10716) );
	dfxtp_1 DFF_1382_Q_reg( .D(n5768), .CLK(CLK), .Q(n10913) );
	dfxtp_1 DFF_1290_Q_reg( .D(n5702), .CLK(CLK), .Q(n10910) );
	dfxtp_1 DFF_193_Q_reg( .D(n4906), .CLK(CLK), .Q(n10906) );
	dfxtp_1 DFF_424_Q_reg( .D(n5079), .CLK(CLK), .Q(n10908) );
	dfxtp_1 DFF_1193_Q_reg( .D(n5627), .CLK(CLK), .Q(n10705) );
	dfxtp_1 DFF_452_Q_reg( .D(n5100), .CLK(CLK), .Q(n10278) );
	dfxtp_1 DFF_566_Q_reg( .D(n4648), .CLK(CLK), .Q(g17577) );
	dfxtp_1 DFF_155_Q_reg( .D(n4879), .CLK(CLK), .Q(n10588) );
	dfxtp_1 DFF_222_Q_reg( .D(n4927), .CLK(CLK), .Q(n10657) );
	dfxtp_1 DFF_892_Q_reg( .D(n5405), .CLK(CLK), .Q(n10181) );
	dfxtp_1 DFF_894_Q_reg( .D(n5407), .CLK(CLK), .Q(n10169) );
	dfxtp_1 DFF_139_Q_reg( .D(n4870), .CLK(CLK), .Q(n10366) );
	dfxtp_1 DFF_833_Q_reg( .D(n5359), .CLK(CLK), .Q(n10367) );
	dfxtp_1 DFF_286_Q_reg( .D(n4979), .CLK(CLK), .Q(n10369) );
	dfxtp_1 DFF_1312_Q_reg( .D(n5717), .CLK(CLK), .Q(n10370) );
	dfxtp_1 DFF_195_Q_reg( .D(n4908), .CLK(CLK), .Q(n10590) );
	dfxtp_1 DFF_706_Q_reg( .D(n5269), .CLK(CLK), .Q(n10443) );
	dfxtp_1 DFF_1204_Q_reg( .D(n5637), .CLK(CLK), .Q(n10592) );
	dfxtp_1 DFF_42_Q_reg( .D(n4794), .CLK(CLK), .Q(n10695) );
	dfxtp_1 DFF_847_Q_reg( .D(n5371), .CLK(CLK), .Q(n10347) );
	dfxtp_1 DFF_412_Q_reg( .D(n5072), .CLK(CLK), .Q(n10348) );
	dfxtp_1 DFF_1199_Q_reg( .D(n5632), .CLK(CLK), .Q(n10305) );
	dfxtp_1 DFF_849_Q_reg( .D(n5372), .CLK(CLK), .Q(n10403) );
	dfxtp_1 DFF_440_Q_reg( .D(n5089), .CLK(CLK), .Q(n10660) );
	dfxtp_1 DFF_1016_Q_reg( .D(n5496), .CLK(CLK), .Q(n10364) );
	dfxtp_1 DFF_289_Q_reg( .D(n4982), .CLK(CLK), .Q(n10156) );
	dfxtp_1 DFF_1098_Q_reg( .D(n5559), .CLK(CLK), .Q(n10159) );
	dfxtp_1 DFF_54_Q_reg( .D(n4804), .CLK(CLK), .Q(n10164) );
	dfxtp_1 DFF_1273_Q_reg( .D(n5689), .CLK(CLK), .Q(n10153) );
	dfxtp_1 DFF_717_Q_reg( .D(n5276), .CLK(CLK), .Q(n10237) );
	dfxtp_1 DFF_1361_Q_reg( .D(n5751), .CLK(CLK), .Q(n10356) );
	dfxtp_1 DFF_1019_Q_reg( .D(n5499), .CLK(CLK), .Q(n10520) );
	dfxtp_1 DFF_1094_Q_reg( .D(n5555), .CLK(CLK), .Q(n10441) );
	dfxtp_1 DFF_167_Q_reg( .D(n4888), .CLK(CLK), .Q(n10440) );
	dfxtp_1 DFF_98_Q_reg( .D(n4840), .CLK(CLK), .Q(n10431) );
	dfxtp_1 DFF_182_Q_reg( .D(n4898), .CLK(CLK), .Q(n10430) );
	dfxtp_1 DFF_395_Q_reg( .D(n5058), .CLK(CLK), .Q(n10688) );
	dfxtp_1 DFF_1221_Q_reg( .D(n5651), .CLK(CLK), .Q(n10656) );
	dfxtp_1 DFF_353_Q_reg( .D(n5030), .CLK(CLK), .Q(n10371) );
	dfxtp_1 DFF_828_Q_reg( .D(n4753), .CLK(CLK), .Q(g23683) );
	dfxtp_1 DFF_1404_Q_reg( .D(n5786), .CLK(CLK), .Q(n10416) );
	dfxtp_1 DFF_512_Q_reg( .D(n5144), .CLK(CLK), .Q(n10343) );
	dfxtp_1 DFF_1327_Q_reg( .D(n5727), .CLK(CLK), .Q(n10177) );
	dfxtp_1 DFF_965_Q_reg( .D(n5461), .CLK(CLK), .Q(n10297) );
	dfxtp_1 DFF_661_Q_reg( .D(n5240), .CLK(CLK), .Q(n10385) );
	dfxtp_1 DFF_560_Q_reg( .D(n5171), .CLK(CLK), .Q(n10532) );
	dfxtp_1 DFF_1082_Q_reg( .D(n5544), .CLK(CLK), .Q(n10553) );
	dfxtp_1 DFF_1310_Q_reg( .D(n5715), .CLK(CLK), .Q(n10554) );
	dfxtp_1 DFF_989_Q_reg( .D(n5478), .CLK(CLK), .Q(n10344) );
	dfxtp_1 DFF_812_Q_reg( .D(n5349), .CLK(CLK), .Q(n10398) );
	dfxtp_1 DFF_74_Q_reg( .D(n4821), .CLK(CLK), .Q(n10391) );
	dfxtp_1 DFF_751_Q_reg( .D(n5305), .CLK(CLK), .Q(n10392) );
	dfxtp_1 DFF_772_Q_reg( .D(n5319), .CLK(CLK), .Q(n10345) );
	dfxtp_1 DFF_295_Q_reg( .D(n95), .CLK(CLK), .Q(n10718) );
	dfxtp_1 DFF_372_Q_reg( .D(n75), .CLK(CLK), .Q(n10717) );
	dfxtp_1 DFF_802_Q_reg( .D(n5341), .CLK(CLK), .Q(n10924) );
	dfxtp_1 DFF_293_Q_reg( .D(n4986), .CLK(CLK), .Q(n10484) );
	dfxtp_1 DFF_506_Q_reg( .D(n5138), .CLK(CLK), .Q(n10533) );
	dfxtp_1 DFF_269_Q_reg( .D(n4679), .CLK(CLK), .Q(g8719) );
	dfxtp_1 DFF_331_Q_reg( .D(n36), .CLK(CLK), .Q(n10920) );
	dfxtp_1 DFF_408_Q_reg( .D(n5068), .CLK(CLK), .Q(n10914) );
	dfxtp_1 DFF_863_Q_reg( .D(n5382), .CLK(CLK), .Q(n10531) );
	dfxtp_1 DFF_1115_Q_reg( .D(n5567), .CLK(CLK), .Q(n10478) );
	dfxtp_1 DFF_1020_Q_reg( .D(n5804), .CLK(CLK), .Q(n10552) );
	dfxtp_1 DFF_37_Q_reg( .D(n4790), .CLK(CLK), .Q(n10546) );
	dfxtp_1 DFF_1069_Q_reg( .D(n5538), .CLK(CLK), .Q(n10548) );
	dfxtp_1 DFF_1167_Q_reg( .D(n5606), .CLK(CLK), .Q(n10547) );
	dfxtp_1 DFF_406_Q_reg( .D(n5066), .CLK(CLK), .Q(n10545) );
	dfxtp_1 DFF_402_Q_reg( .D(n5064), .CLK(CLK), .Q(n10287) );
	dfxtp_1 DFF_1127_Q_reg( .D(n5575), .CLK(CLK), .Q(n10286) );
	dfxtp_1 DFF_573_Q_reg( .D(n5178), .CLK(CLK), .Q(n10358) );
	dfxtp_1 DFF_568_Q_reg( .D(n5175), .CLK(CLK), .Q(n10674) );
	dfxtp_1 DFF_1328_Q_reg( .D(n5728), .CLK(CLK), .Q(n10677) );
	dfxtp_1 DFF_804_Q_reg( .D(n5343), .CLK(CLK), .Q(n10676) );
	dfxtp_1 DFF_1129_Q_reg( .D(n5577), .CLK(CLK), .Q(n10678) );
	dfxtp_1 DFF_1281_Q_reg( .D(n5695), .CLK(CLK), .Q(n10681) );
	dfxtp_1 DFF_777_Q_reg( .D(n5323), .CLK(CLK), .Q(n10679) );
	dfxtp_1 DFF_726_Q_reg( .D(n5284), .CLK(CLK), .Q(n10675) );
	dfxtp_1 DFF_977_Q_reg( .D(n5468), .CLK(CLK), .Q(n10680) );
	dfxtp_1 DFF_1053_Q_reg( .D(n5525), .CLK(CLK), .Q(n10339) );
	dfxtp_1 DFF_1136_Q_reg( .D(n5583), .CLK(CLK), .Q(n10306) );
	dfxtp_1 DFF_1323_Q_reg( .D(n5723), .CLK(CLK), .Q(n10285) );
	dfxtp_1 DFF_135_Q_reg( .D(n4867), .CLK(CLK), .Q(n10426) );
	dfxtp_1 DFF_403_Q_reg( .D(n5065), .CLK(CLK), .Q(n10258) );
	dfxtp_1 DFF_1425_Q_reg( .D(n37), .CLK(CLK), .Q(g20049) );
	dfxtp_1 DFF_1045_Q_reg( .D(n5519), .CLK(CLK), .Q(n10354) );
	dfxtp_1 DFF_237_Q_reg( .D(n4939), .CLK(CLK), .Q(n10168) );
	dfxtp_1 DFF_115_Q_reg( .D(n4853), .CLK(CLK), .Q(n10279) );
	dfxtp_1 DFF_1248_Q_reg( .D(n4653), .CLK(CLK), .Q(g17688) );
	dfxtp_1 DFF_797_Q_reg( .D(n4632), .CLK(CLK), .Q(g17739) );
	dfxtp_1 DFF_656_Q_reg( .D(n5235), .CLK(CLK), .Q(n10220) );
	dfxtp_1 DFF_546_Q_reg( .D(n5163), .CLK(CLK), .Q(n10901) );
	dfxtp_1 DFF_1196_Q_reg( .D(n4636), .CLK(CLK), .Q(g17778) );
	dfxtp_1 DFF_927_Q_reg( .D(n4633), .CLK(CLK), .Q(g17674) );
	dfxtp_1 DFF_942_Q_reg( .D(n4634), .CLK(CLK), .Q(g16744) );
	dfxtp_1 DFF_48_Q_reg( .D(n4799), .CLK(CLK), .Q(n10526) );
	dfxtp_1 DFF_760_Q_reg( .D(n5311), .CLK(CLK), .Q(n10185) );
	dfxtp_1 DFF_120_Q_reg( .D(n4857), .CLK(CLK), .Q(n10276) );
	dfxtp_1 DFF_941_Q_reg( .D(n5441), .CLK(CLK), .Q(n10281) );
	dfxtp_1 DFF_953_Q_reg( .D(n5451), .CLK(CLK), .Q(n10402) );
	dfxtp_1 DFF_181_Q_reg( .D(n4644), .CLK(CLK), .Q(g16659) );
	dfxtp_1 DFF_81_Q_reg( .D(n4640), .CLK(CLK), .Q(g16656) );
	dfxtp_1 DFF_966_Q_reg( .D(n5462), .CLK(CLK), .Q(n10528) );
	dfxtp_1 DFF_328_Q_reg( .D(n5014), .CLK(CLK), .Q(n10399) );
	dfxtp_1 DFF_79_Q_reg( .D(n4825), .CLK(CLK), .Q(n10506) );
	dfxtp_1 DFF_734_Q_reg( .D(n5292), .CLK(CLK), .Q(n10272) );
	dfxtp_1 DFF_925_Q_reg( .D(n5430), .CLK(CLK), .Q(n10271) );
	dfxtp_1 DFF_784_Q_reg( .D(n5328), .CLK(CLK), .Q(n10275) );
	dfxtp_1 DFF_1010_Q_reg( .D(n5492), .CLK(CLK), .Q(n10250) );
	dfxtp_1 DFF_1141_Q_reg( .D(n5588), .CLK(CLK), .Q(n10251) );
	dfxtp_1 DFF_305_Q_reg( .D(n4630), .CLK(CLK), .Q(g16775) );
	dfxtp_1 DFF_244_Q_reg( .D(n4946), .CLK(CLK), .Q(n10273) );
	dfxtp_1 DFF_463_Q_reg( .D(n5109), .CLK(CLK), .Q(n10898) );
	dfxtp_1 DFF_58_Q_reg( .D(n4806), .CLK(CLK), .Q(n10902) );
	dfxtp_1 DFF_1066_Q_reg( .D(n5535), .CLK(CLK), .Q(n10899) );
	dfxtp_1 DFF_240_Q_reg( .D(n4942), .CLK(CLK), .Q(n10593) );
	dfxtp_1 DFF_263_Q_reg( .D(n4646), .CLK(CLK), .Q(g17580) );
	dfxtp_1 DFF_906_Q_reg( .D(n4651), .CLK(CLK), .Q(g17519) );
	dfxtp_1 DFF_220_Q_reg( .D(n4645), .CLK(CLK), .Q(g16627) );
	dfxtp_1 DFF_110_Q_reg( .D(n4642), .CLK(CLK), .Q(g17607) );
	dfxtp_1 DFF_315_Q_reg( .D(n4647), .CLK(CLK), .Q(g17649) );
	dfxtp_1 DFF_474_Q_reg( .D(n4631), .CLK(CLK), .Q(g17760) );
	dfxtp_1 DFF_1229_Q_reg( .D(n5656), .CLK(CLK), .Q(n10555) );
	dfxtp_1 DFF_1372_Q_reg( .D(n5760), .CLK(CLK), .Q(n10903) );
	dfxtp_1 DFF_694_Q_reg( .D(n5261), .CLK(CLK), .Q(n10896) );
	dfxtp_1 DFF_170_Q_reg( .D(n4890), .CLK(CLK), .Q(n10897) );
	dfxtp_1 DFF_1346_Q_reg( .D(n5740), .CLK(CLK), .Q(n10900) );
	dfxtp_1 DFF_910_Q_reg( .D(n5417), .CLK(CLK), .Q(n10203) );
	dfxtp_1 DFF_385_Q_reg( .D(n5051), .CLK(CLK), .Q(n10207) );
	dfxtp_1 DFF_20_Q_reg( .D(n4776), .CLK(CLK), .Q(n10206) );
	dfxtp_1 DFF_522_Q_reg( .D(n5148), .CLK(CLK), .Q(n10201) );
	dfxtp_1 DFF_467_Q_reg( .D(n5112), .CLK(CLK), .Q(n10208) );
	dfxtp_1 DFF_1408_Q_reg( .D(n5789), .CLK(CLK), .Q(n10209) );
	dfxtp_1 DFF_737_Q_reg( .D(n4649), .CLK(CLK), .Q(g17646) );
	dfxtp_1 DFF_117_Q_reg( .D(n4629), .CLK(CLK), .Q(g17711) );
	dfxtp_1 DFF_496_Q_reg( .D(n5130), .CLK(CLK), .Q(n10463) );
	dfxtp_1 DFF_673_Q_reg( .D(n5246), .CLK(CLK), .Q(n10465) );
	dfxtp_1 DFF_407_Q_reg( .D(n5067), .CLK(CLK), .Q(n10274) );
	dfxtp_1 DFF_35_Q_reg( .D(n4789), .CLK(CLK), .Q(n10295) );
	dfxtp_1 DFF_410_Q_reg( .D(n5070), .CLK(CLK), .Q(n10270) );
	dfxtp_1 DFF_1293_Q_reg( .D(n4654), .CLK(CLK), .Q(g16603) );
	dfxtp_1 DFF_871_Q_reg( .D(n62), .CLK(CLK), .Q(n10621) );
	dfxtp_1 DFF_118_Q_reg( .D(n4855), .CLK(CLK), .Q(n10192) );
	dfxtp_1 DFF_429_Q_reg( .D(n5082), .CLK(CLK), .Q(n10193) );
	dfxtp_1 DFF_517_Q_reg( .D(n5145), .CLK(CLK), .Q(n10195) );
	dfxtp_1 DFF_536_Q_reg( .D(n5157), .CLK(CLK), .Q(n10196) );
	dfxtp_1 DFF_511_Q_reg( .D(n5143), .CLK(CLK), .Q(n10915) );
	dfxtp_1 DFF_690_Q_reg( .D(n5258), .CLK(CLK), .Q(n10360) );
	dfxtp_1 DFF_1038_Q_reg( .D(n4635), .CLK(CLK), .Q(g16718) );
	dfxtp_1 DFF_445_Q_reg( .D(n5094), .CLK(CLK), .Q(n10382) );
	dfxtp_1 DFF_505_Q_reg( .D(n5137), .CLK(CLK), .Q(n10265) );
	dfxtp_1 DFF_432_Q_reg( .D(n5084), .CLK(CLK), .Q(n10536) );
	dfxtp_1 DFF_1194_Q_reg( .D(n5628), .CLK(CLK), .Q(n10404) );
	dfxtp_1 DFF_646_Q_reg( .D(n5228), .CLK(CLK), .Q(n10266) );
	dfxtp_1 DFF_1379_Q_reg( .D(n5765), .CLK(CLK), .Q(n10361) );
	dfxtp_1 DFF_1275_Q_reg( .D(n4639), .CLK(CLK), .Q(g12923) );
	dfxtp_1 DFF_547_Q_reg( .D(n5164), .CLK(CLK), .Q(n10509) );
	dfxtp_1 DFF_1390_Q_reg( .D(n5774), .CLK(CLK), .Q(n10267) );
	dfxtp_1 DFF_790_Q_reg( .D(n5332), .CLK(CLK), .Q(n10200) );
	dfxtp_1 DFF_1395_Q_reg( .D(n5778), .CLK(CLK), .Q(n10691) );
	dfxtp_1 DFF_232_Q_reg( .D(n4935), .CLK(CLK), .Q(n10693) );
	dfxtp_1 DFF_571_Q_reg( .D(n5177), .CLK(CLK), .Q(n10692) );
	dfxtp_1 DFF_888_Q_reg( .D(n5401), .CLK(CLK), .Q(n10694) );
	dfxtp_1 DFF_446_Q_reg( .D(n5095), .CLK(CLK), .Q(n10697) );
	dfxtp_1 DFF_1243_Q_reg( .D(n5667), .CLK(CLK), .Q(n10696) );
	dfxtp_1 DFF_824_Q_reg( .D(n4661), .CLK(CLK), .Q(g8358) );
	dfxtp_1 DFF_831_Q_reg( .D(n4656), .CLK(CLK), .Q(g8839) );
	dfxtp_1 DFF_60_Q_reg( .D(n4598), .CLK(CLK), .Q(g7946) );
	dfxtp_1 DFF_62_Q_reg( .D(n4809), .CLK(CLK), .Q(n10290) );
	dfxtp_1 DFF_366_Q_reg( .D(n5039), .CLK(CLK), .Q(n10183) );
	dfxtp_1 DFF_1283_Q_reg( .D(n5697), .CLK(CLK), .Q(n10194) );
	dfxtp_1 DFF_724_Q_reg( .D(n5283), .CLK(CLK), .Q(n10380) );
	dfxtp_1 DFF_1103_Q_reg( .D(n5560), .CLK(CLK), .Q(n10405) );
	dfxtp_1 DFF_606_Q_reg( .D(n5203), .CLK(CLK), .Q(n10457) );
	dfxtp_1 DFF_67_Q_reg( .D(n4814), .CLK(CLK), .Q(n10456) );
	dfxtp_1 DFF_1143_Q_reg( .D(n5589), .CLK(CLK), .Q(n10238) );
	dfxtp_1 DFF_819_Q_reg( .D(n4684), .CLK(CLK), .Q(g11349) );
	dfxtp_1 DFF_1001_Q_reg( .D(n4685), .CLK(CLK), .Q(g11418) );
	dfxtp_1 DFF_46_Q_reg( .D(n4677), .CLK(CLK), .Q(g12300) );
	dfxtp_1 DFF_554_Q_reg( .D(n4682), .CLK(CLK), .Q(g12422) );
	dfxtp_1 DFF_1161_Q_reg( .D(n5601), .CLK(CLK), .Q(n10537) );
	dfxtp_1 DFF_660_Q_reg( .D(n5239), .CLK(CLK), .Q(n10515) );
	dfxtp_1 DFF_137_Q_reg( .D(n4869), .CLK(CLK), .Q(n10282) );
	dfxtp_1 DFF_595_Q_reg( .D(n5196), .CLK(CLK), .Q(n10257) );
	dfxtp_1 DFF_1133_Q_reg( .D(n5580), .CLK(CLK), .Q(n10346) );
	dfxtp_1 DFF_853_Q_reg( .D(n5374), .CLK(CLK), .Q(n10245) );
	dfxtp_1 DFF_218_Q_reg( .D(n4925), .CLK(CLK), .Q(n10277) );
	dfxtp_1 DFF_1046_Q_reg( .D(n5520), .CLK(CLK), .Q(n10283) );
	dfxtp_1 DFF_159_Q_reg( .D(n57), .CLK(CLK), .Q(n10922) );
	dfxtp_1 DFF_798_Q_reg( .D(n5339), .CLK(CLK), .Q(n10669) );
	dfxtp_1 DFF_296_Q_reg( .D(n4988), .CLK(CLK), .Q(n10284) );
	dfxtp_1 DFF_774_Q_reg( .D(n5321), .CLK(CLK), .Q(n10256) );
	dfxtp_1 DFF_591_Q_reg( .D(n5193), .CLK(CLK), .Q(n10161) );
	dfxtp_1 DFF_1370_Q_reg( .D(n5758), .CLK(CLK), .Q(n10685) );
	dfxtp_1 DFF_667_Q_reg( .D(n5242), .CLK(CLK), .Q(n10340) );
	dfxtp_1 DFF_1148_Q_reg( .D(n5805), .CLK(CLK), .Q(n10923) );
	dfxtp_1 DFF_214_Q_reg( .D(n4922), .CLK(CLK), .Q(n10248) );
	dfxtp_1 DFF_68_Q_reg( .D(n4815), .CLK(CLK), .Q(n10204) );
	dfxtp_1 DFF_1150_Q_reg( .D(n5594), .CLK(CLK), .Q(n10202) );
	dfxtp_1 DFF_962_Q_reg( .D(n5803), .CLK(CLK), .Q(n10152) );
	dfxtp_1 DFF_1034_Q_reg( .D(n5510), .CLK(CLK), .Q(n10320) );
	dfxtp_1 DFF_1342_Q_reg( .D(n5737), .CLK(CLK), .Q(n10686) );
	dfxtp_1 DFF_400_Q_reg( .D(n5063), .CLK(CLK), .Q(n10502) );
	dfxtp_1 DFF_875_Q_reg( .D(n5391), .CLK(CLK), .Q(n10684) );
	dfxtp_1 DFF_449_Q_reg( .D(n5098), .CLK(CLK), .Q(n10188) );
	dfxtp_1 DFF_878_Q_reg( .D(n5394), .CLK(CLK), .Q(n10191) );
	dfxtp_1 DFF_346_Q_reg( .D(n5025), .CLK(CLK), .Q(n10178) );
	dfxtp_1 DFF_500_Q_reg( .D(n5134), .CLK(CLK), .Q(n10254) );
	dfxtp_1 DFF_671_Q_reg( .D(n5245), .CLK(CLK), .Q(n10252) );
	dfxtp_1 DFF_265_Q_reg( .D(n4963), .CLK(CLK), .Q(n10249) );
	dfxtp_1 DFF_759_Q_reg( .D(n5310), .CLK(CLK), .Q(n10253) );
	dfxtp_1 DFF_622_Q_reg( .D(n5212), .CLK(CLK), .Q(n10293) );
	dfxtp_1 DFF_891_Q_reg( .D(n5404), .CLK(CLK), .Q(n10182) );
	dfxtp_1 DFF_1054_Q_reg( .D(n5526), .CLK(CLK), .Q(n10268) );
	dfxtp_1 DFF_933_Q_reg( .D(n5437), .CLK(CLK), .Q(n10318) );
	dfxtp_1 DFF_1184_Q_reg( .D(n5620), .CLK(CLK), .Q(n10323) );
	dfxtp_1 DFF_713_Q_reg( .D(n5273), .CLK(CLK), .Q(n10247) );
	dfxtp_1 DFF_883_Q_reg( .D(n5397), .CLK(CLK), .Q(n10543) );
	dfxtp_1 DFF_807_Q_reg( .D(n5344), .CLK(CLK), .Q(n10719) );
	dfxtp_1 DFF_886_Q_reg( .D(n5399), .CLK(CLK), .Q(n10259) );
	dfxtp_1 DFF_47_Q_reg( .D(n4798), .CLK(CLK), .Q(n10330) );
	dfxtp_1 DFF_799_Q_reg( .D(n5340), .CLK(CLK), .Q(n10219) );
	dfxtp_1 DFF_1145_Q_reg( .D(n5591), .CLK(CLK), .Q(n10199) );
	dfxtp_1 DFF_675_Q_reg( .D(n4619), .CLK(CLK), .Q(g7916) );
	dfxtp_1 DFF_529_Q_reg( .D(n4624), .CLK(CLK), .Q(g13895) );
	dfxtp_1 DFF_326_Q_reg( .D(n4621), .CLK(CLK), .Q(g14738) );
	dfxtp_1 DFF_635_Q_reg( .D(n5221), .CLK(CLK), .Q(n10198) );
	dfxtp_1 DFF_1065_Q_reg( .D(n5534), .CLK(CLK), .Q(n10151) );
	dfxtp_1 DFF_401_Q_reg( .D(n4622), .CLK(CLK), .Q(g13966) );
	dfxtp_1 DFF_468_Q_reg( .D(n4623), .CLK(CLK), .Q(g13926) );
	dfxtp_1 DFF_669_Q_reg( .D(n5243), .CLK(CLK), .Q(n10406) );
	dfxtp_1 DFF_1173_Q_reg( .D(n5610), .CLK(CLK), .Q(n10160) );
	dfxtp_1 DFF_1324_Q_reg( .D(n5724), .CLK(CLK), .Q(n10362) );
	dfxtp_1 DFF_1335_Q_reg( .D(n4627), .CLK(CLK), .Q(g14694) );
	dfxtp_1 DFF_806_Q_reg( .D(n4626), .CLK(CLK), .Q(g14828) );
	dfxtp_1 DFF_655_Q_reg( .D(n4625), .CLK(CLK), .Q(g14662) );
	dfxtp_1 DFF_188_Q_reg( .D(n4620), .CLK(CLK), .Q(g14779) );
	dfxtp_1 DFF_209_Q_reg( .D(n4917), .CLK(CLK), .Q(n10239) );
	dfxtp_1 DFF_769_Q_reg( .D(n5316), .CLK(CLK), .Q(n10240) );
	dfxtp_1 DFF_272_Q_reg( .D(n4967), .CLK(CLK), .Q(n10243) );
	dfxtp_1 DFF_1413_Q_reg( .D(n5793), .CLK(CLK), .Q(n10241) );
	dfxtp_1 DFF_111_Q_reg( .D(n4850), .CLK(CLK), .Q(n10242) );
	dfxtp_1 DFF_30_Q_reg( .D(n4676), .CLK(CLK), .Q(g12350) );
	dfxtp_1 DFF_1158_Q_reg( .D(n4686), .CLK(CLK), .Q(g12470) );
	dfxtp_1 DFF_165_Q_reg( .D(n4678), .CLK(CLK), .Q(g12238) );
	dfxtp_1 DFF_1420_Q_reg( .D(n4687), .CLK(CLK), .Q(g11388) );
	dfxtp_1 DFF_1232_Q_reg( .D(n5659), .CLK(CLK), .Q(n10921) );
	dfxtp_1 DFF_1084_Q_reg( .D(n5546), .CLK(CLK), .Q(n10246) );
	dfxtp_1 DFF_99_Q_reg( .D(n4841), .CLK(CLK), .Q(n10197) );
	dfxtp_1 DFF_845_Q_reg( .D(n5369), .CLK(CLK), .Q(n10338) );
	dfxtp_1 DFF_551_Q_reg( .D(n5166), .CLK(CLK), .Q(n10342) );
	dfxtp_1 DFF_746_Q_reg( .D(n5300), .CLK(CLK), .Q(n10244) );
	dfxtp_1 DFF_860_Q_reg( .D(n5380), .CLK(CLK), .Q(n10328) );
	dfxtp_1 DFF_948_Q_reg( .D(n5446), .CLK(CLK), .Q(n10508) );
	dfxtp_1 DFF_914_Q_reg( .D(n5421), .CLK(CLK), .Q(n10289) );
	dfxtp_1 DFF_386_Q_reg( .D(n5052), .CLK(CLK), .Q(n10514) );
	dfxtp_1 DFF_1242_Q_reg( .D(n5666), .CLK(CLK), .Q(n10507) );
	dfxtp_1 DFF_18_Q_reg( .D(n4774), .CLK(CLK), .Q(n10264) );
	dfxtp_1 DFF_996_Q_reg( .D(n5483), .CLK(CLK), .Q(n10262) );
	dfxtp_1 DFF_620_Q_reg( .D(n5211), .CLK(CLK), .Q(n10263) );
	dfxtp_1 DFF_339_Q_reg( .D(n4637), .CLK(CLK), .Q(g12919) );
	dfxtp_1 DFF_63_Q_reg( .D(n4810), .CLK(CLK), .Q(n10269) );
	dfxtp_1 DFF_648_Q_reg( .D(n5230), .CLK(CLK), .Q(n10302) );
	dfxtp_1 DFF_771_Q_reg( .D(n5318), .CLK(CLK), .Q(n10459) );
	dfxtp_1 DFF_411_Q_reg( .D(n5071), .CLK(CLK), .Q(n10163) );
	dfxtp_1 DFF_562_Q_reg( .D(n5172), .CLK(CLK), .Q(n10331) );
	dfxtp_1 DFF_1091_Q_reg( .D(n5552), .CLK(CLK), .Q(n10334) );
	dfxtp_1 DFF_103_Q_reg( .D(n4844), .CLK(CLK), .Q(n10336) );
	dfxtp_1 DFF_148_Q_reg( .D(n4874), .CLK(CLK), .Q(n10332) );
	dfxtp_1 DFF_681_Q_reg( .D(n5250), .CLK(CLK), .Q(n10333) );
	dfxtp_1 DFF_1295_Q_reg( .D(n5705), .CLK(CLK), .Q(n10335) );
	dfxtp_1 DFF_794_Q_reg( .D(n5336), .CLK(CLK), .Q(n10292) );
	dfxtp_1 DFF_1375_Q_reg( .D(n5762), .CLK(CLK), .Q(n10337) );
	dfxtp_1 DFF_1233_Q_reg( .D(n5660), .CLK(CLK), .Q(n10260) );
	dfxtp_1 DFF_1047_Q_reg( .D(n5521), .CLK(CLK), .Q(n10261) );
	dfxtp_1 DFF_351_Q_reg( .D(n5029), .CLK(CLK), .Q(n10288) );
	dfxtp_1 DFF_698_Q_reg( .D(n5264), .CLK(CLK), .Q(n10179) );
	dfxtp_1 DFF_990_Q_reg( .D(n5479), .CLK(CLK), .Q(n10326) );
	dfxtp_1 DFF_541_Q_reg( .D(n5159), .CLK(CLK), .Q(n10187) );
	dfxtp_1 DFF_748_Q_reg( .D(n5302), .CLK(CLK), .Q(n10236) );
	dfxtp_1 DFF_1080_Q_reg( .D(n5543), .CLK(CLK), .Q(n10235) );
	inv_2 U6662( .A(1'b1), .Y(g34597) );
	inv_2 U6664( .A(1'b0), .Y(g34240) );
	inv_2 U6666( .A(1'b0), .Y(g34239) );
	inv_2 U6668( .A(1'b0), .Y(g34238) );
	inv_2 U6670( .A(1'b0), .Y(g34237) );
	inv_2 U6672( .A(1'b0), .Y(g34236) );
	inv_2 U6674( .A(1'b0), .Y(g34235) );
	inv_2 U6676( .A(1'b0), .Y(g34234) );
	inv_2 U6678( .A(1'b0), .Y(g34233) );
	inv_2 U6680( .A(1'b0), .Y(g34232) );
	inv_2 U6682( .A(1'b0), .Y(g33950) );
	inv_2 U6684( .A(1'b0), .Y(g33949) );
	inv_2 U6686( .A(1'b0), .Y(g33948) );
	inv_2 U6688( .A(1'b0), .Y(g33947) );
	inv_2 U6690( .A(1'b0), .Y(g33946) );
	inv_2 U6692( .A(1'b0), .Y(g33945) );
	inv_2 U6694( .A(1'b0), .Y(g32454) );
	inv_2 U6696( .A(1'b0), .Y(g32429) );
	inv_2 U6698( .A(1'b0), .Y(g25590) );
	inv_2 U6700( .A(1'b0), .Y(g25589) );
	inv_2 U6702( .A(1'b0), .Y(g25588) );
	inv_2 U6704( .A(1'b0), .Y(g25587) );
	inv_2 U6706( .A(1'b0), .Y(g25586) );
	inv_2 U6708( .A(1'b0), .Y(g25585) );
	inv_2 U6710( .A(1'b0), .Y(g25584) );
	inv_2 U6712( .A(1'b0), .Y(g25583) );
	inv_2 U6714( .A(1'b0), .Y(g25582) );
	inv_2 U6716( .A(1'b0), .Y(g24151) );
	nor2_4 U6718( .A(g35), .B(n6363), .Y(n6437) );
	buf_1 U6719( .A(n6165), .X(n6196) );
	buf_1 U6720( .A(n6165), .X(n6197) );
	buf_1 U6721( .A(n6167), .X(n6203) );
	buf_1 U6722( .A(n6169), .X(n6209) );
	buf_1 U6723( .A(n6169), .X(n6208) );
	buf_1 U6724( .A(n6169), .X(n6210) );
	buf_1 U6725( .A(n6167), .X(n6204) );
	buf_1 U6726( .A(n6168), .X(n6207) );
	buf_1 U6727( .A(n6170), .X(n6211) );
	buf_1 U6728( .A(n6168), .X(n6205) );
	buf_1 U6729( .A(n6168), .X(n6206) );
	inv_2 U6730( .A(n6328), .Y(n6278) );
	buf_1 U6731( .A(n6167), .X(n6202) );
	buf_1 U6732( .A(n6165), .X(n6198) );
	buf_1 U6733( .A(n6170), .X(n6212) );
	buf_1 U6734( .A(n6166), .X(n6199) );
	buf_1 U6735( .A(n6166), .X(n6201) );
	buf_1 U6736( .A(n6166), .X(n6200) );
	inv_2 U6737( .A(n6329), .Y(n6277) );
	inv_2 U6738( .A(n6320), .Y(n6301) );
	inv_2 U6739( .A(n6321), .Y(n6299) );
	inv_2 U6740( .A(n6320), .Y(n6300) );
	buf_1 U6741( .A(n6174), .X(n6225) );
	buf_1 U6742( .A(n6171), .X(n6215) );
	buf_1 U6743( .A(n6172), .X(n6219) );
	buf_1 U6744( .A(n6170), .X(n6213) );
	buf_1 U6745( .A(n6171), .X(n6214) );
	buf_1 U6746( .A(n6171), .X(n6216) );
	buf_1 U6747( .A(n6172), .X(n6217) );
	buf_1 U6748( .A(n6172), .X(n6218) );
	inv_2 U6749( .A(n6318), .Y(n6306) );
	inv_2 U6750( .A(n6321), .Y(n6298) );
	inv_2 U6751( .A(n6318), .Y(n6307) );
	buf_1 U6752( .A(n6173), .X(n6220) );
	inv_2 U6753( .A(n6322), .Y(n6295) );
	inv_2 U6754( .A(n6321), .Y(n6297) );
	inv_2 U6755( .A(n6322), .Y(n6296) );
	buf_1 U6756( .A(n6176), .X(n6230) );
	buf_1 U6757( .A(n6178), .X(n6237) );
	buf_1 U6758( .A(n6178), .X(n6235) );
	buf_1 U6759( .A(n6175), .X(n6227) );
	buf_1 U6760( .A(n6179), .X(n6238) );
	buf_1 U6761( .A(n6177), .X(n6234) );
	buf_1 U6762( .A(n6175), .X(n6228) );
	buf_1 U6763( .A(n6175), .X(n6226) );
	buf_1 U6764( .A(n6179), .X(n6240) );
	buf_1 U6765( .A(n6177), .X(n6233) );
	buf_1 U6766( .A(n6176), .X(n6231) );
	buf_1 U6767( .A(n6176), .X(n6229) );
	buf_1 U6768( .A(n6177), .X(n6232) );
	buf_1 U6769( .A(n6179), .X(n6239) );
	buf_1 U6770( .A(n6178), .X(n6236) );
	inv_2 U6771( .A(n6317), .Y(n6309) );
	inv_2 U6772( .A(n6317), .Y(n6308) );
	buf_1 U6773( .A(n6173), .X(n6222) );
	buf_1 U6774( .A(n6174), .X(n6224) );
	buf_1 U6775( .A(n6173), .X(n6221) );
	buf_1 U6776( .A(n6174), .X(n6223) );
	inv_2 U6777( .A(n6322), .Y(n6294) );
	inv_2 U6778( .A(n6315), .Y(n6314) );
	inv_2 U6779( .A(n6320), .Y(n6302) );
	inv_2 U6780( .A(n6324), .Y(n6291) );
	inv_2 U6781( .A(n6327), .Y(n6281) );
	inv_2 U6782( .A(n6324), .Y(n6290) );
	inv_2 U6783( .A(n6327), .Y(n6283) );
	inv_2 U6784( .A(n6326), .Y(n6286) );
	inv_2 U6785( .A(n6323), .Y(n6292) );
	inv_2 U6786( .A(n6326), .Y(n6285) );
	inv_2 U6787( .A(n6328), .Y(n6280) );
	inv_2 U6788( .A(n6326), .Y(n6284) );
	inv_2 U6789( .A(n6328), .Y(n6279) );
	inv_2 U6790( .A(n6325), .Y(n6289) );
	inv_2 U6791( .A(n6325), .Y(n6287) );
	inv_2 U6792( .A(n6327), .Y(n6282) );
	inv_2 U6793( .A(n6323), .Y(n6293) );
	inv_2 U6794( .A(n6325), .Y(n6288) );
	inv_2 U6795( .A(n6315), .Y(n6313) );
	inv_2 U6796( .A(n6316), .Y(n6312) );
	inv_2 U6797( .A(n6319), .Y(n6303) );
	inv_2 U6798( .A(n6318), .Y(n6305) );
	inv_2 U6799( .A(n6319), .Y(n6304) );
	inv_2 U6800( .A(n6316), .Y(n6310) );
	inv_2 U6801( .A(n6316), .Y(n6311) );
	buf_1 U6802( .A(n6164), .X(n6195) );
	buf_1 U6803( .A(n6164), .X(n6194) );
	buf_1 U6804( .A(n6164), .X(n6193) );
	buf_1 U6805( .A(n6180), .X(n6241) );
	buf_1 U6806( .A(n6180), .X(n6242) );
	buf_1 U6807( .A(n6182), .X(n6247) );
	buf_1 U6808( .A(n6181), .X(n6246) );
	buf_1 U6809( .A(n6180), .X(n6243) );
	buf_1 U6810( .A(n6181), .X(n6245) );
	buf_1 U6811( .A(n6181), .X(n6244) );
	buf_1 U6812( .A(n6267), .X(n6330) );
	buf_1 U6813( .A(n6271), .X(n6341) );
	buf_1 U6814( .A(n6272), .X(n6344) );
	buf_1 U6815( .A(n6271), .X(n6343) );
	buf_1 U6816( .A(n6271), .X(n6342) );
	buf_1 U6817( .A(n6267), .X(n6331) );
	buf_1 U6818( .A(n6268), .X(n6334) );
	buf_1 U6819( .A(n6269), .X(n6336) );
	buf_1 U6820( .A(n6269), .X(n6335) );
	buf_1 U6821( .A(n6268), .X(n6333) );
	buf_1 U6822( .A(n6268), .X(n6332) );
	buf_1 U6823( .A(n6269), .X(n6337) );
	buf_1 U6824( .A(n6267), .X(n6329) );
	buf_1 U6825( .A(n6272), .X(n6345) );
	buf_1 U6826( .A(n6266), .X(n6326) );
	buf_1 U6827( .A(n6266), .X(n6328) );
	buf_1 U6828( .A(n6265), .X(n6324) );
	buf_1 U6829( .A(n6266), .X(n6327) );
	buf_1 U6830( .A(n6264), .X(n6323) );
	buf_1 U6831( .A(n6264), .X(n6321) );
	buf_1 U6832( .A(n6265), .X(n6325) );
	buf_1 U6833( .A(n6263), .X(n6318) );
	buf_1 U6834( .A(n6262), .X(n6315) );
	buf_1 U6835( .A(n6262), .X(n6317) );
	buf_1 U6836( .A(n6262), .X(n6316) );
	buf_1 U6837( .A(n6264), .X(n6322) );
	buf_1 U6838( .A(n6263), .X(n6320) );
	buf_1 U6839( .A(n6263), .X(n6319) );
	buf_1 U6840( .A(n6270), .X(n6338) );
	buf_1 U6841( .A(n6270), .X(n6339) );
	buf_1 U6842( .A(n6182), .X(n6248) );
	buf_1 U6843( .A(n6270), .X(n6340) );
	buf_1 U6844( .A(n6272), .X(n6346) );
	buf_1 U6845( .A(n6186), .X(n6173) );
	buf_1 U6846( .A(n6185), .X(n6174) );
	buf_1 U6847( .A(n6187), .X(n6169) );
	buf_1 U6848( .A(n6185), .X(n6175) );
	buf_1 U6849( .A(n6186), .X(n6171) );
	buf_1 U6850( .A(n6185), .X(n6176) );
	buf_1 U6851( .A(n6188), .X(n6167) );
	buf_1 U6852( .A(n6186), .X(n6172) );
	buf_1 U6853( .A(n6184), .X(n6177) );
	buf_1 U6854( .A(n6187), .X(n6170) );
	buf_1 U6855( .A(n6188), .X(n6166) );
	buf_1 U6856( .A(n6187), .X(n6168) );
	buf_1 U6857( .A(n6184), .X(n6179) );
	buf_1 U6858( .A(n6184), .X(n6178) );
	buf_1 U6859( .A(n6188), .X(n6165) );
	buf_1 U6860( .A(n6274), .X(n6268) );
	buf_1 U6861( .A(n6191), .X(n6185) );
	buf_1 U6862( .A(n6275), .X(n6266) );
	buf_1 U6863( .A(n6275), .X(n6264) );
	buf_1 U6864( .A(n6275), .X(n6265) );
	buf_1 U6865( .A(n6274), .X(n6269) );
	buf_1 U6866( .A(n6273), .X(n6272) );
	buf_1 U6867( .A(n6273), .X(n6271) );
	buf_1 U6868( .A(n6274), .X(n6267) );
	buf_1 U6869( .A(n6191), .X(n6186) );
	buf_1 U6870( .A(n6276), .X(n6262) );
	buf_1 U6871( .A(n6190), .X(n6187) );
	buf_1 U6872( .A(n6273), .X(n6270) );
	buf_1 U6873( .A(n6191), .X(n6184) );
	buf_1 U6874( .A(n6190), .X(n6188) );
	buf_1 U6875( .A(n6276), .X(n6263) );
	buf_1 U6876( .A(n6183), .X(n6180) );
	buf_1 U6877( .A(n6183), .X(n6181) );
	buf_1 U6878( .A(n6189), .X(n6164) );
	buf_1 U6879( .A(n6190), .X(n6189) );
	buf_1 U6880( .A(n6183), .X(n6182) );
	buf_1 U6881( .A(n6426), .X(n6249) );
	buf_1 U6882( .A(n6426), .X(n6252) );
	buf_1 U6883( .A(n6426), .X(n6251) );
	buf_1 U6884( .A(n6426), .X(n6250) );
	buf_1 U6885( .A(n6426), .X(n6259) );
	buf_1 U6886( .A(n6426), .X(n6253) );
	buf_1 U6887( .A(n6426), .X(n6260) );
	buf_1 U6888( .A(n6426), .X(n6258) );
	buf_1 U6889( .A(n6426), .X(n6257) );
	buf_1 U6890( .A(n6426), .X(n6256) );
	buf_1 U6891( .A(n6426), .X(n6254) );
	buf_1 U6892( .A(n6426), .X(n6255) );
	buf_1 U6893( .A(n6426), .X(n6261) );
	buf_1 U6894( .A(n6192), .X(n6183) );
	buf_1 U6895( .A(n6390), .X(n6192) );
	buf_1 U6896( .A(n6457), .X(n6275) );
	buf_1 U6897( .A(n6457), .X(n6274) );
	buf_1 U6898( .A(n6390), .X(n6191) );
	buf_1 U6899( .A(n6457), .X(n6273) );
	buf_1 U6900( .A(n6390), .X(n6190) );
	buf_1 U6901( .A(n6457), .X(n6276) );
	inv_2 U6902( .A(n6373), .Y(n6349) );
	inv_2 U6903( .A(n6373), .Y(n6348) );
	inv_2 U6904( .A(n6370), .Y(n6350) );
	inv_2 U6905( .A(n6373), .Y(n6347) );
	inv_2 U6906( .A(n6370), .Y(n6368) );
	inv_2 U6907( .A(n6371), .Y(n6364) );
	inv_2 U6908( .A(n6371), .Y(n6365) );
	inv_2 U6909( .A(n6371), .Y(n6366) );
	inv_2 U6910( .A(n6372), .Y(n6363) );
	inv_2 U6911( .A(n6371), .Y(n6351) );
	inv_2 U6912( .A(n6370), .Y(n6367) );
	inv_2 U6913( .A(n6372), .Y(n6362) );
	inv_2 U6914( .A(n6372), .Y(n6361) );
	inv_2 U6915( .A(n6372), .Y(n6352) );
	inv_2 U6916( .A(n6370), .Y(n6359) );
	inv_2 U6917( .A(n6371), .Y(n6358) );
	inv_2 U6918( .A(n6385), .Y(n6357) );
	inv_2 U6919( .A(n6384), .Y(n6355) );
	inv_2 U6920( .A(n6387), .Y(n6354) );
	inv_2 U6921( .A(n6386), .Y(n6356) );
	inv_2 U6922( .A(n6372), .Y(n6353) );
	inv_2 U6923( .A(n6373), .Y(n6360) );
	inv_2 U6924( .A(n6370), .Y(n6369) );
	inv_2 U6925( .A(RST), .Y(n6377) );
	inv_2 U6926( .A(RST), .Y(n6374) );
	inv_2 U6927( .A(RST), .Y(n6376) );
	inv_2 U6928( .A(RST), .Y(n6375) );
	inv_2 U6929( .A(RST), .Y(n6382) );
	inv_2 U6930( .A(RST), .Y(n6383) );
	inv_2 U6931( .A(RST), .Y(n6378) );
	inv_2 U6932( .A(RST), .Y(n6379) );
	inv_2 U6933( .A(RST), .Y(n6380) );
	inv_2 U6934( .A(RST), .Y(n6381) );
	inv_2 U6935( .A(RST), .Y(n6373) );
	inv_2 U6936( .A(RST), .Y(n6371) );
	inv_2 U6937( .A(RST), .Y(n6370) );
	inv_2 U6938( .A(RST), .Y(n6372) );
	inv_2 U6939( .A(RST), .Y(n6387) );
	inv_2 U6940( .A(RST), .Y(n6385) );
	inv_2 U6941( .A(RST), .Y(n6384) );
	inv_2 U6942( .A(RST), .Y(n6386) );
	buf_1 U6943( .A(g34839), .X(g34956) );
	buf_1 U6944( .A(g33894), .X(g34788) );
	buf_1 U6945( .A(g31521), .X(g34435) );
	buf_1 U6946( .A(g26801), .X(g32975) );
	buf_1 U6947( .A(g25167), .X(g31863) );
	buf_1 U6948( .A(g25259), .X(g31862) );
	buf_1 U6949( .A(g25219), .X(g31861) );
	buf_1 U6950( .A(g31665), .X(g34437) );
	buf_1 U6951( .A(g31656), .X(g34436) );
	buf_1 U6952( .A(g23683), .X(g30332) );
	buf_1 U6953( .A(g23759), .X(g30331) );
	buf_1 U6954( .A(g23002), .X(g30327) );
	buf_1 U6955( .A(g21292), .X(g29221) );
	buf_1 U6956( .A(g21245), .X(g29220) );
	buf_1 U6957( .A(g20654), .X(g29219) );
	buf_1 U6958( .A(g21270), .X(g29217) );
	buf_1 U6959( .A(g21176), .X(g29216) );
	buf_1 U6960( .A(g20901), .X(g29215) );
	buf_1 U6961( .A(g20652), .X(g29214) );
	buf_1 U6962( .A(g20557), .X(g29213) );
	buf_1 U6963( .A(g20899), .X(g29212) );
	buf_1 U6964( .A(g20763), .X(g29211) );
	buf_1 U6965( .A(g20049), .X(g29210) );
	buf_1 U6966( .A(g28753), .X(g33959) );
	buf_1 U6967( .A(g27831), .X(g33533) );
	buf_1 U6968( .A(g25114), .X(g31860) );
	buf_1 U6969( .A(g44), .X(g24185) );
	buf_1 U6970( .A(g135), .X(g24184) );
	buf_1 U6971( .A(g134), .X(g24183) );
	buf_1 U6972( .A(g127), .X(g24182) );
	buf_1 U6973( .A(g126), .X(g24181) );
	buf_1 U6974( .A(g125), .X(g24180) );
	buf_1 U6975( .A(g124), .X(g24179) );
	buf_1 U6976( .A(g120), .X(g24178) );
	buf_1 U6977( .A(g116), .X(g24177) );
	buf_1 U6978( .A(g115), .X(g24176) );
	buf_1 U6979( .A(g114), .X(g24175) );
	buf_1 U6980( .A(g113), .X(g24174) );
	buf_1 U6981( .A(g100), .X(g24173) );
	buf_1 U6982( .A(g99), .X(g24172) );
	buf_1 U6983( .A(g92), .X(g24171) );
	buf_1 U6984( .A(g91), .X(g24170) );
	buf_1 U6985( .A(g90), .X(g24169) );
	buf_1 U6986( .A(g84), .X(g24168) );
	buf_1 U6987( .A(g73), .X(g24167) );
	buf_1 U6988( .A(g72), .X(g24166) );
	buf_1 U6989( .A(g64), .X(g24165) );
	buf_1 U6990( .A(g57), .X(g24164) );
	buf_1 U6991( .A(g56), .X(g24163) );
	buf_1 U6992( .A(g54), .X(g24162) );
	buf_1 U6993( .A(g53), .X(g24161) );
	buf_1 U6994( .A(g23652), .X(g30330) );
	buf_1 U6995( .A(g23612), .X(g30329) );
	buf_1 U6996( .A(g36), .X(g21698) );
	buf_1 U6997( .A(g18881), .X(g29218) );
	buf_1 U6998( .A(g6746), .X(g18101) );
	buf_1 U6999( .A(g6751), .X(g18100) );
	buf_1 U7000( .A(g6745), .X(g18099) );
	buf_1 U7001( .A(g6744), .X(g18098) );
	buf_1 U7002( .A(g6747), .X(g18097) );
	buf_1 U7003( .A(g6750), .X(g18096) );
	buf_1 U7004( .A(g6749), .X(g18095) );
	buf_1 U7005( .A(g6748), .X(g18094) );
	buf_1 U7006( .A(g6753), .X(g18092) );
	a21oi_1 U7007( .A1(n6388), .A2(n6389), .B1(n6308), .Y(n5805) );
	xnor2_1 U7008( .A(n10923), .B(g7946), .Y(n6388) );
	o21ai_0 U7009( .A1(n6233), .A2(n6391), .B1(n6392), .Y(n5804) );
	mux2i_1 U7010( .A0(n6393), .A1(n6394), .S(n6395), .Y(n6392) );
	nor2_1 U7011( .A(n6396), .B(n6397), .Y(n6394) );
	nor3_1 U7012( .A(n6398), .B(n10552), .C(n6368), .Y(n6393) );
	o221ai_1 U7013( .A1(n6212), .A2(n6399), .B1(n10152), .B2(n6312), .C1(n6400), .Y(n5803) );
	inv_1 U7014( .A(n10917), .Y(n6399) );
	or3_1 U7015( .A(n6401), .B(n6402), .C(n6403), .X(n5802) );
	o22ai_1 U7016( .A1(n6404), .A2(n6405), .B1(n6196), .B2(n6406), .Y(n6403) );
	a21oi_1 U7017( .A1(n6407), .A2(n6408), .B1(n6307), .Y(n6402) );
	nor3_1 U7018( .A(n6409), .B(g7916), .C(n6368), .Y(n6401) );
	o21ai_0 U7019( .A1(n6227), .A2(n6410), .B1(n6411), .Y(n5801) );
	mux2i_1 U7020( .A0(n6412), .A1(n6413), .S(n6414), .Y(n6411) );
	nor2_1 U7021( .A(n6415), .B(n6299), .Y(n6413) );
	and2_0 U7022( .A(n6415), .B(n6416), .X(n6412) );
	mux2i_1 U7023( .A0(n6417), .A1(n6418), .S(n6410), .Y(n6415) );
	nor2_1 U7024( .A(n10177), .B(n6419), .Y(n6418) );
	nor2_1 U7025( .A(n6420), .B(n6421), .Y(n6417) );
	nor2_1 U7026( .A(n6359), .B(n6422), .Y(n5800) );
	o21ai_0 U7027( .A1(n6228), .A2(n6423), .B1(n6424), .Y(n5799) );
	a22oi_1 U7028( .A1(n10784), .A2(n6425), .B1(n6249), .B2(n6427), .Y(n6424) );
	o21ai_0 U7029( .A1(n6229), .A2(n6022), .B1(n6428), .Y(n5798) );
	mux2i_1 U7030( .A0(n6429), .A1(n6430), .S(n6431), .Y(n6428) );
	nor2_1 U7031( .A(n10263), .B(n6432), .Y(n6431) );
	nor2_1 U7032( .A(n6277), .B(n5998), .Y(n6429) );
	o32ai_1 U7033( .A1(n5908), .A2(n6433), .A3(n6313), .B1(n6434), .B2(n6435), .Y(n5797) );
	nor2_1 U7034( .A(n6436), .B(n6437), .Y(n6434) );
	nor4_1 U7035( .A(n11959), .B(n6367), .C(n6438), .D(n6439), .Y(n6436) );
	a21oi_1 U7036( .A1(n6440), .A2(n6435), .B1(n6439), .Y(n6433) );
	o21ai_0 U7037( .A1(n6441), .A2(n6096), .B1(n6442), .Y(n5796) );
	mux2i_1 U7038( .A0(n6443), .A1(n6444), .S(n6445), .Y(n6442) );
	nor2_1 U7039( .A(n10325), .B(n6446), .Y(n6444) );
	nand2_1 U7040( .A(n6221), .B(n6447), .Y(n6443) );
	o22ai_1 U7041( .A1(n6210), .A2(n6448), .B1(n6449), .B2(n6295), .Y(n5795) );
	nor2_1 U7042( .A(g4242), .B(n10453), .Y(n6449) );
	inv_1 U7043( .A(n10665), .Y(n6448) );
	o22ai_1 U7044( .A1(n6210), .A2(n6067), .B1(n6277), .B2(n6450), .Y(n5794) );
	mux2i_1 U7045( .A0(n6451), .A1(n10213), .S(n10506), .Y(n6450) );
	o32ai_1 U7046( .A1(n6452), .A2(n10262), .A3(n6453), .B1(n6454), .B2(n6455), .Y(n5793) );
	o21ai_0 U7047( .A1(n10241), .A2(n6456), .B1(n6343), .Y(n6452) );
	o21ai_0 U7048( .A1(n6230), .A2(n6458), .B1(n6459), .Y(n5792) );
	mux2i_1 U7049( .A0(n6460), .A1(n6461), .S(n6462), .Y(n6459) );
	o21ai_0 U7050( .A1(n6230), .A2(n5987), .B1(n6463), .Y(n5791) );
	mux2i_1 U7051( .A0(n6464), .A1(n6249), .S(n6465), .Y(n6463) );
	nor2_1 U7052( .A(n6466), .B(n6467), .Y(n6465) );
	nor2_1 U7053( .A(n6308), .B(n6468), .Y(n6464) );
	nand2_1 U7054( .A(n6469), .B(n6470), .Y(n5790) );
	nand3_1 U7055( .A(n6471), .B(n6373), .C(n6472), .Y(n6470) );
	mux2i_1 U7056( .A0(n6473), .A1(n6474), .S(n10903), .Y(n6469) );
	nand2_1 U7057( .A(n6221), .B(n6475), .Y(n6474) );
	nand3_1 U7058( .A(n6380), .B(n6476), .C(n6477), .Y(n6475) );
	nor2_1 U7059( .A(n6478), .B(n6476), .Y(n6473) );
	o22ai_1 U7060( .A1(n6479), .A2(n6480), .B1(n6481), .B2(n6482), .Y(n5789) );
	a21oi_1 U7061( .A1(n6483), .A2(n6480), .B1(n6437), .Y(n6481) );
	o221ai_1 U7062( .A1(n6484), .A2(n6485), .B1(n6486), .B2(n6225), .C1(n6487), .Y(n5788) );
	nand3_1 U7063( .A(n10456), .B(g35), .C(n61), .Y(n6487) );
	o21ai_0 U7064( .A1(n6230), .A2(n5972), .B1(n6488), .Y(n5787) );
	mux2i_1 U7065( .A0(n6489), .A1(n6250), .S(n6490), .Y(n6488) );
	nor2_1 U7066( .A(n6491), .B(n6492), .Y(n6490) );
	nor2_1 U7067( .A(n6309), .B(n6493), .Y(n6489) );
	a21oi_1 U7068( .A1(n6198), .A2(n6494), .B1(n5915), .Y(n5786) );
	or2_0 U7069( .A(n6495), .B(n6369), .X(n6494) );
	o22ai_1 U7070( .A1(n6296), .A2(n6496), .B1(n6195), .B2(n5906), .Y(n5785) );
	o21ai_0 U7071( .A1(n6230), .A2(n6497), .B1(n6498), .Y(n5784) );
	mux2i_1 U7072( .A0(n6499), .A1(n6249), .S(n6500), .Y(n6498) );
	nor2_1 U7073( .A(n6501), .B(n6502), .Y(n6500) );
	nor2_1 U7074( .A(n6311), .B(n6503), .Y(n6499) );
	o32ai_1 U7075( .A1(n6310), .A2(n10417), .A3(n6504), .B1(n6201), .B2(n6505), .Y(n5783) );
	o21ai_0 U7076( .A1(n6368), .A2(n6506), .B1(n6248), .Y(n5782) );
	mux2i_1 U7077( .A0(n11779), .A1(g113), .S(n6507), .Y(n6506) );
	nor2_1 U7078( .A(n10660), .B(n6508), .Y(n6507) );
	o32ai_1 U7079( .A1(n6054), .A2(n6350), .A3(n6509), .B1(n6510), .B2(n6511), .Y(n5781) );
	mux2i_1 U7080( .A0(n6512), .A1(n6513), .S(n11845), .Y(n5780) );
	a21oi_1 U7081( .A1(n6378), .A2(n6514), .B1(n6437), .Y(n6513) );
	nand2_1 U7082( .A(n91), .B(g35), .Y(n6512) );
	nor2_1 U7083( .A(n6514), .B(n6363), .Y(n91) );
	inv_1 U7084( .A(g10306), .Y(n6514) );
	and2_0 U7085( .A(n6387), .B(g9555), .X(n5779) );
	o21ai_0 U7086( .A1(n6230), .A2(n5877), .B1(n6515), .Y(n5778) );
	mux2_1 U7087( .A0(n6516), .A1(n6517), .S(n10691), .X(n6515) );
	o21ai_0 U7088( .A1(n6230), .A2(n6037), .B1(n6518), .Y(n5777) );
	mux2i_1 U7089( .A0(n6519), .A1(n6520), .S(n6521), .Y(n6518) );
	nor2_1 U7090( .A(n6455), .B(n6522), .Y(n6521) );
	nor2_1 U7091( .A(n6310), .B(n6023), .Y(n6519) );
	o32ai_1 U7092( .A1(n6523), .A2(n6524), .A3(n6313), .B1(n6525), .B2(n6526), .Y(n5776) );
	a21oi_1 U7093( .A1(n6527), .A2(n10669), .B1(n6437), .Y(n6525) );
	nor2_1 U7094( .A(n6359), .B(n6524), .Y(n6527) );
	o22ai_1 U7095( .A1(n6211), .A2(n6070), .B1(n6528), .B2(n6295), .Y(n5775) );
	nor2_1 U7096( .A(n10233), .B(n10655), .Y(n6528) );
	o221ai_1 U7097( .A1(n6529), .A2(n6530), .B1(n6214), .B2(n6531), .C1(n6532), .Y(n5774) );
	o21ai_0 U7098( .A1(n6533), .A2(n6534), .B1(n10267), .Y(n6532) );
	nor3_1 U7099( .A(n6535), .B(n10520), .C(n6307), .Y(n6533) );
	nor2_1 U7100( .A(n6359), .B(n6536), .Y(n5773) );
	o22ai_1 U7101( .A1(n11781), .A2(n6302), .B1(n6194), .B2(n6537), .Y(n5772) );
	o21ai_0 U7102( .A1(n6231), .A2(n6538), .B1(n6539), .Y(n5771) );
	mux2i_1 U7103( .A0(n6540), .A1(n6249), .S(n6541), .Y(n6539) );
	nor2_1 U7104( .A(n6466), .B(n6542), .Y(n6541) );
	nor2_1 U7105( .A(n6313), .B(n6543), .Y(n6540) );
	o22ai_1 U7106( .A1(n6211), .A2(n6064), .B1(n6544), .B2(n6296), .Y(n5770) );
	o32ai_1 U7107( .A1(n6055), .A2(n6350), .A3(n6545), .B1(n6546), .B2(n6547), .Y(n5769) );
	o32ai_1 U7108( .A1(n6298), .A2(n6548), .A3(n6549), .B1(n6202), .B2(n6550), .Y(n5768) );
	a21oi_1 U7109( .A1(n6551), .A2(n6552), .B1(n10913), .Y(n6549) );
	nor3_1 U7110( .A(n6553), .B(n6404), .C(n6554), .Y(n6548) );
	xnor2_1 U7111( .A(n10282), .B(n6555), .Y(n6553) );
	nor2_1 U7112( .A(n6197), .B(n6556), .Y(n5767) );
	o21ai_0 U7113( .A1(n6232), .A2(n5989), .B1(n6557), .Y(n5766) );
	mux2i_1 U7114( .A0(n6558), .A1(n6559), .S(n6560), .Y(n6557) );
	and2_0 U7115( .A(n6561), .B(n6562), .X(n6560) );
	nor2_1 U7116( .A(n6312), .B(n6024), .Y(n6558) );
	nor2_1 U7117( .A(n6563), .B(n6564), .Y(n5765) );
	xnor2_1 U7118( .A(n6565), .B(n10361), .Y(n6563) );
	o21ai_0 U7119( .A1(n6232), .A2(n6566), .B1(n6567), .Y(n5764) );
	mux2i_1 U7120( .A0(n6568), .A1(n6250), .S(n6569), .Y(n6567) );
	nor2_1 U7121( .A(n6542), .B(n6570), .Y(n6569) );
	nor2_1 U7122( .A(n6295), .B(n6571), .Y(n6568) );
	o221ai_1 U7123( .A1(n6572), .A2(n6308), .B1(n6215), .B2(n6573), .C1(n6574), .Y(n5763) );
	nand4_1 U7124( .A(n10481), .B(n6575), .C(n6576), .D(n6577), .Y(n6574) );
	nor2_1 U7125( .A(n6359), .B(n6578), .Y(n6576) );
	a21oi_1 U7126( .A1(n10241), .A2(g35), .B1(n10262), .Y(n6578) );
	a21oi_1 U7127( .A1(n10481), .A2(n6579), .B1(n6580), .Y(n6572) );
	a21oi_1 U7128( .A1(n6577), .A2(n6575), .B1(n6581), .Y(n6580) );
	a21oi_1 U7129( .A1(n6582), .A2(n6583), .B1(n6584), .Y(n6581) );
	nand2_1 U7130( .A(n6585), .B(n6586), .Y(n6575) );
	o221ai_1 U7131( .A1(n6587), .A2(n6588), .B1(n6215), .B2(n5966), .C1(n6589), .Y(n5762) );
	a21oi_1 U7132( .A1(n10176), .A2(n6590), .B1(n6591), .Y(n6589) );
	o21ai_0 U7133( .A1(n6232), .A2(n6592), .B1(n6593), .Y(n5761) );
	mux2i_1 U7134( .A0(n6594), .A1(n6595), .S(n6596), .Y(n6593) );
	and2_0 U7135( .A(n6597), .B(n6598), .X(n6595) );
	nor2_1 U7136( .A(n6597), .B(n6599), .Y(n6594) );
	o21ai_0 U7137( .A1(n6233), .A2(n6476), .B1(n6600), .Y(n5760) );
	a22oi_1 U7138( .A1(n6601), .A2(n6602), .B1(n6603), .B2(n10903), .Y(n6600) );
	xnor2_1 U7139( .A(n6604), .B(n6605), .Y(n6601) );
	nand2_1 U7140( .A(n10903), .B(n6606), .Y(n6604) );
	nand3_1 U7141( .A(g16624), .B(n6607), .C(n10379), .Y(n6606) );
	mux2i_1 U7142( .A0(n6608), .A1(n6609), .S(n10717), .Y(n5759) );
	a21oi_1 U7143( .A1(n6378), .A2(n6610), .B1(n6437), .Y(n6609) );
	nand2_1 U7144( .A(n10214), .B(n6335), .Y(n6608) );
	o21ai_0 U7145( .A1(n6233), .A2(n5947), .B1(n6611), .Y(n5758) );
	mux2i_1 U7146( .A0(n6612), .A1(n6613), .S(n10685), .Y(n6611) );
	nor2_1 U7147( .A(n6288), .B(n6614), .Y(n6612) );
	inv_1 U7148( .A(n6615), .Y(n5757) );
	a221oi_1 U7149( .A1(n6616), .A2(n10636), .B1(n6437), .B2(n10323), .C1(n6617), .Y(n6615) );
	inv_1 U7150( .A(n6618), .Y(n6617) );
	o21ai_0 U7151( .A1(n6232), .A2(n5869), .B1(n6619), .Y(n5756) );
	mux2i_1 U7152( .A0(n6620), .A1(n6621), .S(n6622), .Y(n6619) );
	inv_1 U7153( .A(n6623), .Y(n6621) );
	o21ai_0 U7154( .A1(n6232), .A2(n5927), .B1(n6624), .Y(n5755) );
	mux2i_1 U7155( .A0(n6625), .A1(n6249), .S(n6626), .Y(n6624) );
	nor2_1 U7156( .A(n6627), .B(n6628), .Y(n6626) );
	nor2_1 U7157( .A(n6289), .B(n6629), .Y(n6625) );
	o22ai_1 U7158( .A1(n5954), .A2(n6630), .B1(n6631), .B2(n6632), .Y(n5754) );
	o211ai_1 U7159( .A1(n6203), .A2(n6633), .B1(n6400), .C1(n6634), .Y(n5753) );
	mux2i_1 U7160( .A0(n6635), .A1(n6636), .S(n6637), .Y(n6634) );
	nor2_1 U7161( .A(n6359), .B(n6638), .Y(n6636) );
	and2_0 U7162( .A(n6638), .B(n6345), .X(n6635) );
	o21ai_0 U7163( .A1(n6232), .A2(n6639), .B1(n6640), .Y(n5752) );
	a22oi_1 U7164( .A1(n10797), .A2(n6613), .B1(g26801), .B2(n6249), .Y(n6640) );
	inv_1 U7165( .A(n6510), .Y(n6613) );
	o21ai_0 U7166( .A1(n6232), .A2(n6641), .B1(n6642), .Y(n5751) );
	mux2i_1 U7167( .A0(n6643), .A1(n6644), .S(n6645), .Y(n6642) );
	nor2_1 U7168( .A(n6646), .B(n6647), .Y(n6644) );
	and2_0 U7169( .A(n6647), .B(n6648), .X(n6643) );
	o21ai_0 U7170( .A1(n6232), .A2(n5878), .B1(n6649), .Y(n5750) );
	mux2i_1 U7171( .A0(n6650), .A1(n6651), .S(n6652), .Y(n6649) );
	nor2_1 U7172( .A(n6293), .B(n6653), .Y(n6651) );
	o221ai_1 U7173( .A1(n6654), .A2(n6655), .B1(n6215), .B2(n6656), .C1(n6657), .Y(n5749) );
	inv_1 U7174( .A(n10686), .Y(n6656) );
	inv_1 U7175( .A(n10646), .Y(n6655) );
	o22ai_1 U7176( .A1(n6303), .A2(n6658), .B1(n6194), .B2(n6659), .Y(n5748) );
	o21ai_0 U7177( .A1(n6232), .A2(n6660), .B1(n6661), .Y(n5747) );
	a22oi_1 U7178( .A1(n10823), .A2(n6662), .B1(n6663), .B2(n6249), .Y(n6661) );
	o21ai_0 U7179( .A1(n6231), .A2(n6664), .B1(n6665), .Y(n5746) );
	mux2i_1 U7180( .A0(n6666), .A1(n6250), .S(n6667), .Y(n6665) );
	nor2_1 U7181( .A(n6668), .B(n6669), .Y(n6667) );
	nor2_1 U7182( .A(n6292), .B(n5925), .Y(n6666) );
	o21ai_0 U7183( .A1(n6231), .A2(n6670), .B1(n6671), .Y(n5745) );
	mux2i_1 U7184( .A0(n6672), .A1(n6250), .S(n6673), .Y(n6671) );
	nor2_1 U7185( .A(n6502), .B(n6674), .Y(n6673) );
	nor2_1 U7186( .A(n6285), .B(n6675), .Y(n6672) );
	o21ai_0 U7187( .A1(n6231), .A2(n6676), .B1(n6677), .Y(n5744) );
	mux2i_1 U7188( .A0(n6678), .A1(n6250), .S(n6679), .Y(n6677) );
	nor2_1 U7189( .A(n6680), .B(n6681), .Y(n6679) );
	nor2_1 U7190( .A(n6279), .B(n6682), .Y(n6678) );
	o221ai_1 U7191( .A1(n6683), .A2(n19450), .B1(n6684), .B2(n6685), .C1(n6686), .Y(n5743) );
	o21ai_0 U7192( .A1(n6231), .A2(n6687), .B1(n6688), .Y(n5742) );
	a22oi_1 U7193( .A1(n10745), .A2(n6689), .B1(n6690), .B2(n6249), .Y(n6688) );
	o21ai_0 U7194( .A1(n6231), .A2(n6691), .B1(n6692), .Y(n5741) );
	mux2i_1 U7195( .A0(n6603), .A1(n6693), .S(n6694), .Y(n6692) );
	nor2_1 U7196( .A(n6695), .B(n6696), .Y(n6693) );
	inv_1 U7197( .A(n6602), .Y(n6696) );
	o21ai_0 U7198( .A1(n6231), .A2(n6697), .B1(n6698), .Y(n5740) );
	a22oi_1 U7199( .A1(n6699), .A2(n6700), .B1(n6701), .B2(n10900), .Y(n6698) );
	xnor2_1 U7200( .A(n6702), .B(n6703), .Y(n6699) );
	nand2_1 U7201( .A(n10900), .B(n6704), .Y(n6702) );
	o221ai_1 U7202( .A1(n6705), .A2(n5891), .B1(n6706), .B2(n6707), .C1(n6708), .Y(n5739) );
	a21oi_1 U7203( .A1(n6709), .A2(n6381), .B1(n6437), .Y(n6705) );
	o32ai_1 U7204( .A1(n6710), .A2(n6278), .A3(n6711), .B1(n6712), .B2(n6713), .Y(n5738) );
	a21oi_1 U7205( .A1(n6714), .A2(n6381), .B1(n6437), .Y(n6712) );
	o21ai_0 U7206( .A1(n6033), .A2(n6715), .B1(n6716), .Y(n6710) );
	o21ai_0 U7207( .A1(n6231), .A2(n6038), .B1(n6717), .Y(n5737) );
	mux2i_1 U7208( .A0(n6718), .A1(n6719), .S(n10686), .Y(n6717) );
	nor2_1 U7209( .A(n6285), .B(n6720), .Y(n6718) );
	o21ai_0 U7210( .A1(n6230), .A2(n6721), .B1(n6722), .Y(n5736) );
	mux2i_1 U7211( .A0(n6723), .A1(n6724), .S(n6725), .Y(n6722) );
	nor2_1 U7212( .A(n6726), .B(n6727), .Y(n6724) );
	and2_0 U7213( .A(n6346), .B(n6726), .X(n6723) );
	nor2_1 U7214( .A(n10183), .B(n10151), .Y(n6726) );
	o22ai_1 U7215( .A1(n6303), .A2(n6728), .B1(n6194), .B2(n6729), .Y(n5735) );
	inv_1 U7216( .A(n10453), .Y(n6729) );
	o21ai_0 U7217( .A1(n6230), .A2(n6088), .B1(n6730), .Y(n5734) );
	mux2i_1 U7218( .A0(n6731), .A1(n6732), .S(n6733), .Y(n6730) );
	nor2_1 U7219( .A(n10564), .B(n6363), .Y(n6732) );
	nor2_1 U7220( .A(n6734), .B(n6735), .Y(n6731) );
	o221ai_1 U7221( .A1(n6736), .A2(n5918), .B1(n10333), .B2(n6737), .C1(n6738), .Y(n5733) );
	mux2i_1 U7222( .A0(n6739), .A1(n6740), .S(n6741), .Y(n6738) );
	nor4_1 U7223( .A(n6742), .B(n6743), .C(n6744), .D(n6745), .Y(n6740) );
	nand2_1 U7224( .A(n6224), .B(n6737), .Y(n6739) );
	a211oi_1 U7225( .A1(n6329), .A2(n6743), .B1(n6746), .C1(n6747), .Y(n6736) );
	o22ai_1 U7226( .A1(n6303), .A2(n6748), .B1(n6194), .B2(n6749), .Y(n5732) );
	o32ai_1 U7227( .A1(n6056), .A2(n6350), .A3(n6750), .B1(n6751), .B2(n6752), .Y(n5731) );
	o221ai_1 U7228( .A1(n5896), .A2(n6753), .B1(n6213), .B2(n6754), .C1(n6755), .Y(n5730) );
	a21oi_1 U7229( .A1(n6756), .A2(n6757), .B1(n6758), .Y(n6755) );
	nor2_1 U7230( .A(n10332), .B(n6759), .Y(n6756) );
	nand3_1 U7231( .A(n6760), .B(n6761), .C(n6762), .Y(n5729) );
	nand2_1 U7232( .A(g4546), .B(n6763), .Y(n6762) );
	o21ai_0 U7233( .A1(n6764), .A2(n6765), .B1(n6766), .Y(n5728) );
	mux2i_1 U7234( .A0(n6767), .A1(n6768), .S(n10546), .Y(n6766) );
	nand2_1 U7235( .A(n6223), .B(n6769), .Y(n6768) );
	nand3_1 U7236( .A(n6770), .B(n6373), .C(n6771), .Y(n6769) );
	nor2_1 U7237( .A(n6286), .B(n6770), .Y(n6767) );
	nand2_1 U7238( .A(n10677), .B(n6772), .Y(n6770) );
	o211ai_1 U7239( .A1(n6203), .A2(n6773), .B1(n6774), .C1(n6775), .Y(n5727) );
	mux2i_1 U7240( .A0(n6776), .A1(n6777), .S(n6420), .Y(n6775) );
	nor2_1 U7241( .A(n6359), .B(n6421), .Y(n6777) );
	nor3_1 U7242( .A(n6727), .B(n6778), .C(n6779), .Y(n6776) );
	mux2i_1 U7243( .A0(n6780), .A1(n6781), .S(n10197), .Y(n5726) );
	a21oi_1 U7244( .A1(n6782), .A2(n6783), .B1(n6437), .Y(n6781) );
	or2_0 U7245( .A(n6784), .B(n6783), .X(n6780) );
	o21ai_0 U7246( .A1(n6229), .A2(n6785), .B1(n6786), .Y(n5725) );
	mux2i_1 U7247( .A0(n6787), .A1(n6250), .S(n6788), .Y(n6786) );
	nor2_1 U7248( .A(n6491), .B(n6789), .Y(n6788) );
	nor2_1 U7249( .A(n6296), .B(n6790), .Y(n6787) );
	mux2i_1 U7250( .A0(n6791), .A1(n6792), .S(n6793), .Y(n5724) );
	nand2_1 U7251( .A(n6794), .B(n10362), .Y(n6792) );
	a21oi_1 U7252( .A1(n6648), .A2(n6641), .B1(n6437), .Y(n6791) );
	o21ai_0 U7253( .A1(n6229), .A2(n6795), .B1(n6796), .Y(n5723) );
	mux2i_1 U7254( .A0(n6797), .A1(n6798), .S(n6799), .Y(n6796) );
	and2_0 U7255( .A(n6387), .B(n6800), .X(n6798) );
	nor2_1 U7256( .A(n6800), .B(n6298), .Y(n6797) );
	nor4_1 U7257( .A(n6801), .B(n6802), .C(n6795), .D(n10440), .Y(n6800) );
	o22ai_1 U7258( .A1(n6304), .A2(n6803), .B1(n6193), .B2(n6804), .Y(n5722) );
	o21ai_0 U7259( .A1(n6229), .A2(n5977), .B1(n6805), .Y(n5721) );
	mux2i_1 U7260( .A0(n6806), .A1(n6250), .S(n6807), .Y(n6805) );
	nor2_1 U7261( .A(n6680), .B(n6808), .Y(n6807) );
	nor2_1 U7262( .A(n6313), .B(n6809), .Y(n6806) );
	o21ai_0 U7263( .A1(n6810), .A2(n6811), .B1(n6812), .Y(n5720) );
	mux2i_1 U7264( .A0(n6813), .A1(n6814), .S(n6815), .Y(n6812) );
	nor2_1 U7265( .A(n6816), .B(n6817), .Y(n6814) );
	nand2_1 U7266( .A(n6223), .B(n6818), .Y(n6813) );
	nand3_1 U7267( .A(n6819), .B(n6373), .C(n6816), .Y(n6818) );
	o22ai_1 U7268( .A1(n6209), .A2(n6820), .B1(n6821), .B2(n6297), .Y(n5719) );
	nor2_1 U7269( .A(n10939), .B(n6822), .Y(n6821) );
	o22ai_1 U7270( .A1(n6209), .A2(n6823), .B1(n6299), .B2(n6824), .Y(n5718) );
	mux2i_1 U7271( .A0(n6825), .A1(n6826), .S(n6827), .Y(n6824) );
	nor2_1 U7272( .A(n10404), .B(n6825), .Y(n6826) );
	inv_1 U7273( .A(n6828), .Y(n6825) );
	o21ai_0 U7274( .A1(n6229), .A2(n6829), .B1(n6830), .Y(n5717) );
	mux2i_1 U7275( .A0(n6831), .A1(n6832), .S(n6833), .Y(n6830) );
	and2_0 U7276( .A(n6834), .B(n6835), .X(n6832) );
	o211ai_1 U7277( .A1(n6836), .A2(n6837), .B1(n6838), .C1(n6839), .Y(n5716) );
	nand3_1 U7278( .A(n11941), .B(n6840), .C(n6841), .Y(n6838) );
	a21oi_1 U7279( .A1(n6842), .A2(n6843), .B1(n6437), .Y(n6836) );
	o221ai_1 U7280( .A1(n6037), .A2(n6844), .B1(n6845), .B2(n6846), .C1(n6847), .Y(n5715) );
	a22oi_1 U7281( .A1(n10554), .A2(n6848), .B1(n10335), .B2(n6437), .Y(n6847) );
	inv_1 U7282( .A(n6849), .Y(n6846) );
	a221oi_1 U7283( .A1(n10723), .A2(n6850), .B1(n6851), .B2(n11780), .C1(n6852), .Y(n6845) );
	o32ai_1 U7284( .A1(n6853), .A2(n11950), .A3(n10335), .B1(n10174), .B2(n6854), .Y(n6852) );
	a22oi_1 U7285( .A1(n11809), .A2(n10335), .B1(n11822), .B2(n11950), .Y(n6854) );
	o21ai_0 U7286( .A1(n6229), .A2(n5974), .B1(n6855), .Y(n5714) );
	mux2i_1 U7287( .A0(n6856), .A1(n6250), .S(n6857), .Y(n6855) );
	nor2_1 U7288( .A(n6628), .B(n6858), .Y(n6857) );
	nor2_1 U7289( .A(n6278), .B(n6859), .Y(n6856) );
	o21ai_0 U7290( .A1(n6228), .A2(n6043), .B1(n6860), .Y(n5713) );
	mux2i_1 U7291( .A0(n6861), .A1(n6862), .S(n6863), .Y(n6860) );
	nor2_1 U7292( .A(n6290), .B(n6864), .Y(n6862) );
	o21ai_0 U7293( .A1(n6228), .A2(n6865), .B1(n6866), .Y(n5712) );
	inv_1 U7294( .A(n6867), .Y(n6866) );
	o22ai_1 U7295( .A1(n6868), .A2(n6869), .B1(n6870), .B2(n6871), .Y(n6867) );
	nor2_1 U7296( .A(n6359), .B(n6872), .Y(n5711) );
	o21ai_0 U7297( .A1(n6654), .A2(n6873), .B1(n6874), .Y(n5710) );
	mux2i_1 U7298( .A0(n6875), .A1(n6876), .S(n10646), .Y(n6874) );
	nand2_1 U7299( .A(n6224), .B(n6657), .Y(n6876) );
	nand3_1 U7300( .A(n6477), .B(n6374), .C(n10686), .Y(n6657) );
	nor2_1 U7301( .A(n10686), .B(n6478), .Y(n6875) );
	nor2_1 U7302( .A(n6877), .B(n6301), .Y(n5709) );
	nor4_1 U7303( .A(n6878), .B(n6879), .C(n6880), .D(n6881), .Y(n6877) );
	nand3_1 U7304( .A(n10245), .B(n6882), .C(n10160), .Y(n6878) );
	o32ai_1 U7305( .A1(n6310), .A2(g8342), .A3(n6883), .B1(n6199), .B2(n6884), .Y(n5708) );
	a21oi_1 U7306( .A1(g8279), .A2(n6884), .B1(n10618), .Y(n6883) );
	inv_1 U7307( .A(n10617), .Y(n6884) );
	o21ai_0 U7308( .A1(n6227), .A2(n5994), .B1(n6885), .Y(n5707) );
	mux2i_1 U7309( .A0(n6886), .A1(n6250), .S(n6887), .Y(n6885) );
	nor2_1 U7310( .A(n6888), .B(n6669), .Y(n6887) );
	nor2_1 U7311( .A(n6290), .B(n6015), .Y(n6886) );
	o221ai_1 U7312( .A1(n6683), .A2(n19451), .B1(n6684), .B2(n6685), .C1(n6889), .Y(n5706) );
	inv_1 U7313( .A(n6763), .Y(n6683) );
	o221ai_1 U7314( .A1(n6890), .A2(n6891), .B1(n6218), .B2(n5963), .C1(n6892), .Y(n5705) );
	a21oi_1 U7315( .A1(n6849), .A2(n10174), .B1(n6893), .Y(n6892) );
	o21ai_0 U7316( .A1(n6227), .A2(n6894), .B1(n6895), .Y(n5704) );
	mux2i_1 U7317( .A0(n6896), .A1(n6250), .S(n6897), .Y(n6895) );
	nor2_1 U7318( .A(n6898), .B(n6899), .Y(n6897) );
	nor2_1 U7319( .A(n6290), .B(n6900), .Y(n6896) );
	o21ai_0 U7320( .A1(n6227), .A2(n6901), .B1(n6902), .Y(n5703) );
	mux2i_1 U7321( .A0(n6903), .A1(n6250), .S(n6904), .Y(n6902) );
	nor2_1 U7322( .A(n6905), .B(n6906), .Y(n6904) );
	nor2_1 U7323( .A(n6291), .B(n6907), .Y(n6903) );
	o32ai_1 U7324( .A1(n6310), .A2(n6908), .A3(n6909), .B1(n6199), .B2(n6910), .Y(n5702) );
	a21oi_1 U7325( .A1(n6911), .A2(n6551), .B1(n10910), .Y(n6909) );
	nor3_1 U7326( .A(n6912), .B(n6554), .C(n6407), .Y(n6908) );
	xnor2_1 U7327( .A(n10284), .B(n6555), .Y(n6912) );
	o22ai_1 U7328( .A1(n6303), .A2(n5897), .B1(n6193), .B2(n6748), .Y(n5701) );
	o221ai_1 U7329( .A1(n6913), .A2(n6914), .B1(n6218), .B2(n5885), .C1(n6915), .Y(n5700) );
	nand3_1 U7330( .A(n10525), .B(n6374), .C(n6916), .Y(n6915) );
	o21ai_0 U7331( .A1(n6917), .A2(n6918), .B1(n6919), .Y(n6914) );
	inv_1 U7332( .A(n6920), .Y(n57) );
	a21oi_1 U7333( .A1(n6437), .A2(n10656), .B1(n5433), .Y(n6920) );
	a21oi_1 U7334( .A1(n6197), .A2(n6921), .B1(n5911), .Y(n5699) );
	or2_0 U7335( .A(n6504), .B(n6369), .X(n6921) );
	nor2_1 U7336( .A(n6505), .B(n6922), .Y(n6504) );
	o21ai_0 U7337( .A1(n6510), .A2(n6041), .B1(n6923), .Y(n5698) );
	mux2i_1 U7338( .A0(n6924), .A1(n6925), .S(n6511), .Y(n6923) );
	inv_1 U7339( .A(n10651), .Y(n6511) );
	nor3_1 U7340( .A(n6614), .B(n11909), .C(n6306), .Y(n6925) );
	inv_1 U7341( .A(g26801), .Y(n6614) );
	nand2_1 U7342( .A(n6224), .B(n6926), .Y(n6924) );
	nand3_1 U7343( .A(n11909), .B(n6374), .C(g26801), .Y(n6926) );
	o22ai_1 U7344( .A1(n6211), .A2(n6927), .B1(n6928), .B2(n6929), .Y(n5697) );
	o21ai_0 U7345( .A1(n6930), .A2(n6931), .B1(n6382), .Y(n6929) );
	a21oi_1 U7346( .A1(n6932), .A2(n6933), .B1(n6934), .Y(n6931) );
	mux2i_1 U7347( .A0(n6935), .A1(n10194), .S(n6936), .Y(n6928) );
	o22ai_1 U7348( .A1(n6304), .A2(n6937), .B1(n6193), .B2(n5897), .Y(n5696) );
	o21ai_0 U7349( .A1(n6706), .A2(n6938), .B1(n6939), .Y(n5695) );
	mux2i_1 U7350( .A0(n6940), .A1(n6941), .S(n10548), .Y(n6939) );
	nand2_1 U7351( .A(n6223), .B(n6942), .Y(n6941) );
	nand3_1 U7352( .A(n6943), .B(n6374), .C(n6709), .Y(n6942) );
	nor2_1 U7353( .A(n6278), .B(n6943), .Y(n6940) );
	nand2_1 U7354( .A(n10681), .B(n6944), .Y(n6943) );
	o21ai_0 U7355( .A1(n6226), .A2(n5937), .B1(n6945), .Y(n5694) );
	mux2i_1 U7356( .A0(n6946), .A1(n6250), .S(n6947), .Y(n6945) );
	nor2_1 U7357( .A(n6467), .B(n6502), .Y(n6947) );
	nor2_1 U7358( .A(n6293), .B(n6670), .Y(n6946) );
	inv_1 U7359( .A(n10835), .Y(n6670) );
	o21ai_0 U7360( .A1(n6226), .A2(n6948), .B1(n6949), .Y(n5693) );
	mux2_1 U7361( .A0(n6950), .A1(n6951), .S(n11878), .X(n6949) );
	o21ai_0 U7362( .A1(n6952), .A2(n6052), .B1(n6953), .Y(n5692) );
	mux2i_1 U7363( .A0(n6954), .A1(n6955), .S(n6956), .Y(n6953) );
	nor3_1 U7364( .A(n6957), .B(n10697), .C(n6306), .Y(n6955) );
	nand2_1 U7365( .A(n6224), .B(n6958), .Y(n6954) );
	nand3_1 U7366( .A(n6959), .B(n6374), .C(n10697), .Y(n6958) );
	o221ai_1 U7367( .A1(n6960), .A2(n6961), .B1(n6219), .B2(n6962), .C1(n6963), .Y(n5691) );
	inv_1 U7368( .A(n10320), .Y(n6962) );
	inv_1 U7369( .A(n10633), .Y(n6961) );
	o221ai_1 U7370( .A1(n6964), .A2(n6965), .B1(n6220), .B2(n6966), .C1(n6967), .Y(n5690) );
	nand3_1 U7371( .A(n6968), .B(n5932), .C(n6969), .Y(n6967) );
	o21ai_0 U7372( .A1(n6970), .A2(n6968), .B1(n6344), .Y(n6965) );
	xnor2_1 U7373( .A(n6555), .B(n10306), .Y(n6968) );
	o32ai_1 U7374( .A1(n6971), .A2(n10153), .A3(n6972), .B1(n6198), .B2(n5898), .Y(n5689) );
	o21ai_0 U7375( .A1(n6225), .A2(n5883), .B1(n6973), .Y(n5688) );
	o22ai_1 U7376( .A1(n6304), .A2(n6804), .B1(n6193), .B2(n6974), .Y(n5687) );
	o221ai_1 U7377( .A1(n6975), .A2(n6976), .B1(n6220), .B2(n6977), .C1(n6978), .Y(n5686) );
	nand2_1 U7378( .A(n6338), .B(n6979), .Y(n6976) );
	o32ai_1 U7379( .A1(n6980), .A2(n6350), .A3(n6981), .B1(n6982), .B2(n6983), .Y(n5685) );
	inv_1 U7380( .A(n10691), .Y(n6980) );
	inv_1 U7381( .A(n6984), .Y(n5684) );
	a221oi_1 U7382( .A1(n6620), .A2(n10631), .B1(n6437), .B2(n10318), .C1(n6985), .Y(n6984) );
	inv_1 U7383( .A(n6986), .Y(n6985) );
	o32ai_1 U7384( .A1(n6987), .A2(n6350), .A3(n6988), .B1(n6952), .B2(n6989), .Y(n5683) );
	inv_1 U7385( .A(n10484), .Y(n6987) );
	o21ai_0 U7386( .A1(n6227), .A2(n6990), .B1(n6991), .Y(n5682) );
	mux2i_1 U7387( .A0(n6992), .A1(n6251), .S(n6993), .Y(n6991) );
	nor2_1 U7388( .A(n6994), .B(n6995), .Y(n6993) );
	nor2_1 U7389( .A(n6292), .B(n6996), .Y(n6992) );
	o21ai_0 U7390( .A1(n6226), .A2(n6997), .B1(n6998), .Y(n5681) );
	mux2i_1 U7391( .A0(n6999), .A1(n6250), .S(n7000), .Y(n6998) );
	nor2_1 U7392( .A(n6570), .B(n6674), .Y(n7000) );
	nor2_1 U7393( .A(n6288), .B(n6538), .Y(n6999) );
	inv_1 U7394( .A(n10841), .Y(n6538) );
	o21ai_0 U7395( .A1(n6225), .A2(n6047), .B1(n7001), .Y(n5680) );
	mux2i_1 U7396( .A0(n7002), .A1(n7003), .S(n7004), .Y(n7001) );
	nor2_1 U7397( .A(n6287), .B(n7005), .Y(n7003) );
	o21ai_0 U7398( .A1(n6546), .A2(n6040), .B1(n7006), .Y(n5679) );
	mux2i_1 U7399( .A0(n7007), .A1(n7008), .S(n6547), .Y(n7006) );
	inv_1 U7400( .A(n10652), .Y(n6547) );
	nor3_1 U7401( .A(n6653), .B(n11911), .C(n6306), .Y(n7008) );
	nand2_1 U7402( .A(n6223), .B(n7009), .Y(n7007) );
	nand3_1 U7403( .A(n11911), .B(n6374), .C(n7010), .Y(n7009) );
	o21ai_0 U7404( .A1(n6226), .A2(n7011), .B1(n7012), .Y(n5678) );
	mux2i_1 U7405( .A0(n7013), .A1(n6251), .S(n7014), .Y(n7012) );
	nor2_1 U7406( .A(n7015), .B(n7016), .Y(n7014) );
	nor2_1 U7407( .A(n6279), .B(n7017), .Y(n7013) );
	o21ai_0 U7408( .A1(n6227), .A2(n7018), .B1(n7019), .Y(n5677) );
	a22oi_1 U7409( .A1(n11771), .A2(n7020), .B1(n7021), .B2(n7022), .Y(n7019) );
	o21ai_0 U7410( .A1(n6226), .A2(n5980), .B1(n7023), .Y(n5676) );
	mux2i_1 U7411( .A0(n7024), .A1(n6251), .S(n7025), .Y(n7023) );
	nor2_1 U7412( .A(n6905), .B(n7026), .Y(n7025) );
	nor2_1 U7413( .A(n6292), .B(n7027), .Y(n7024) );
	o221ai_1 U7414( .A1(n7028), .A2(n7029), .B1(n6219), .B2(n7030), .C1(n7031), .Y(n5675) );
	o21ai_0 U7415( .A1(n7032), .A2(n6746), .B1(n11863), .Y(n7031) );
	inv_1 U7416( .A(n7033), .Y(n7032) );
	o21ai_0 U7417( .A1(n7029), .A2(n7034), .B1(n6343), .Y(n7033) );
	a21oi_1 U7418( .A1(n7035), .A2(n7036), .B1(n7037), .Y(n7028) );
	nor4_1 U7419( .A(n10249), .B(n7034), .C(n7038), .D(n7039), .Y(n7037) );
	a21oi_1 U7420( .A1(n10259), .A2(n7040), .B1(n6308), .Y(n7035) );
	o22ai_1 U7421( .A1(n6208), .A2(n7041), .B1(n7042), .B2(n6297), .Y(n5674) );
	nor2_1 U7422( .A(n10587), .B(n7043), .Y(n7042) );
	o21ai_0 U7423( .A1(n6227), .A2(n7044), .B1(n7045), .Y(n5673) );
	mux2i_1 U7424( .A0(n7046), .A1(n7047), .S(n6927), .Y(n7045) );
	and2_0 U7425( .A(n6935), .B(n7048), .X(n7047) );
	nand2_1 U7426( .A(n7049), .B(n7050), .Y(n6935) );
	inv_1 U7427( .A(n10416), .Y(n7044) );
	o21ai_0 U7428( .A1(n6226), .A2(n7051), .B1(n7052), .Y(n5672) );
	mux2i_1 U7429( .A0(n7053), .A1(n7054), .S(n10916), .Y(n7052) );
	nor2_1 U7430( .A(n7055), .B(n7056), .Y(n7054) );
	and2_0 U7431( .A(n7055), .B(n7057), .X(n7053) );
	and2_0 U7432( .A(n7058), .B(n10427), .X(n7055) );
	o221ai_1 U7433( .A1(n7059), .A2(n6810), .B1(n6218), .B2(n7060), .C1(n7061), .Y(n5671) );
	o21ai_0 U7434( .A1(n6226), .A2(n6025), .B1(n7062), .Y(n5670) );
	mux2i_1 U7435( .A0(n7063), .A1(n7064), .S(n7065), .Y(n7062) );
	nor2_1 U7436( .A(n10260), .B(n7066), .Y(n7065) );
	nor2_1 U7437( .A(n6292), .B(n5984), .Y(n7063) );
	inv_1 U7438( .A(n7067), .Y(n5669) );
	o21ai_0 U7439( .A1(n11775), .A2(n11859), .B1(n6343), .Y(n7067) );
	o21ai_0 U7440( .A1(n6226), .A2(n5982), .B1(n7068), .Y(n5668) );
	mux2i_1 U7441( .A0(n7069), .A1(n6251), .S(n7070), .Y(n7068) );
	nor2_1 U7442( .A(n7071), .B(n7072), .Y(n7070) );
	nor2_1 U7443( .A(n6293), .B(n5971), .Y(n7069) );
	o21ai_0 U7444( .A1(n6227), .A2(n5942), .B1(n7073), .Y(n5667) );
	mux2_1 U7445( .A0(n7074), .A1(n7075), .S(n10696), .X(n7073) );
	nor2_1 U7446( .A(n6292), .B(n7076), .Y(n5666) );
	o21ai_0 U7447( .A1(n6226), .A2(n7077), .B1(n7078), .Y(n5665) );
	mux2i_1 U7448( .A0(n7079), .A1(n7080), .S(n7081), .Y(n7078) );
	nor2_1 U7449( .A(n6360), .B(n7082), .Y(n7080) );
	and2_0 U7450( .A(n7082), .B(n7083), .X(n7079) );
	o32ai_1 U7451( .A1(n6311), .A2(n7084), .A3(n7085), .B1(n6198), .B2(n7086), .Y(n5664) );
	a21oi_1 U7452( .A1(n7087), .A2(n7088), .B1(n10581), .Y(n7085) );
	nor4_1 U7453( .A(n10239), .B(n6742), .C(n7089), .D(n7090), .Y(n7084) );
	o22ai_1 U7454( .A1(n6208), .A2(n7091), .B1(n6277), .B2(n7092), .Y(n5663) );
	o22ai_1 U7455( .A1(n10412), .A2(n7093), .B1(n7094), .B2(n7095), .Y(n7092) );
	nor3_1 U7456( .A(n7096), .B(n7097), .C(n7098), .Y(n7093) );
	o221ai_1 U7457( .A1(n7099), .A2(n5893), .B1(n7100), .B2(n6891), .C1(n7101), .Y(n5662) );
	a21oi_1 U7458( .A1(n7102), .A2(n6370), .B1(n6437), .Y(n7099) );
	o21ai_0 U7459( .A1(n6226), .A2(n7103), .B1(n7104), .Y(n5661) );
	mux2i_1 U7460( .A0(n7105), .A1(n7106), .S(n7107), .Y(n7104) );
	nor2_1 U7461( .A(n10390), .B(n6363), .Y(n7106) );
	nor2_1 U7462( .A(n7108), .B(n7109), .Y(n7105) );
	o221ai_1 U7463( .A1(n7110), .A2(n7111), .B1(n6218), .B2(n7089), .C1(n7112), .Y(n5660) );
	or3_1 U7464( .A(n7113), .B(n6369), .C(n7066), .X(n7112) );
	o22ai_1 U7465( .A1(n6207), .A2(n7114), .B1(n7115), .B2(n6297), .Y(n5659) );
	xnor2_1 U7466( .A(n10669), .B(n10921), .Y(n7115) );
	o21ai_0 U7467( .A1(n6226), .A2(n6036), .B1(n7116), .Y(n5658) );
	mux2i_1 U7468( .A0(n7117), .A1(n7118), .S(n7119), .Y(n7116) );
	nor2_1 U7469( .A(n7120), .B(n7121), .Y(n7119) );
	nor2_1 U7470( .A(n6292), .B(n6021), .Y(n7117) );
	o22ai_1 U7471( .A1(n6207), .A2(n7122), .B1(n6277), .B2(n7123), .Y(n5657) );
	nor2_1 U7472( .A(n6360), .B(n7124), .Y(n5656) );
	and2_0 U7473( .A(n6387), .B(g9553), .X(n5655) );
	o21ai_0 U7474( .A1(n6228), .A2(n5934), .B1(n7125), .Y(n5654) );
	mux2i_1 U7475( .A0(n7126), .A1(n7127), .S(n7128), .Y(n7125) );
	nor2_1 U7476( .A(n7129), .B(n7130), .Y(n7127) );
	nor2_1 U7477( .A(n7131), .B(n6299), .Y(n7126) );
	o221ai_1 U7478( .A1(n6441), .A2(n6445), .B1(n6219), .B2(n7132), .C1(n6447), .Y(n5653) );
	nand3_1 U7479( .A(n7133), .B(n6374), .C(n10325), .Y(n6447) );
	inv_1 U7480( .A(n10638), .Y(n6445) );
	o21ai_0 U7481( .A1(n6227), .A2(n7134), .B1(n7135), .Y(n5652) );
	a22oi_1 U7482( .A1(n7136), .A2(n7137), .B1(n7138), .B2(n10847), .Y(n7135) );
	o22ai_1 U7483( .A1(n7139), .A2(n6302), .B1(n7140), .B2(n7141), .Y(n5651) );
	a21oi_1 U7484( .A1(n6378), .A2(n7142), .B1(n6437), .Y(n7140) );
	a21oi_1 U7485( .A1(n10473), .A2(n7141), .B1(n7143), .Y(n7139) );
	xnor2_1 U7486( .A(n7144), .B(n10519), .Y(n7143) );
	o21ai_0 U7487( .A1(n6227), .A2(n6571), .B1(n7145), .Y(n5650) );
	mux2i_1 U7488( .A0(n7146), .A1(n6251), .S(n7147), .Y(n7145) );
	nor2_1 U7489( .A(n6501), .B(n6570), .Y(n7147) );
	nor2_1 U7490( .A(n6293), .B(n7148), .Y(n7146) );
	inv_1 U7491( .A(n10840), .Y(n6571) );
	o21ai_0 U7492( .A1(n6228), .A2(n5941), .B1(n7149), .Y(n5649) );
	mux2i_1 U7493( .A0(n7150), .A1(n7151), .S(n7152), .Y(n7149) );
	nor2_1 U7494( .A(n6294), .B(n5931), .Y(n7151) );
	nor2_1 U7495( .A(n11947), .B(n6363), .Y(n7150) );
	o221ai_1 U7496( .A1(n7153), .A2(n5876), .B1(n6216), .B2(n7154), .C1(n7155), .Y(n5648) );
	nand3_1 U7497( .A(n7156), .B(n7157), .C(n7158), .Y(n7155) );
	xnor2_1 U7498( .A(n7159), .B(n10679), .Y(n7157) );
	a21oi_1 U7499( .A1(n6332), .A2(n7160), .B1(n7161), .Y(n7153) );
	o221ai_1 U7500( .A1(n7162), .A2(n7163), .B1(n6218), .B2(n7164), .C1(n7165), .Y(n5647) );
	inv_1 U7501( .A(n10684), .Y(n7164) );
	inv_1 U7502( .A(n10642), .Y(n7163) );
	o32ai_1 U7503( .A1(n6311), .A2(n10419), .A3(n7166), .B1(n6199), .B2(n7167), .Y(n5646) );
	o21ai_0 U7504( .A1(n7168), .A2(n6093), .B1(n7169), .Y(n5645) );
	mux2i_1 U7505( .A0(n7170), .A1(n7171), .S(n7172), .Y(n7169) );
	nor2_1 U7506( .A(n10322), .B(n6844), .Y(n7171) );
	nand2_1 U7507( .A(n6224), .B(n7173), .Y(n7170) );
	o21ai_0 U7508( .A1(n6227), .A2(n7174), .B1(n7175), .Y(n5644) );
	mux2i_1 U7509( .A0(n7176), .A1(n6251), .S(n7177), .Y(n7175) );
	nor2_1 U7510( .A(n6868), .B(n7178), .Y(n7177) );
	nor2_1 U7511( .A(n6293), .B(n5939), .Y(n7176) );
	o21ai_0 U7512( .A1(n6228), .A2(n7179), .B1(n7180), .Y(n5643) );
	mux2_1 U7513( .A0(n7181), .A1(n7182), .S(n11909), .X(n7180) );
	o21ai_0 U7514( .A1(n6228), .A2(n6019), .B1(n7183), .Y(n5642) );
	mux2i_1 U7515( .A0(n7184), .A1(n6251), .S(n7185), .Y(n7183) );
	nor2_1 U7516( .A(n6467), .B(n7186), .Y(n7185) );
	nor2_1 U7517( .A(n6294), .B(n7187), .Y(n7184) );
	and2_0 U7518( .A(g4520), .B(n6383), .X(n5641) );
	o21ai_0 U7519( .A1(n6228), .A2(n6675), .B1(n7188), .Y(n5640) );
	mux2i_1 U7520( .A0(n7189), .A1(n6251), .S(n7190), .Y(n7188) );
	nor2_1 U7521( .A(n6542), .B(n7186), .Y(n7190) );
	nor2_1 U7522( .A(n6293), .B(n7191), .Y(n7189) );
	a21oi_1 U7523( .A1(n7192), .A2(n7193), .B1(n6308), .Y(n5639) );
	o211ai_1 U7524( .A1(n7194), .A2(n7195), .B1(n7196), .C1(n7197), .Y(n7193) );
	mux2i_1 U7525( .A0(n7198), .A1(n7199), .S(n6691), .Y(n7195) );
	inv_1 U7526( .A(n10420), .Y(n6691) );
	mux2i_1 U7527( .A0(n7200), .A1(n7201), .S(n5909), .Y(n7194) );
	o21ai_0 U7528( .A1(n7197), .A2(n7202), .B1(n10596), .Y(n7192) );
	o21ai_0 U7529( .A1(n6228), .A2(n7203), .B1(n7204), .Y(n5638) );
	a22oi_1 U7530( .A1(n11787), .A2(n7046), .B1(n7048), .B2(n7205), .Y(n7204) );
	o32ai_1 U7531( .A1(n7206), .A2(n10592), .A3(n6313), .B1(n6200), .B2(n7207), .Y(n5637) );
	o21ai_0 U7532( .A1(n7208), .A2(n6044), .B1(n7209), .Y(n5636) );
	mux2i_1 U7533( .A0(n7210), .A1(n7211), .S(n10897), .Y(n7209) );
	nand2_1 U7534( .A(n6224), .B(n7212), .Y(n7211) );
	nand3_1 U7535( .A(n6379), .B(n7213), .C(n7214), .Y(n7212) );
	nor2_1 U7536( .A(n7215), .B(n7213), .Y(n7210) );
	o32ai_1 U7537( .A1(n6311), .A2(n7216), .A3(n7217), .B1(n6200), .B2(n7218), .Y(n5635) );
	a21oi_1 U7538( .A1(n7219), .A2(n7220), .B1(n10584), .Y(n7217) );
	nor4_1 U7539( .A(n10242), .B(n7221), .C(n7222), .D(n7223), .Y(n7216) );
	o21ai_0 U7540( .A1(n6228), .A2(n7224), .B1(n7225), .Y(n5634) );
	mux2i_1 U7541( .A0(n7226), .A1(n6251), .S(n7227), .Y(n7225) );
	nor2_1 U7542( .A(n7228), .B(n7229), .Y(n7227) );
	nor2_1 U7543( .A(n6294), .B(n7230), .Y(n7226) );
	o21ai_0 U7544( .A1(n6229), .A2(n7231), .B1(n7232), .Y(n5633) );
	mux2i_1 U7545( .A0(n7233), .A1(n7234), .S(n7235), .Y(n7232) );
	nor2_1 U7546( .A(n6360), .B(n7236), .Y(n7234) );
	and2_0 U7547( .A(n7236), .B(n7237), .X(n7233) );
	o22ai_1 U7548( .A1(n7238), .A2(n7239), .B1(n7240), .B2(n7241), .Y(n5632) );
	a21oi_1 U7549( .A1(n7242), .A2(n7238), .B1(n6437), .Y(n7240) );
	o21ai_0 U7550( .A1(n6751), .A2(n7243), .B1(n7244), .Y(n5631) );
	mux2i_1 U7551( .A0(n7245), .A1(n7246), .S(n6752), .Y(n7244) );
	inv_1 U7552( .A(n10649), .Y(n6752) );
	nor3_1 U7553( .A(n6864), .B(n11919), .C(n6307), .Y(n7246) );
	nand2_1 U7554( .A(n6224), .B(n7247), .Y(n7245) );
	nand3_1 U7555( .A(n11919), .B(n6375), .C(n7248), .Y(n7247) );
	inv_1 U7556( .A(n10661), .Y(n7243) );
	o21ai_0 U7557( .A1(n6229), .A2(n7249), .B1(n7250), .Y(n5630) );
	mux2i_1 U7558( .A0(n7251), .A1(n6251), .S(n7252), .Y(n7250) );
	nor2_1 U7559( .A(n6502), .B(n6542), .Y(n7252) );
	nand3_1 U7560( .A(n7253), .B(n7254), .C(n6674), .Y(n6542) );
	nor2_1 U7561( .A(n6293), .B(n6497), .Y(n7251) );
	nor3_1 U7562( .A(n7255), .B(n6351), .C(n7256), .Y(n5629) );
	a21oi_1 U7563( .A1(n10854), .A2(n6545), .B1(n7257), .Y(n7256) );
	nor3_1 U7564( .A(n7258), .B(n7259), .C(n7010), .Y(n7255) );
	o32ai_1 U7565( .A1(n7260), .A2(n6828), .A3(n6313), .B1(n7261), .B2(n6827), .Y(n5628) );
	inv_1 U7566( .A(n10445), .Y(n6827) );
	a21oi_1 U7567( .A1(n7262), .A2(n6828), .B1(n6437), .Y(n7261) );
	nor2_1 U7568( .A(n10404), .B(n6363), .Y(n7262) );
	o22ai_1 U7569( .A1(n6305), .A2(n7263), .B1(n6193), .B2(n7264), .Y(n5627) );
	o221ai_1 U7570( .A1(n6305), .A2(n7265), .B1(n6213), .B2(n7266), .C1(n7267), .Y(n5626) );
	mux2i_1 U7571( .A0(n7268), .A1(n7269), .S(n7270), .Y(n7267) );
	nor2_1 U7572( .A(n6360), .B(n7271), .Y(n7269) );
	nor3_1 U7573( .A(n6727), .B(n7272), .C(n7273), .Y(n7268) );
	and2_0 U7574( .A(n6386), .B(g8353), .X(n5625) );
	o32ai_1 U7575( .A1(n7274), .A2(n7275), .A3(n7276), .B1(n7277), .B2(n6197), .Y(n5624) );
	o21ai_0 U7576( .A1(n7278), .A2(n11788), .B1(n6343), .Y(n7274) );
	nor3_1 U7577( .A(n7279), .B(n7280), .C(n7281), .Y(n7278) );
	a21oi_1 U7578( .A1(n6198), .A2(n7282), .B1(n5910), .Y(n5623) );
	or2_0 U7579( .A(n7283), .B(n6369), .X(n7282) );
	o21ai_0 U7580( .A1(n6229), .A2(n6032), .B1(n7284), .Y(n5622) );
	mux2i_1 U7581( .A0(n7285), .A1(n7286), .S(n7287), .Y(n7284) );
	and2_0 U7582( .A(n10362), .B(n7288), .X(n7287) );
	nor2_1 U7583( .A(n6293), .B(n6031), .Y(n7285) );
	o21ai_0 U7584( .A1(n6229), .A2(n6790), .B1(n7289), .Y(n5621) );
	mux2i_1 U7585( .A0(n7290), .A1(n6251), .S(n7291), .Y(n7289) );
	nor2_1 U7586( .A(n6491), .B(n6870), .Y(n7291) );
	nor2_1 U7587( .A(n6293), .B(n5993), .Y(n7290) );
	inv_1 U7588( .A(n10799), .Y(n6790) );
	o21ai_0 U7589( .A1(n6229), .A2(n6045), .B1(n7292), .Y(n5620) );
	mux2i_1 U7590( .A0(n7293), .A1(n7294), .S(n10323), .Y(n7292) );
	nor2_1 U7591( .A(n6293), .B(n7295), .Y(n7293) );
	o22ai_1 U7592( .A1(n6205), .A2(n7296), .B1(n7297), .B2(n6295), .Y(n5619) );
	nor3_1 U7593( .A(n7298), .B(n10452), .C(n7299), .Y(n7297) );
	nor2_1 U7594( .A(n6360), .B(n7300), .Y(n5618) );
	o21ai_0 U7595( .A1(n6229), .A2(n5997), .B1(n7301), .Y(n5617) );
	mux2i_1 U7596( .A0(n7302), .A1(n7303), .S(n7304), .Y(n7301) );
	nor2_1 U7597( .A(n7305), .B(n7306), .Y(n7304) );
	nor2_1 U7598( .A(n6283), .B(n7307), .Y(n7302) );
	o21ai_0 U7599( .A1(n6045), .A2(n7308), .B1(n7309), .Y(n5616) );
	mux2i_1 U7600( .A0(n7310), .A1(n7311), .S(n7312), .Y(n7309) );
	nor3_1 U7601( .A(n7295), .B(n10695), .C(n6307), .Y(n7311) );
	inv_1 U7602( .A(n7313), .Y(n7295) );
	nand2_1 U7603( .A(n6224), .B(n7314), .Y(n7310) );
	nand3_1 U7604( .A(n7313), .B(n6374), .C(n10695), .Y(n7314) );
	o22ai_1 U7605( .A1(n6204), .A2(n7315), .B1(n7316), .B2(n6294), .Y(n5615) );
	nor2_1 U7606( .A(n11936), .B(n7317), .Y(n7316) );
	o21ai_0 U7607( .A1(n6230), .A2(n5971), .B1(n7318), .Y(n5614) );
	mux2i_1 U7608( .A0(n7319), .A1(n6251), .S(n7320), .Y(n7318) );
	nor2_1 U7609( .A(n7071), .B(n7321), .Y(n7320) );
	nor2_1 U7610( .A(n6283), .B(n6660), .Y(n7319) );
	inv_1 U7611( .A(n10499), .Y(n6660) );
	and2_0 U7612( .A(n6386), .B(g8403), .X(n5613) );
	o21ai_0 U7613( .A1(n6230), .A2(n7322), .B1(n7323), .Y(n5612) );
	mux2i_1 U7614( .A0(n7324), .A1(n6251), .S(n7325), .Y(n7323) );
	nor2_1 U7615( .A(n6282), .B(n7326), .Y(n7324) );
	o21ai_0 U7616( .A1(n6230), .A2(n7327), .B1(n7328), .Y(n5611) );
	mux2i_1 U7617( .A0(n7329), .A1(n6252), .S(n7330), .Y(n7328) );
	nor2_1 U7618( .A(n7331), .B(n7332), .Y(n7330) );
	nor2_1 U7619( .A(n6280), .B(n7333), .Y(n7329) );
	o21ai_0 U7620( .A1(n6230), .A2(n7334), .B1(n7335), .Y(n5610) );
	mux2i_1 U7621( .A0(n7336), .A1(n7337), .S(n7338), .Y(n7335) );
	and2_0 U7622( .A(n7339), .B(n7340), .X(n7337) );
	nor2_1 U7623( .A(n7340), .B(n7341), .Y(n7336) );
	o21ai_0 U7624( .A1(n6230), .A2(n7159), .B1(n7342), .Y(n5609) );
	a22oi_1 U7625( .A1(n11770), .A2(n7294), .B1(n7313), .B2(n6430), .Y(n7342) );
	inv_1 U7626( .A(n7308), .Y(n7294) );
	o21ai_0 U7627( .A1(n6230), .A2(n5991), .B1(n7343), .Y(n5608) );
	mux2i_1 U7628( .A0(n7344), .A1(n7345), .S(n7346), .Y(n7343) );
	nor3_1 U7629( .A(n7030), .B(n7347), .C(n7038), .Y(n7346) );
	nor2_1 U7630( .A(n6280), .B(n7348), .Y(n7344) );
	o21ai_0 U7631( .A1(n6231), .A2(n7349), .B1(n7350), .Y(n5607) );
	mux2i_1 U7632( .A0(n7351), .A1(n6252), .S(n7352), .Y(n7350) );
	nor2_1 U7633( .A(n7353), .B(n7331), .Y(n7352) );
	nor2_1 U7634( .A(n6279), .B(n7354), .Y(n7351) );
	o221ai_1 U7635( .A1(n6035), .A2(n7074), .B1(n7355), .B2(n7356), .C1(n7357), .Y(n5606) );
	a22oi_1 U7636( .A1(n10547), .A2(n7358), .B1(n10337), .B2(n6437), .Y(n7357) );
	inv_1 U7637( .A(n6590), .Y(n7356) );
	a221oi_1 U7638( .A1(n10725), .A2(n7359), .B1(n11854), .B2(n7360), .C1(n7361), .Y(n7355) );
	o32ai_1 U7639( .A1(n7362), .A2(n11958), .A3(n10337), .B1(n10176), .B2(n7363), .Y(n7361) );
	a22oi_1 U7640( .A1(n11855), .A2(n10337), .B1(n11848), .B2(n11958), .Y(n7363) );
	o21ai_0 U7641( .A1(n6231), .A2(n6543), .B1(n7364), .Y(n5605) );
	mux2i_1 U7642( .A0(n7365), .A1(n6252), .S(n7366), .Y(n7364) );
	nor2_1 U7643( .A(n6466), .B(n6501), .Y(n7366) );
	nor2_1 U7644( .A(n6279), .B(n6006), .Y(n7365) );
	o21ai_0 U7645( .A1(n6231), .A2(n7367), .B1(n7368), .Y(n5604) );
	a22oi_1 U7646( .A1(n10329), .A2(n7369), .B1(n11937), .B2(n7370), .Y(n7368) );
	o21ai_0 U7647( .A1(n7075), .A2(n6094), .B1(n7371), .Y(n5603) );
	mux2i_1 U7648( .A0(n7372), .A1(n7373), .S(n7374), .Y(n7371) );
	nor2_1 U7649( .A(n10324), .B(n7074), .Y(n7373) );
	nand2_1 U7650( .A(n7375), .B(n6334), .Y(n7074) );
	nand2_1 U7651( .A(n6223), .B(n7376), .Y(n7372) );
	o32ai_1 U7652( .A1(n6311), .A2(n10416), .A3(n6495), .B1(n6201), .B2(n7377), .Y(n5602) );
	nor2_1 U7653( .A(n7377), .B(n7378), .Y(n6495) );
	o22ai_1 U7654( .A1(n6204), .A2(n7379), .B1(n7380), .B2(n6297), .Y(n5601) );
	xnor2_1 U7655( .A(n7381), .B(n10537), .Y(n7380) );
	o21ai_0 U7656( .A1(n6231), .A2(n7382), .B1(n7383), .Y(n5600) );
	mux2i_1 U7657( .A0(n7384), .A1(n6252), .S(n7385), .Y(n7383) );
	nor2_1 U7658( .A(n6995), .B(n7386), .Y(n7385) );
	nor2_1 U7659( .A(n6279), .B(n5921), .Y(n7384) );
	o22ai_1 U7660( .A1(n6205), .A2(n7387), .B1(n6277), .B2(n7388), .Y(n5599) );
	o22ai_1 U7661( .A1(n10411), .A2(n7389), .B1(n7390), .B2(n7391), .Y(n7388) );
	nor3_1 U7662( .A(n7392), .B(n7393), .C(n7281), .Y(n7389) );
	nor2_1 U7663( .A(n6279), .B(n7394), .Y(n5598) );
	o32ai_1 U7664( .A1(n6057), .A2(n6350), .A3(n7395), .B1(n7396), .B2(n7397), .Y(n5597) );
	o21ai_0 U7665( .A1(n6232), .A2(n6711), .B1(n7398), .Y(n5596) );
	mux2i_1 U7666( .A0(n7399), .A1(n7400), .S(n7401), .Y(n7398) );
	nor2_1 U7667( .A(n7402), .B(n7130), .Y(n7400) );
	nor2_1 U7668( .A(n6280), .B(n7403), .Y(n7399) );
	o22ai_1 U7669( .A1(n6305), .A2(n7404), .B1(n6194), .B2(n6937), .Y(n5595) );
	mux2i_1 U7670( .A0(n7405), .A1(n7406), .S(n7407), .Y(n5594) );
	nand2_1 U7671( .A(n7408), .B(n10202), .Y(n7406) );
	a21oi_1 U7672( .A1(n7409), .A2(n7410), .B1(n6437), .Y(n7405) );
	nor2_1 U7673( .A(n6360), .B(n7411), .Y(n5593) );
	o32ai_1 U7674( .A1(n7412), .A2(n7142), .A3(n7413), .B1(n6367), .B2(n6078), .Y(n5592) );
	o22ai_1 U7675( .A1(n6204), .A2(n7414), .B1(n7415), .B2(n6298), .Y(n5591) );
	nor2_1 U7676( .A(n7416), .B(n7417), .Y(n7415) );
	xnor2_1 U7677( .A(n7418), .B(n7419), .Y(n7417) );
	o32ai_1 U7678( .A1(n6062), .A2(n7420), .A3(n6313), .B1(n7421), .B2(n7422), .Y(n5590) );
	nor2_1 U7679( .A(n7423), .B(n6437), .Y(n7421) );
	nor4_1 U7680( .A(n11939), .B(n6367), .C(n7424), .D(n7425), .Y(n7423) );
	a21oi_1 U7681( .A1(n10518), .A2(n7422), .B1(n7425), .Y(n7420) );
	inv_1 U7682( .A(n10423), .Y(n7422) );
	o32ai_1 U7683( .A1(n7426), .A2(n10259), .A3(n7036), .B1(n7030), .B2(n7427), .Y(n5589) );
	o21ai_0 U7684( .A1(n10238), .A2(n7428), .B1(n6343), .Y(n7426) );
	o221ai_1 U7685( .A1(n7429), .A2(n7430), .B1(n6215), .B2(n5969), .C1(n7431), .Y(n5588) );
	or4_1 U7686( .A(n7121), .B(n6314), .C(n7432), .D(n7433), .X(n7431) );
	inv_1 U7687( .A(n7434), .Y(n5587) );
	a21oi_1 U7688( .A1(n6620), .A2(n11921), .B1(n7435), .Y(n7434) );
	mux2_1 U7689( .A0(n7436), .A1(n7437), .S(n10631), .X(n7435) );
	nand2_1 U7690( .A(n6223), .B(n6986), .Y(n7437) );
	nand3_1 U7691( .A(n7438), .B(n6375), .C(n10318), .Y(n6986) );
	nor2_1 U7692( .A(n10318), .B(n6623), .Y(n7436) );
	nor2_1 U7693( .A(n6280), .B(n7438), .Y(n6620) );
	o32ai_1 U7694( .A1(n7439), .A2(n7440), .A3(n6313), .B1(n7441), .B2(n5953), .Y(n5586) );
	a21oi_1 U7695( .A1(n7440), .A2(n6381), .B1(n6437), .Y(n7441) );
	and2_0 U7696( .A(n7288), .B(n6641), .X(n7440) );
	nor2_1 U7697( .A(n7442), .B(n10182), .Y(n7288) );
	nor3_1 U7698( .A(n7443), .B(n6350), .C(n7444), .Y(n5585) );
	a21oi_1 U7699( .A1(n10851), .A2(n6750), .B1(n7257), .Y(n7444) );
	nor3_1 U7700( .A(n7445), .B(n7259), .C(n7248), .Y(n7443) );
	o21ai_0 U7701( .A1(n6232), .A2(n5988), .B1(n7446), .Y(n5584) );
	mux2i_1 U7702( .A0(n7447), .A1(n7021), .S(n7448), .Y(n7446) );
	nor2_1 U7703( .A(n7449), .B(n7450), .Y(n7448) );
	nor2_1 U7704( .A(n6280), .B(n7451), .Y(n7447) );
	o21ai_0 U7705( .A1(n6232), .A2(n6964), .B1(n7452), .Y(n5583) );
	mux2i_1 U7706( .A0(n7453), .A1(n7454), .S(n7455), .Y(n7452) );
	and2_0 U7707( .A(n6386), .B(n7456), .X(n7454) );
	nor2_1 U7708( .A(n7456), .B(n6300), .Y(n7453) );
	nor4_1 U7709( .A(n6964), .B(n6970), .C(n6550), .D(n10441), .Y(n7456) );
	inv_1 U7710( .A(n10911), .Y(n6964) );
	o21ai_0 U7711( .A1(n6232), .A2(n5990), .B1(n7457), .Y(n5582) );
	mux2i_1 U7712( .A0(n7458), .A1(n7118), .S(n7459), .Y(n7457) );
	nor2_1 U7713( .A(n7120), .B(n7460), .Y(n7459) );
	inv_1 U7714( .A(n7461), .Y(n7120) );
	nor2_1 U7715( .A(n6281), .B(n7462), .Y(n7458) );
	o32ai_1 U7716( .A1(n7463), .A2(n6350), .A3(n7464), .B1(n7465), .B2(n7466), .Y(n5581) );
	o32ai_1 U7717( .A1(n6311), .A2(n10179), .A3(n7467), .B1(n6201), .B2(n7468), .Y(n5580) );
	xnor2_1 U7718( .A(n7469), .B(n10346), .Y(n7467) );
	o22ai_1 U7719( .A1(n6484), .A2(n6202), .B1(n6304), .B2(n7470), .Y(n5579) );
	mux2i_1 U7720( .A0(n10467), .A1(n10456), .S(n7471), .Y(n7470) );
	nor2_1 U7721( .A(n7281), .B(n7472), .Y(n7471) );
	o32ai_1 U7722( .A1(n6311), .A2(n10413), .A3(n7473), .B1(n6201), .B2(n7474), .Y(n5578) );
	o21ai_0 U7723( .A1(n6891), .A2(n7475), .B1(n7476), .Y(n5577) );
	mux2i_1 U7724( .A0(n7477), .A1(n7478), .S(n10554), .Y(n7476) );
	nand2_1 U7725( .A(n6223), .B(n7479), .Y(n7478) );
	nand3_1 U7726( .A(n7480), .B(n6374), .C(n7102), .Y(n7479) );
	nor2_1 U7727( .A(n6281), .B(n7480), .Y(n7477) );
	nand2_1 U7728( .A(n10678), .B(n7481), .Y(n7480) );
	o21ai_0 U7729( .A1(n6232), .A2(n6682), .B1(n7482), .Y(n5576) );
	mux2i_1 U7730( .A0(n7483), .A1(n6252), .S(n7484), .Y(n7482) );
	nor2_1 U7731( .A(n6680), .B(n7485), .Y(n7484) );
	nor2_1 U7732( .A(n6281), .B(n5976), .Y(n7483) );
	o221ai_1 U7733( .A1(n7486), .A2(n7487), .B1(n6216), .B2(n6074), .C1(n7488), .Y(n5575) );
	nand3_1 U7734( .A(n6340), .B(n7489), .C(n7490), .Y(n7488) );
	o21ai_0 U7735( .A1(n6233), .A2(n7059), .B1(n7491), .Y(n5574) );
	inv_1 U7736( .A(n7492), .Y(n7491) );
	o22ai_1 U7737( .A1(n7061), .A2(n7060), .B1(n5950), .B2(n6630), .Y(n7492) );
	inv_1 U7738( .A(n10857), .Y(n7059) );
	o22ai_1 U7739( .A1(n6305), .A2(n5872), .B1(n6194), .B2(n5955), .Y(n5573) );
	o21ai_0 U7740( .A1(n6225), .A2(n5928), .B1(n7493), .Y(n5572) );
	mux2i_1 U7741( .A0(n7494), .A1(n6252), .S(n7495), .Y(n7493) );
	nor2_1 U7742( .A(n6628), .B(n7496), .Y(n7495) );
	nor2_1 U7743( .A(n6281), .B(n7497), .Y(n7494) );
	o21ai_0 U7744( .A1(n5947), .A2(n7182), .B1(n7498), .Y(n5571) );
	mux2i_1 U7745( .A0(n7499), .A1(n7500), .S(n10900), .Y(n7498) );
	nand2_1 U7746( .A(n6222), .B(n7501), .Y(n7500) );
	nand3_1 U7747( .A(n6381), .B(n6697), .C(n7502), .Y(n7501) );
	nor2_1 U7748( .A(n6697), .B(n7181), .Y(n7499) );
	o21ai_0 U7749( .A1(n6233), .A2(n6900), .B1(n7503), .Y(n5570) );
	mux2i_1 U7750( .A0(n7504), .A1(n6255), .S(n7505), .Y(n7503) );
	nor2_1 U7751( .A(n6899), .B(n7506), .Y(n7505) );
	nor2_1 U7752( .A(n6282), .B(n5922), .Y(n7504) );
	o22ai_1 U7753( .A1(n7507), .A2(n7508), .B1(n7509), .B2(n7510), .Y(n5569) );
	a21oi_1 U7754( .A1(n7511), .A2(n10621), .B1(n6437), .Y(n7509) );
	nor2_1 U7755( .A(n10571), .B(n7512), .Y(n7511) );
	a21oi_1 U7756( .A1(n7513), .A2(n7510), .B1(n62), .Y(n7507) );
	o22ai_1 U7757( .A1(n6205), .A2(n7514), .B1(n7515), .B2(n6297), .Y(n5568) );
	o22ai_1 U7758( .A1(n7516), .A2(n6302), .B1(n7517), .B2(n7038), .Y(n5567) );
	a21oi_1 U7759( .A1(n7518), .A2(n10478), .B1(n6437), .Y(n7517) );
	nor2_1 U7760( .A(n6361), .B(n7519), .Y(n7518) );
	a22oi_1 U7761( .A1(n7519), .A2(n7520), .B1(n10478), .B2(n7521), .Y(n7516) );
	o21ai_0 U7762( .A1(n7030), .A2(n7519), .B1(n7522), .Y(n7521) );
	o21ai_0 U7763( .A1(n10478), .A2(n7347), .B1(n7523), .Y(n7520) );
	mux2_1 U7764( .A0(n7524), .A1(n10688), .S(n7525), .X(n7519) );
	nand2_1 U7765( .A(n7526), .B(n7527), .Y(n7524) );
	o32ai_1 U7766( .A1(n7528), .A2(n6349), .A3(n7529), .B1(n7530), .B2(n7018), .Y(n5566) );
	o221ai_1 U7767( .A1(n7531), .A2(n7532), .B1(n6216), .B2(n7533), .C1(n7534), .Y(n5565) );
	nand3_1 U7768( .A(n6340), .B(n7535), .C(n10522), .Y(n7534) );
	o21ai_0 U7769( .A1(n6917), .A2(n7536), .B1(n7537), .Y(n7532) );
	o21ai_0 U7770( .A1(n6233), .A2(n7538), .B1(n7539), .Y(n5564) );
	mux2i_1 U7771( .A0(n7540), .A1(n7541), .S(n7542), .Y(n7539) );
	nor2_1 U7772( .A(n7543), .B(n7544), .Y(n7540) );
	o22ai_1 U7773( .A1(n6810), .A2(n7545), .B1(n6811), .B2(n7546), .Y(n5563) );
	o22ai_1 U7774( .A1(n6071), .A2(n6784), .B1(n7547), .B2(n7548), .Y(n5562) );
	inv_1 U7775( .A(n10931), .Y(n7548) );
	a21oi_1 U7776( .A1(n6782), .A2(n7549), .B1(n6437), .Y(n7547) );
	o21ai_0 U7777( .A1(n6233), .A2(n7550), .B1(n7551), .Y(n5561) );
	a22oi_1 U7778( .A1(n7136), .A2(n7552), .B1(n10735), .B2(n7138), .Y(n7551) );
	o32ai_1 U7779( .A1(n7553), .A2(n7554), .A3(n6313), .B1(n7555), .B2(n7556), .Y(n5560) );
	a21oi_1 U7780( .A1(n7557), .A2(n7554), .B1(n6437), .Y(n7555) );
	nor2_1 U7781( .A(n10405), .B(n6363), .Y(n7557) );
	o32ai_1 U7782( .A1(n6871), .A2(n10159), .A3(n6492), .B1(n6202), .B2(n5903), .Y(n5559) );
	inv_1 U7783( .A(n7558), .Y(n6871) );
	o21ai_0 U7784( .A1(n6232), .A2(n6026), .B1(n7559), .Y(n5558) );
	mux2i_1 U7785( .A0(n7560), .A1(n6559), .S(n7561), .Y(n7559) );
	nor2_1 U7786( .A(n10265), .B(n7562), .Y(n7561) );
	nor2_1 U7787( .A(n6281), .B(n5989), .Y(n7560) );
	o21ai_0 U7788( .A1(n6232), .A2(n7563), .B1(n7564), .Y(n5557) );
	a22oi_1 U7789( .A1(n7565), .A2(n11772), .B1(n7566), .B2(n7118), .Y(n7564) );
	o21ai_0 U7790( .A1(n6232), .A2(n5992), .B1(n7567), .Y(n5556) );
	mux2i_1 U7791( .A0(n7568), .A1(n6252), .S(n7569), .Y(n7567) );
	nor2_1 U7792( .A(n7570), .B(n6868), .Y(n7569) );
	nor2_1 U7793( .A(n6282), .B(n5999), .Y(n7568) );
	o32ai_1 U7794( .A1(n7571), .A2(n7572), .A3(n6312), .B1(n7573), .B2(n5932), .Y(n5555) );
	o221ai_1 U7795( .A1(n7574), .A2(n5963), .B1(n10335), .B2(n7101), .C1(n7575), .Y(n5554) );
	mux2i_1 U7796( .A0(n7576), .A1(n7577), .S(n7100), .Y(n7575) );
	nor4_1 U7797( .A(n6744), .B(n7578), .C(n6890), .D(n7579), .Y(n7577) );
	nand2_1 U7798( .A(n6222), .B(n7101), .Y(n7576) );
	inv_1 U7799( .A(n6893), .Y(n7101) );
	a211oi_1 U7800( .A1(n6330), .A2(n7579), .B1(n6746), .C1(n6848), .Y(n7574) );
	o221ai_1 U7801( .A1(n7580), .A2(n6309), .B1(n7544), .B2(n7581), .C1(n7582), .Y(n5553) );
	o21ai_0 U7802( .A1(n6437), .A2(n64), .B1(n11861), .Y(n7582) );
	inv_1 U7803( .A(n7583), .Y(n7580) );
	o21ai_0 U7804( .A1(g12923), .A2(n11861), .B1(g19357), .Y(n7583) );
	o221ai_1 U7805( .A1(n6764), .A2(n7584), .B1(n6215), .B2(n5873), .C1(n7585), .Y(n5552) );
	a21oi_1 U7806( .A1(n7586), .A2(n10173), .B1(n7587), .Y(n7585) );
	o21ai_0 U7807( .A1(n6231), .A2(n7588), .B1(n7589), .Y(n5551) );
	mux2i_1 U7808( .A0(n7590), .A1(n7591), .S(n7592), .Y(n7589) );
	nor2_1 U7809( .A(n10394), .B(n6364), .Y(n7591) );
	nor2_1 U7810( .A(n7108), .B(n7593), .Y(n7590) );
	o221ai_1 U7811( .A1(n7594), .A2(n7595), .B1(n6215), .B2(n7596), .C1(n7597), .Y(n5550) );
	o21ai_0 U7812( .A1(n7598), .A2(n6746), .B1(n11866), .Y(n7597) );
	a21oi_1 U7813( .A1(g27831), .A2(n7599), .B1(n6314), .Y(n7598) );
	nand2_1 U7814( .A(g27831), .B(n7599), .Y(n7595) );
	mux2i_1 U7815( .A0(n7600), .A1(n7601), .S(n7602), .Y(n7594) );
	and2_0 U7816( .A(n6386), .B(n11944), .X(n5549) );
	o32ai_1 U7817( .A1(n7603), .A2(n6349), .A3(n7604), .B1(n7605), .B2(n7606), .Y(n5548) );
	inv_1 U7818( .A(n10694), .Y(n7603) );
	o21ai_0 U7819( .A1(n6231), .A2(n7607), .B1(n7608), .Y(n5547) );
	mux2i_1 U7820( .A0(n7609), .A1(n6252), .S(n7610), .Y(n7608) );
	nor2_1 U7821( .A(n7229), .B(n7611), .Y(n7610) );
	nor2_1 U7822( .A(n6282), .B(n5924), .Y(n7609) );
	o21ai_0 U7823( .A1(n6231), .A2(n7612), .B1(n7613), .Y(n5546) );
	mux2i_1 U7824( .A0(n7614), .A1(n7615), .S(n7616), .Y(n7613) );
	nor3_1 U7825( .A(n7617), .B(n10246), .C(n6368), .Y(n7615) );
	nor2_1 U7826( .A(n7618), .B(n6564), .Y(n7614) );
	o21ai_0 U7827( .A1(n6231), .A2(n6031), .B1(n7619), .Y(n5545) );
	mux2i_1 U7828( .A0(n7620), .A1(n7286), .S(n7621), .Y(n7619) );
	nor2_1 U7829( .A(n6645), .B(n7442), .Y(n7621) );
	nor2_1 U7830( .A(n6282), .B(n5952), .Y(n7620) );
	o221ai_1 U7831( .A1(n6623), .A2(n6027), .B1(n7622), .B2(n7623), .C1(n7624), .Y(n5544) );
	a22oi_1 U7832( .A1(n10553), .A2(n7625), .B1(n10331), .B2(n6437), .Y(n7624) );
	inv_1 U7833( .A(n7626), .Y(n7623) );
	a221oi_1 U7834( .A1(n7627), .A2(n11782), .B1(n7628), .B2(n11853), .C1(n7629), .Y(n7622) );
	o32ai_1 U7835( .A1(n7630), .A2(n11946), .A3(n10331), .B1(n10299), .B2(n7631), .Y(n7629) );
	a22oi_1 U7836( .A1(n10331), .A2(n11792), .B1(n11813), .B2(n11946), .Y(n7631) );
	nand2_1 U7837( .A(n7438), .B(n6334), .Y(n6623) );
	nor3_1 U7838( .A(n7632), .B(n7633), .C(n5894), .Y(n7438) );
	o22ai_1 U7839( .A1(n6206), .A2(n6637), .B1(n7634), .B2(n6396), .Y(n5543) );
	xnor2_1 U7840( .A(n10235), .B(n7635), .Y(n7634) );
	o21ai_0 U7841( .A1(n7162), .A2(n7636), .B1(n7637), .Y(n5542) );
	mux2i_1 U7842( .A0(n7638), .A1(n7639), .S(n10642), .Y(n7637) );
	nand2_1 U7843( .A(n6221), .B(n7165), .Y(n7639) );
	nand3_1 U7844( .A(n7640), .B(n6375), .C(n10684), .Y(n7165) );
	nor2_1 U7845( .A(n10684), .B(n7641), .Y(n7638) );
	o21ai_0 U7846( .A1(n6231), .A2(n6050), .B1(n7642), .Y(n5541) );
	mux2i_1 U7847( .A0(n7020), .A1(n7643), .S(n7644), .Y(n7642) );
	nor2_1 U7848( .A(n6282), .B(n7645), .Y(n7643) );
	inv_1 U7849( .A(n7530), .Y(n7020) );
	o21ai_0 U7850( .A1(n7646), .A2(n6048), .B1(n7647), .Y(n5540) );
	mux2i_1 U7851( .A0(n7648), .A1(n7649), .S(n7650), .Y(n7647) );
	nor3_1 U7852( .A(n7651), .B(n10690), .C(n6306), .Y(n7649) );
	nand2_1 U7853( .A(n6221), .B(n7652), .Y(n7648) );
	nand3_1 U7854( .A(n10690), .B(n6375), .C(n7653), .Y(n7652) );
	o221ai_1 U7855( .A1(n5893), .A2(n6891), .B1(n6214), .B2(n7654), .C1(n7655), .Y(n5539) );
	a21oi_1 U7856( .A1(n7656), .A2(n6849), .B1(n6893), .Y(n7655) );
	nor3_1 U7857( .A(n7578), .B(n7657), .C(n7579), .Y(n6893) );
	nor2_1 U7858( .A(n10335), .B(n6851), .Y(n7656) );
	inv_1 U7859( .A(n6848), .Y(n6891) );
	o221ai_1 U7860( .A1(n6446), .A2(n6028), .B1(n7658), .B2(n7659), .C1(n7660), .Y(n5538) );
	a22oi_1 U7861( .A1(n10548), .A2(n7661), .B1(n10292), .B2(n6437), .Y(n7660) );
	inv_1 U7862( .A(n7662), .Y(n7659) );
	a221oi_1 U7863( .A1(n10738), .A2(n7663), .B1(n10930), .B2(g25167), .C1( n7664), .Y(n7658) );
	o32ai_1 U7864( .A1(n7307), .A2(n11953), .A3(n10292), .B1(n10301), .B2(n7665), .Y(n7664) );
	a22oi_1 U7865( .A1(n11830), .A2(n10292), .B1(n11820), .B2(n11953), .Y(n7665) );
	o22ai_1 U7866( .A1(n6206), .A2(n7410), .B1(n7666), .B2(n7667), .Y(n5537) );
	a211oi_1 U7867( .A1(n10349), .A2(n7407), .B1(n7668), .C1(n7325), .Y(n7666) );
	nor2_1 U7868( .A(n7669), .B(n7407), .Y(n7325) );
	nor2_1 U7869( .A(n6282), .B(n6974), .Y(n5536) );
	o21ai_0 U7870( .A1(n6230), .A2(n7670), .B1(n7671), .Y(n5535) );
	a22oi_1 U7871( .A1(n7672), .A2(n7048), .B1(n10899), .B2(n7046), .Y(n7671) );
	nor2_1 U7872( .A(n6283), .B(n6932), .Y(n7046) );
	nor2_1 U7873( .A(n6936), .B(n6301), .Y(n7048) );
	xnor2_1 U7874( .A(n7673), .B(n7205), .Y(n7672) );
	nand2_1 U7875( .A(n7674), .B(n7675), .Y(n7205) );
	mux2i_1 U7876( .A0(n7676), .A1(n7677), .S(n7678), .Y(n7675) );
	xnor2_1 U7877( .A(n7377), .B(g12300), .Y(n7678) );
	nand3_1 U7878( .A(n7679), .B(n7680), .C(n7681), .Y(n7677) );
	nand3_1 U7879( .A(n11783), .B(g17711), .C(n6930), .Y(n7681) );
	nand3_1 U7880( .A(n11812), .B(g14694), .C(n7682), .Y(n7680) );
	nand3_1 U7881( .A(g17580), .B(n10496), .C(n7683), .Y(n7679) );
	nand3_1 U7882( .A(n7684), .B(n7685), .C(n7686), .Y(n7676) );
	nand3_1 U7883( .A(n7687), .B(g17711), .C(n11951), .Y(n7686) );
	nand3_1 U7884( .A(n7682), .B(g17580), .C(n10790), .Y(n7685) );
	nand3_1 U7885( .A(n7683), .B(g14694), .C(n11952), .Y(n7684) );
	inv_1 U7886( .A(n6933), .Y(n7683) );
	mux2_1 U7887( .A0(n7688), .A1(n7689), .S(n7377), .X(n7674) );
	a221oi_1 U7888( .A1(n6930), .A2(n7690), .B1(n7687), .B2(n7691), .C1(n7692), .Y(n7689) );
	o32ai_1 U7889( .A1(n7693), .A2(n5925), .A3(n7694), .B1(n7695), .B2(n6933), .Y(n7692) );
	a22oi_1 U7890( .A1(n10778), .A2(g13049), .B1(n10779), .B2(n10224), .Y(n7695) );
	o22ai_1 U7891( .A1(n6664), .A2(n7696), .B1(n7697), .B2(n7698), .Y(n7691) );
	o22ai_1 U7892( .A1(n7699), .A2(n7700), .B1(n7701), .B2(n7702), .Y(n7690) );
	a221oi_1 U7893( .A1(n6930), .A2(n7703), .B1(n7687), .B2(n7704), .C1(n7705), .Y(n7688) );
	o32ai_1 U7894( .A1(n5938), .A2(n6933), .A3(n7693), .B1(n7706), .B2(n7694), .Y(n7705) );
	a22oi_1 U7895( .A1(n10788), .A2(g13049), .B1(n10789), .B2(n10224), .Y(n7706) );
	o22ai_1 U7896( .A1(n7699), .A2(n7707), .B1(n7203), .B2(n7701), .Y(n7704) );
	inv_1 U7897( .A(n10784), .Y(n7203) );
	o22ai_1 U7898( .A1(n7696), .A2(n7708), .B1(n7697), .B2(n7709), .Y(n7703) );
	nand2_1 U7899( .A(n10899), .B(n7710), .Y(n7673) );
	o32ai_1 U7900( .A1(n6311), .A2(g9553), .A3(n7711), .B1(n6202), .B2(n7712), .Y(n5534) );
	a21oi_1 U7901( .A1(g9497), .A2(n7712), .B1(n10151), .Y(n7711) );
	inv_1 U7902( .A(n10614), .Y(n7712) );
	o221ai_1 U7903( .A1(n5891), .A2(n6706), .B1(n6213), .B2(n7713), .C1(n7714), .Y(n5533) );
	a21oi_1 U7904( .A1(n7715), .A2(n7662), .B1(n7716), .Y(n7714) );
	nor2_1 U7905( .A(n10292), .B(n7663), .Y(n7715) );
	o221ai_1 U7906( .A1(n7717), .A2(n5965), .B1(n10336), .B2(n7718), .C1(n7719), .Y(n5532) );
	mux2i_1 U7907( .A0(n7720), .A1(n7721), .S(n7722), .Y(n7719) );
	nor4_1 U7908( .A(n7222), .B(n7723), .C(n6744), .D(n7724), .Y(n7721) );
	nand2_1 U7909( .A(n6220), .B(n7718), .Y(n7720) );
	a211oi_1 U7910( .A1(n6330), .A2(n7724), .B1(n7161), .C1(n6746), .Y(n7717) );
	and2_0 U7911( .A(n6385), .B(g8291), .X(n5531) );
	o22ai_1 U7912( .A1(n6206), .A2(n7725), .B1(n7726), .B2(n6734), .Y(n5530) );
	xnor2_1 U7913( .A(n11954), .B(n7727), .Y(n7726) );
	o21ai_0 U7914( .A1(n6230), .A2(n6907), .B1(n7728), .Y(n5529) );
	mux2i_1 U7915( .A0(n7729), .A1(n6252), .S(n7730), .Y(n7728) );
	nor2_1 U7916( .A(n6905), .B(n7731), .Y(n7730) );
	nor2_1 U7917( .A(n6282), .B(n5979), .Y(n7729) );
	inv_1 U7918( .A(n10773), .Y(n6907) );
	o21ai_0 U7919( .A1(n6230), .A2(n7732), .B1(n7733), .Y(n5528) );
	mux2i_1 U7920( .A0(n7734), .A1(n7735), .S(n7736), .Y(n7733) );
	nor2_1 U7921( .A(n6361), .B(n7737), .Y(n7735) );
	and2_0 U7922( .A(n7737), .B(n6345), .X(n7734) );
	o32ai_1 U7923( .A1(n7738), .A2(n6349), .A3(n7395), .B1(n7396), .B2(n7739), .Y(n5527) );
	o21ai_0 U7924( .A1(n7596), .A2(n7486), .B1(n7740), .Y(n5526) );
	nand4_1 U7925( .A(n6339), .B(n7741), .C(n7489), .D(n7305), .Y(n7740) );
	o21ai_0 U7926( .A1(n7742), .A2(n10286), .B1(n7596), .Y(n7741) );
	o221ai_1 U7927( .A1(n6810), .A2(n7743), .B1(n6213), .B2(n7744), .C1(n7745), .Y(n5525) );
	nand3_1 U7928( .A(n7746), .B(n6535), .C(n10870), .Y(n7745) );
	o21ai_0 U7929( .A1(n6229), .A2(n7747), .B1(n7748), .Y(n5524) );
	mux2i_1 U7930( .A0(n7749), .A1(n6252), .S(n7750), .Y(n7748) );
	nor2_1 U7931( .A(n7015), .B(n7072), .Y(n7750) );
	nor2_1 U7932( .A(n6283), .B(n5929), .Y(n7749) );
	o221ai_1 U7933( .A1(n7751), .A2(n5942), .B1(n6212), .B2(n7752), .C1(n7753), .Y(n5523) );
	nand3_1 U7934( .A(n6590), .B(n7754), .C(n7360), .Y(n7753) );
	xnor2_1 U7935( .A(n7018), .B(n10680), .Y(n7754) );
	inv_1 U7936( .A(n10732), .Y(n7018) );
	a21oi_1 U7937( .A1(n6332), .A2(n7755), .B1(n7358), .Y(n7751) );
	o32ai_1 U7938( .A1(n7756), .A2(n6349), .A3(n7757), .B1(n7758), .B2(n7563), .Y(n5522) );
	o221ai_1 U7939( .A1(n7460), .A2(n7429), .B1(n6212), .B2(n7430), .C1(n7759), .Y(n5521) );
	or3_1 U7940( .A(n7432), .B(n6369), .C(n7760), .X(n7759) );
	o21ai_0 U7941( .A1(n6229), .A2(n7761), .B1(n7762), .Y(n5520) );
	mux2i_1 U7942( .A0(n7763), .A1(n7764), .S(n6966), .Y(n7762) );
	nor2_1 U7943( .A(n6360), .B(n7765), .Y(n7764) );
	and2_0 U7944( .A(n7765), .B(n6345), .X(n7763) );
	nand3_1 U7945( .A(n10912), .B(n7766), .C(n7767), .Y(n7765) );
	inv_1 U7946( .A(n10912), .Y(n7761) );
	o221ai_1 U7947( .A1(n7768), .A2(n7769), .B1(n6216), .B2(n7770), .C1(n7771), .Y(n5519) );
	nand3_1 U7948( .A(n7772), .B(n6330), .C(n10329), .Y(n7771) );
	nor2_1 U7949( .A(n6360), .B(n7773), .Y(n5518) );
	o22ai_1 U7950( .A1(n6630), .A2(n7774), .B1(n7775), .B2(n7061), .Y(n5517) );
	nand2_1 U7951( .A(n7776), .B(n6333), .Y(n7061) );
	o22ai_1 U7952( .A1(n6304), .A2(n7777), .B1(n6195), .B2(n7778), .Y(n5516) );
	o21ai_0 U7953( .A1(n6229), .A2(n6493), .B1(n7779), .Y(n5515) );
	mux2i_1 U7954( .A0(n7780), .A1(n6252), .S(n7781), .Y(n7779) );
	nor2_1 U7955( .A(n6283), .B(n7782), .Y(n7780) );
	inv_1 U7956( .A(n10803), .Y(n6493) );
	nor2_1 U7957( .A(n7783), .B(n6301), .Y(n5514) );
	a21oi_1 U7958( .A1(n10556), .A2(n6715), .B1(n7784), .Y(n7783) );
	mux2i_1 U7959( .A0(n7785), .A1(n7786), .S(n6711), .Y(n7784) );
	nand3_1 U7960( .A(n7787), .B(n7403), .C(n7788), .Y(n7786) );
	nand2_1 U7961( .A(n7789), .B(n7790), .Y(n7785) );
	inv_1 U7962( .A(n6716), .Y(n7789) );
	nand2_1 U7963( .A(n7791), .B(n7403), .Y(n6716) );
	inv_1 U7964( .A(n7402), .Y(n7403) );
	o221ai_1 U7965( .A1(n7792), .A2(n5889), .B1(n7793), .B2(n6587), .C1(n7794), .Y(n5513) );
	a21oi_1 U7966( .A1(n7795), .A2(n6381), .B1(n6437), .Y(n7792) );
	o21ai_0 U7967( .A1(n6229), .A2(n7796), .B1(n7797), .Y(n5512) );
	a22oi_1 U7968( .A1(n7136), .A2(n7713), .B1(n10848), .B2(n7138), .Y(n7797) );
	inv_1 U7969( .A(n10586), .Y(n7713) );
	o22ai_1 U7970( .A1(n6304), .A2(n7798), .B1(n6195), .B2(n7799), .Y(n5511) );
	o21ai_0 U7971( .A1(n6229), .A2(n6046), .B1(n7800), .Y(n5510) );
	mux2i_1 U7972( .A0(n7801), .A1(n7802), .S(n10320), .Y(n7800) );
	nor2_1 U7973( .A(n6283), .B(n7803), .Y(n7801) );
	o21ai_0 U7974( .A1(n6228), .A2(n7804), .B1(n7805), .Y(n5509) );
	mux2i_1 U7975( .A0(n7806), .A1(n6252), .S(n7807), .Y(n7805) );
	nor2_1 U7976( .A(n7669), .B(n7331), .Y(n7807) );
	nor2_1 U7977( .A(n6283), .B(n7808), .Y(n7806) );
	o21ai_0 U7978( .A1(n7809), .A2(n6097), .B1(n7810), .Y(n5508) );
	mux2i_1 U7979( .A0(n7811), .A1(n7812), .S(n7813), .Y(n7810) );
	nor2_1 U7980( .A(n10321), .B(n7814), .Y(n7812) );
	nand2_1 U7981( .A(n6222), .B(n7815), .Y(n7811) );
	o21ai_0 U7982( .A1(n6228), .A2(n6021), .B1(n7816), .Y(n5507) );
	mux2i_1 U7983( .A0(n7817), .A1(n7118), .S(n7818), .Y(n7816) );
	nor2_1 U7984( .A(n10261), .B(n7760), .Y(n7818) );
	nor2_1 U7985( .A(n6283), .B(n5990), .Y(n7817) );
	o21ai_0 U7986( .A1(n6228), .A2(n6783), .B1(n7819), .Y(n5506) );
	mux2i_1 U7987( .A0(n7820), .A1(n7821), .S(n7822), .Y(n7819) );
	and2_0 U7988( .A(n7823), .B(n6782), .X(n7821) );
	nor3_1 U7989( .A(n7824), .B(n6350), .C(n7825), .Y(n6782) );
	nor2_1 U7990( .A(n7823), .B(n6784), .Y(n7820) );
	inv_1 U7991( .A(n7826), .Y(n7823) );
	inv_1 U7992( .A(n10462), .Y(n6783) );
	o221ai_1 U7993( .A1(n7827), .A2(n5862), .B1(n10332), .B2(n7828), .C1(n7829), .Y(n5505) );
	mux2i_1 U7994( .A0(n7830), .A1(n7831), .S(n7832), .Y(n7829) );
	nor4_1 U7995( .A(n7833), .B(n7834), .C(n6744), .D(n7835), .Y(n7831) );
	nand2_1 U7996( .A(n6221), .B(n7828), .Y(n7830) );
	a211oi_1 U7997( .A1(n6330), .A2(n7835), .B1(n7836), .C1(n6746), .Y(n7827) );
	o21ai_0 U7998( .A1(n6228), .A2(n6007), .B1(n7837), .Y(n5504) );
	mux2i_1 U7999( .A0(n7838), .A1(n7118), .S(n7839), .Y(n7837) );
	nor3_1 U8000( .A(n7460), .B(n7433), .C(n7121), .Y(n7839) );
	nor2_1 U8001( .A(n6284), .B(n7840), .Y(n7838) );
	o21ai_0 U8002( .A1(n6228), .A2(n7841), .B1(n7842), .Y(n5503) );
	mux2i_1 U8003( .A0(n7843), .A1(n7345), .S(n7844), .Y(n7842) );
	nor2_1 U8004( .A(n10238), .B(n7845), .Y(n7844) );
	nor2_1 U8005( .A(n6284), .B(n5991), .Y(n7843) );
	o21ai_0 U8006( .A1(n6227), .A2(n7846), .B1(n7847), .Y(n5502) );
	mux2i_1 U8007( .A0(n7848), .A1(n6252), .S(n7849), .Y(n7847) );
	nor2_1 U8008( .A(n7407), .B(n6899), .Y(n7849) );
	nor2_1 U8009( .A(n6284), .B(n7349), .Y(n7848) );
	nor2_1 U8010( .A(n6359), .B(n7850), .Y(n5501) );
	o21ai_0 U8011( .A1(n7162), .A2(n5879), .B1(n7851), .Y(n5500) );
	mux2i_1 U8012( .A0(n7852), .A1(n7853), .S(n10899), .Y(n7851) );
	nand2_1 U8013( .A(n6221), .B(n7854), .Y(n7853) );
	nand3_1 U8014( .A(n6384), .B(n7670), .C(n7640), .Y(n7854) );
	nor2_1 U8015( .A(n7641), .B(n7670), .Y(n7852) );
	o21ai_0 U8016( .A1(n6227), .A2(n7855), .B1(n7856), .Y(n5499) );
	mux2i_1 U8017( .A0(n7857), .A1(n7858), .S(n7859), .Y(n7856) );
	and2_0 U8018( .A(n10439), .B(n7860), .X(n7859) );
	nor3_1 U8019( .A(n7861), .B(n10520), .C(n7862), .Y(n7858) );
	nor2_1 U8020( .A(n7863), .B(n7864), .Y(n7857) );
	inv_1 U8021( .A(n10520), .Y(n7864) );
	o21ai_0 U8022( .A1(n6227), .A2(n7636), .B1(n7865), .Y(n5498) );
	mux2_1 U8023( .A0(n7641), .A1(n7162), .S(n11880), .X(n7865) );
	or2_0 U8024( .A(n6314), .B(n7640), .X(n7162) );
	nand2_1 U8025( .A(n7640), .B(n6333), .Y(n7641) );
	nor2_1 U8026( .A(n7710), .B(n6936), .Y(n7640) );
	nand3_1 U8027( .A(n7687), .B(n10376), .C(g17604), .Y(n7710) );
	inv_1 U8028( .A(n10217), .Y(n7636) );
	o22ai_1 U8029( .A1(n7510), .A2(n7866), .B1(n7867), .B2(n7868), .Y(n5497) );
	inv_1 U8030( .A(n10621), .Y(n7868) );
	a21oi_1 U8031( .A1(n64), .A2(n7510), .B1(n6437), .Y(n7867) );
	inv_1 U8032( .A(n7512), .Y(n64) );
	inv_1 U8033( .A(n62), .Y(n7866) );
	nor2_1 U8034( .A(n7544), .B(n10621), .Y(n62) );
	inv_1 U8035( .A(n10388), .Y(n7510) );
	o22ai_1 U8036( .A1(n6207), .A2(n5956), .B1(n7869), .B2(n6297), .Y(n5496) );
	a211oi_1 U8037( .A1(n10364), .A2(n7870), .B1(n10660), .C1(n7871), .Y(n7869) );
	and2_0 U8038( .A(n6386), .B(g7540), .X(n5495) );
	o21ai_0 U8039( .A1(n6227), .A2(n5973), .B1(n7872), .Y(n5494) );
	mux2i_1 U8040( .A0(n7873), .A1(n6253), .S(n7874), .Y(n7872) );
	nor2_1 U8041( .A(n7875), .B(n7386), .Y(n7874) );
	nor2_1 U8042( .A(n6284), .B(n5985), .Y(n7873) );
	o21ai_0 U8043( .A1(n6227), .A2(n7876), .B1(n7877), .Y(n5493) );
	mux2i_1 U8044( .A0(n7878), .A1(n6253), .S(n7879), .Y(n7877) );
	nor2_1 U8045( .A(n6627), .B(n7880), .Y(n7879) );
	nor2_1 U8046( .A(n6285), .B(n7881), .Y(n7878) );
	o221ai_1 U8047( .A1(n7089), .A2(n7110), .B1(n6218), .B2(n5866), .C1(n7882), .Y(n5492) );
	or4_1 U8048( .A(n7883), .B(n6313), .C(n7113), .D(n7884), .X(n7882) );
	o221ai_1 U8049( .A1(n7885), .A2(n7886), .B1(n6217), .B2(n7887), .C1(n7888), .Y(n5491) );
	o21ai_0 U8050( .A1(n7889), .A2(n6746), .B1(n11868), .Y(n7888) );
	inv_1 U8051( .A(n7890), .Y(n7889) );
	o21ai_0 U8052( .A1(n7886), .A2(n7891), .B1(n6343), .Y(n7890) );
	a21oi_1 U8053( .A1(n7892), .A2(n7893), .B1(n7894), .Y(n7885) );
	nor4_1 U8054( .A(n10253), .B(n7039), .C(n7891), .D(n7895), .Y(n7894) );
	a21oi_1 U8055( .A1(n10263), .A2(n7221), .B1(n6309), .Y(n7892) );
	nor3_1 U8056( .A(n7896), .B(n10326), .C(n7897), .Y(n5490) );
	a22oi_1 U8057( .A1(n6331), .A2(n10703), .B1(n7898), .B2(n7513), .Y(n7897) );
	o21ai_0 U8058( .A1(n6226), .A2(n7899), .B1(n7900), .Y(n5489) );
	mux2i_1 U8059( .A0(n7901), .A1(n6253), .S(n7902), .Y(n7900) );
	nor2_1 U8060( .A(n6888), .B(n7903), .Y(n7902) );
	nor2_1 U8061( .A(n6285), .B(n7698), .Y(n7901) );
	o211ai_1 U8062( .A1(n7904), .A2(n7905), .B1(n7906), .C1(n6839), .Y(n5488) );
	nand3_1 U8063( .A(n6841), .B(n7907), .C(n11801), .Y(n7906) );
	a21oi_1 U8064( .A1(n7908), .A2(n6843), .B1(n6437), .Y(n7904) );
	o21ai_0 U8065( .A1(n6228), .A2(n7909), .B1(n7910), .Y(n5487) );
	mux2_1 U8066( .A0(n7215), .A1(n7208), .S(n11881), .X(n7910) );
	and2_0 U8067( .A(n6385), .B(g14167), .X(n5486) );
	nor2_1 U8068( .A(n6361), .B(n7911), .Y(n5485) );
	o22ai_1 U8069( .A1(n6203), .A2(n7912), .B1(n7913), .B2(n6298), .Y(n5484) );
	nor2_1 U8070( .A(n10878), .B(n11974), .Y(n7913) );
	o221ai_1 U8071( .A1(n6454), .A2(n6573), .B1(n6220), .B2(n7914), .C1(n7915), .Y(n5483) );
	or3_1 U8072( .A(n6453), .B(n6369), .C(n7916), .X(n7915) );
	nor2_1 U8073( .A(n6361), .B(n7917), .Y(n5482) );
	o22ai_1 U8074( .A1(g23002), .A2(n6302), .B1(n6197), .B2(n6658), .Y(n5481) );
	inv_1 U8075( .A(n10927), .Y(n6658) );
	o221ai_1 U8076( .A1(n6764), .A2(n5890), .B1(n6219), .B2(n7918), .C1(n7919), .Y(n5480) );
	a21oi_1 U8077( .A1(n7920), .A2(n7586), .B1(n7587), .Y(n7919) );
	nor2_1 U8078( .A(n10334), .B(n7921), .Y(n7920) );
	nor2_1 U8079( .A(n6361), .B(n7922), .Y(n5479) );
	o221ai_1 U8080( .A1(n6516), .A2(n6029), .B1(n7923), .B2(n7924), .C1(n7925), .Y(n5478) );
	a22oi_1 U8081( .A1(n10344), .A2(n7836), .B1(n10332), .B2(n6437), .Y(n7925) );
	inv_1 U8082( .A(n6757), .Y(n7924) );
	a221oi_1 U8083( .A1(n7926), .A2(n10720), .B1(n11808), .B2(n6759), .C1(n7927), .Y(n7923) );
	o32ai_1 U8084( .A1(n7348), .A2(n11901), .A3(n10332), .B1(n10171), .B2(n7928), .Y(n7927) );
	a22oi_1 U8085( .A1(n11814), .A2(n10332), .B1(n11797), .B2(n11901), .Y(n7928) );
	nor2_1 U8086( .A(n7929), .B(n6300), .Y(n5477) );
	xor2_1 U8087( .A(n7930), .B(n7931), .X(n7929) );
	xor2_1 U8088( .A(n7932), .B(n7933), .X(n7931) );
	xnor2_1 U8089( .A(n7934), .B(n10302), .Y(n7933) );
	xnor2_1 U8090( .A(n7935), .B(n10459), .Y(n7932) );
	xor2_1 U8091( .A(n7936), .B(n7937), .X(n7930) );
	xnor2_1 U8092( .A(n7938), .B(n10187), .Y(n7937) );
	xnor2_1 U8093( .A(n7939), .B(n7367), .Y(n7936) );
	or2_0 U8094( .A(n7940), .B(n7941), .X(n7939) );
	o21ai_0 U8095( .A1(n6951), .A2(n6042), .B1(n7942), .Y(n5476) );
	mux2i_1 U8096( .A0(n7943), .A1(n7944), .S(n10896), .Y(n7942) );
	nand2_1 U8097( .A(n6222), .B(n7945), .Y(n7944) );
	nand3_1 U8098( .A(n6375), .B(n7739), .C(n7946), .Y(n7945) );
	nor2_1 U8099( .A(n6950), .B(n7739), .Y(n7943) );
	o21ai_0 U8100( .A1(n6226), .A2(n7947), .B1(n7948), .Y(n5475) );
	mux2i_1 U8101( .A0(n7949), .A1(n6253), .S(n7950), .Y(n7948) );
	nor2_1 U8102( .A(n6995), .B(n7485), .Y(n7950) );
	nor2_1 U8103( .A(n6286), .B(n7382), .Y(n7949) );
	o22ai_1 U8104( .A1(n6205), .A2(n7822), .B1(n7951), .B2(n6784), .Y(n5474) );
	xnor2_1 U8105( .A(n10931), .B(n7549), .Y(n7951) );
	o32ai_1 U8106( .A1(n6300), .A2(n7952), .A3(n7953), .B1(n6199), .B2(n7362), .Y(n5473) );
	a21oi_1 U8107( .A1(n7359), .A2(n7795), .B1(n10585), .Y(n7953) );
	nor4_1 U8108( .A(n10243), .B(n7954), .C(n7955), .D(n7956), .Y(n7952) );
	o21ai_0 U8109( .A1(n6226), .A2(n7957), .B1(n7958), .Y(n5472) );
	mux2i_1 U8110( .A0(n7959), .A1(n6253), .S(n7960), .Y(n7958) );
	nor2_1 U8111( .A(n7570), .B(n6870), .Y(n7960) );
	nor2_1 U8112( .A(n6286), .B(n5992), .Y(n7959) );
	o21ai_0 U8113( .A1(n6226), .A2(n7961), .B1(n7962), .Y(n5471) );
	mux2i_1 U8114( .A0(n7963), .A1(n6253), .S(n7964), .Y(n7962) );
	nor2_1 U8115( .A(n6482), .B(n7965), .Y(n7964) );
	nor2_1 U8116( .A(n6286), .B(n7966), .Y(n7963) );
	o22ai_1 U8117( .A1(n6207), .A2(n7967), .B1(n6347), .B2(n7968), .Y(n5470) );
	inv_1 U8118( .A(n10602), .Y(n7967) );
	o32ai_1 U8119( .A1(n7969), .A2(n6278), .A3(n7424), .B1(n7970), .B2(n7971), .Y(n5469) );
	a21oi_1 U8120( .A1(n7972), .A2(n6376), .B1(n6437), .Y(n7970) );
	inv_1 U8121( .A(n7973), .Y(n7969) );
	a21oi_1 U8122( .A1(n7972), .A2(n11939), .B1(n7974), .Y(n7973) );
	o21ai_0 U8123( .A1(n6587), .A2(n7752), .B1(n7975), .Y(n5468) );
	mux2i_1 U8124( .A0(n7976), .A1(n7977), .S(n10547), .Y(n7975) );
	nand2_1 U8125( .A(n6222), .B(n7978), .Y(n7977) );
	nand3_1 U8126( .A(n7979), .B(n6375), .C(n7795), .Y(n7978) );
	nor2_1 U8127( .A(n6287), .B(n7979), .Y(n7976) );
	nand2_1 U8128( .A(n10680), .B(n7755), .Y(n7979) );
	inv_1 U8129( .A(n7360), .Y(n7755) );
	inv_1 U8130( .A(n10680), .Y(n7752) );
	o22ai_1 U8131( .A1(n6304), .A2(n7778), .B1(n6196), .B2(n6728), .Y(n5467) );
	inv_1 U8132( .A(n10864), .Y(n7778) );
	o21ai_0 U8133( .A1(n6225), .A2(n6034), .B1(n7980), .Y(n5466) );
	mux2i_1 U8134( .A0(n7981), .A1(n6430), .S(n7982), .Y(n7980) );
	nor2_1 U8135( .A(n7887), .B(n7983), .Y(n7982) );
	nor2_1 U8136( .A(n6287), .B(n6022), .Y(n7981) );
	o22ai_1 U8137( .A1(n6810), .A2(n7984), .B1(n7546), .B2(n6084), .Y(n5465) );
	o21ai_0 U8138( .A1(n6225), .A2(n7985), .B1(n7986), .Y(n5464) );
	mux2i_1 U8139( .A0(n7987), .A1(n6430), .S(n7988), .Y(n7986) );
	nor2_1 U8140( .A(n10242), .B(n6432), .Y(n7988) );
	nor2_1 U8141( .A(n6287), .B(n6020), .Y(n7987) );
	o21ai_0 U8142( .A1(n6227), .A2(n7989), .B1(n7990), .Y(n5463) );
	mux2i_1 U8143( .A0(n7991), .A1(n6253), .S(n7992), .Y(n7990) );
	nor2_1 U8144( .A(n7407), .B(n7332), .Y(n7992) );
	nor2_1 U8145( .A(n6287), .B(n7804), .Y(n7991) );
	o21ai_0 U8146( .A1(n6225), .A2(n7993), .B1(n7994), .Y(n5462) );
	mux2i_1 U8147( .A0(n7995), .A1(n7996), .S(n7997), .Y(n7994) );
	nor2_1 U8148( .A(n10528), .B(n6363), .Y(n7996) );
	nor2_1 U8149( .A(n7108), .B(n7998), .Y(n7995) );
	o22ai_1 U8150( .A1(n6303), .A2(n7999), .B1(n8000), .B2(n6508), .Y(n5461) );
	nor3_1 U8151( .A(n8001), .B(n4705), .C(n6437), .Y(n8000) );
	a21oi_1 U8152( .A1(n11847), .A2(n10297), .B1(n6368), .Y(n8001) );
	o221ai_1 U8153( .A1(n8002), .A2(n5868), .B1(n6220), .B2(n7475), .C1(n8003), .Y(n5460) );
	nand3_1 U8154( .A(n6851), .B(n8004), .C(n6849), .Y(n8003) );
	nor2_1 U8155( .A(n7578), .B(n6300), .Y(n6849) );
	xnor2_1 U8156( .A(n8005), .B(n10678), .Y(n8004) );
	inv_1 U8157( .A(n10678), .Y(n7475) );
	a21oi_1 U8158( .A1(n6331), .A2(n7481), .B1(n6848), .Y(n8002) );
	nor2_1 U8159( .A(n6287), .B(n7102), .Y(n6848) );
	inv_1 U8160( .A(n6851), .Y(n7481) );
	nor2_1 U8161( .A(n7100), .B(n11950), .Y(n6851) );
	o22ai_1 U8162( .A1(n8006), .A2(n7077), .B1(n8007), .B2(n8008), .Y(n5459) );
	a21oi_1 U8163( .A1(n8009), .A2(n4753), .B1(n6437), .Y(n8007) );
	nor2_1 U8164( .A(n10572), .B(n8010), .Y(n8009) );
	inv_1 U8165( .A(n10572), .Y(n7077) );
	a21oi_1 U8166( .A1(n7083), .A2(n8008), .B1(n85), .Y(n8006) );
	o21ai_0 U8167( .A1(n6226), .A2(n5995), .B1(n8011), .Y(n5458) );
	mux2i_1 U8168( .A0(n8012), .A1(n6559), .S(n8013), .Y(n8011) );
	nor2_1 U8169( .A(n8014), .B(n8015), .Y(n8013) );
	nor2_1 U8170( .A(n6287), .B(n7630), .Y(n8012) );
	o21ai_0 U8171( .A1(n6225), .A2(n5975), .B1(n8016), .Y(n5457) );
	mux2i_1 U8172( .A0(n8017), .A1(n7345), .S(n8018), .Y(n8016) );
	nor2_1 U8173( .A(n7038), .B(n8019), .Y(n8018) );
	nor2_1 U8174( .A(n6287), .B(n7841), .Y(n8017) );
	inv_1 U8175( .A(n10720), .Y(n7841) );
	o21ai_0 U8176( .A1(n6226), .A2(n8020), .B1(n8021), .Y(n5456) );
	inv_1 U8177( .A(n8022), .Y(n8021) );
	o22ai_1 U8178( .A1(n8023), .A2(n8024), .B1(n8025), .B2(n6669), .Y(n8022) );
	o21ai_0 U8179( .A1(n6225), .A2(n7333), .B1(n8026), .Y(n5455) );
	mux2i_1 U8180( .A0(n8027), .A1(n6253), .S(n8028), .Y(n8026) );
	nor2_1 U8181( .A(n6898), .B(n7332), .Y(n8028) );
	nor2_1 U8182( .A(n6288), .B(n8029), .Y(n8027) );
	o22ai_1 U8183( .A1(n6208), .A2(n5920), .B1(n6277), .B2(n8030), .Y(n5454) );
	mux2i_1 U8184( .A0(n8031), .A1(n10447), .S(n8032), .Y(n8030) );
	o21ai_0 U8185( .A1(n6244), .A2(n8033), .B1(n8034), .Y(n5453) );
	mux2_1 U8186( .A0(n8035), .A1(n8036), .S(n11884), .X(n8034) );
	o21ai_0 U8187( .A1(n6241), .A2(n8037), .B1(n8038), .Y(n5452) );
	mux2i_1 U8188( .A0(n8039), .A1(n8040), .S(n8041), .Y(n8038) );
	nor2_1 U8189( .A(n10565), .B(n6363), .Y(n8040) );
	nor2_1 U8190( .A(n7544), .B(n8042), .Y(n8039) );
	o21ai_0 U8191( .A1(n6241), .A2(n8043), .B1(n8044), .Y(n5451) );
	mux2i_1 U8192( .A0(n8045), .A1(n8046), .S(n8047), .Y(n8044) );
	nor2_1 U8193( .A(n10402), .B(n6363), .Y(n8046) );
	nor2_1 U8194( .A(n7231), .B(n8048), .Y(n8045) );
	inv_1 U8195( .A(n10402), .Y(n7231) );
	o21ai_0 U8196( .A1(n6241), .A2(n8049), .B1(n8050), .Y(n5450) );
	mux2i_1 U8197( .A0(n8051), .A1(n8052), .S(n8053), .Y(n8050) );
	nor2_1 U8198( .A(n8054), .B(n8055), .Y(n8052) );
	inv_1 U8199( .A(n8056), .Y(n8055) );
	o211ai_1 U8200( .A1(n6203), .A2(n5882), .B1(n6400), .C1(n8057), .Y(n5449) );
	mux2i_1 U8201( .A0(n8058), .A1(n8059), .S(n8060), .Y(n8057) );
	nor2_1 U8202( .A(n6361), .B(n8061), .Y(n8059) );
	nor2_1 U8203( .A(n8062), .B(n6300), .Y(n8058) );
	o21ai_0 U8204( .A1(n6241), .A2(n5993), .B1(n8063), .Y(n5448) );
	mux2i_1 U8205( .A0(n8064), .A1(n6253), .S(n8065), .Y(n8063) );
	nor2_1 U8206( .A(n6491), .B(n6868), .Y(n8065) );
	nor2_1 U8207( .A(n6288), .B(n5972), .Y(n8064) );
	o21ai_0 U8208( .A1(n6241), .A2(n5978), .B1(n8066), .Y(n5447) );
	mux2i_1 U8209( .A0(n8067), .A1(n6253), .S(n8068), .Y(n8066) );
	nor2_1 U8210( .A(n8069), .B(n7611), .Y(n8068) );
	nor2_1 U8211( .A(n6288), .B(n5986), .Y(n8067) );
	nor2_1 U8212( .A(n6288), .B(n8070), .Y(n5446) );
	o21ai_0 U8213( .A1(n6241), .A2(n5923), .B1(n8071), .Y(n5445) );
	mux2i_1 U8214( .A0(n8072), .A1(n6253), .S(n8073), .Y(n8071) );
	nor2_1 U8215( .A(n6808), .B(n8074), .Y(n8073) );
	nor2_1 U8216( .A(n6289), .B(n8075), .Y(n8072) );
	o21ai_0 U8217( .A1(n6241), .A2(n6918), .B1(n8076), .Y(n5444) );
	a22oi_1 U8218( .A1(n7136), .A2(n8077), .B1(n10846), .B2(n7138), .Y(n8076) );
	inv_1 U8219( .A(n10847), .Y(n6918) );
	o21ai_0 U8220( .A1(n6241), .A2(n8078), .B1(n8079), .Y(n5443) );
	mux2i_1 U8221( .A0(n8080), .A1(n6253), .S(n8081), .Y(n8079) );
	nor2_1 U8222( .A(n7496), .B(n8082), .Y(n8081) );
	nor2_1 U8223( .A(n6289), .B(n8083), .Y(n8080) );
	o221ai_1 U8224( .A1(n8084), .A2(n8085), .B1(n6219), .B2(n7883), .C1(n8086), .Y(n5442) );
	o21ai_0 U8225( .A1(n8087), .A2(n6746), .B1(n11864), .Y(n8086) );
	a21oi_1 U8226( .A1(n8088), .A2(n8089), .B1(n6309), .Y(n8087) );
	a21oi_1 U8227( .A1(n8090), .A2(n7113), .B1(n8091), .Y(n8084) );
	nor4_1 U8228( .A(n10250), .B(n7039), .C(n8092), .D(n7111), .Y(n8091) );
	a21oi_1 U8229( .A1(n10260), .A2(n7089), .B1(n6308), .Y(n8090) );
	o22ai_1 U8230( .A1(n6314), .A2(n8093), .B1(n6196), .B2(n8094), .Y(n5441) );
	o21ai_0 U8231( .A1(n6241), .A2(n8095), .B1(n8096), .Y(n5440) );
	mux2i_1 U8232( .A0(n8097), .A1(n6253), .S(n8098), .Y(n8096) );
	nor2_1 U8233( .A(n7903), .B(n8099), .Y(n8098) );
	nor2_1 U8234( .A(n6289), .B(n7709), .Y(n8097) );
	o32ai_1 U8235( .A1(n8100), .A2(n8101), .A3(n8102), .B1(n6199), .B2(n8103), .Y(n5439) );
	inv_1 U8236( .A(n7094), .Y(n8102) );
	o21ai_0 U8237( .A1(n8104), .A2(n11807), .B1(n6343), .Y(n8100) );
	and3_1 U8238( .A(n6911), .B(n7096), .C(g7916), .X(n8104) );
	nor2_1 U8239( .A(n6784), .B(n8105), .Y(n5438) );
	nand3_1 U8240( .A(n8106), .B(n8107), .C(n6331), .Y(n6784) );
	o21ai_0 U8241( .A1(n6241), .A2(n6048), .B1(n8108), .Y(n5437) );
	mux2i_1 U8242( .A0(n8109), .A1(n8110), .S(n10318), .Y(n8108) );
	nor2_1 U8243( .A(n6289), .B(n7651), .Y(n8109) );
	inv_1 U8244( .A(n7653), .Y(n7651) );
	o22ai_1 U8245( .A1(n6207), .A2(n8111), .B1(n8112), .B2(n6296), .Y(n5436) );
	nor2_1 U8246( .A(n10938), .B(n8113), .Y(n8112) );
	o221ai_1 U8247( .A1(n8114), .A2(n8115), .B1(n6219), .B2(n8116), .C1(n8117), .Y(n5435) );
	nand3_1 U8248( .A(n6339), .B(n8118), .C(n10673), .Y(n8117) );
	o21ai_0 U8249( .A1(n6917), .A2(n8116), .B1(n6919), .Y(n8115) );
	inv_1 U8250( .A(n10736), .Y(n8116) );
	o21ai_0 U8251( .A1(n6241), .A2(n6029), .B1(n8119), .Y(n5434) );
	mux2i_1 U8252( .A0(n8120), .A1(n7345), .S(n8121), .Y(n8119) );
	nor2_1 U8253( .A(n7030), .B(n8019), .Y(n8121) );
	inv_1 U8254( .A(n7428), .Y(n8019) );
	nor2_1 U8255( .A(n10249), .B(n7347), .Y(n7428) );
	nor2_1 U8256( .A(n6289), .B(n5996), .Y(n8120) );
	nor2_1 U8257( .A(n5959), .B(n6300), .Y(n5433) );
	o221ai_1 U8258( .A1(n8122), .A2(n5943), .B1(n6218), .B2(n8123), .C1(n8124), .Y(n5432) );
	nand3_1 U8259( .A(n8125), .B(n8126), .C(n8127), .Y(n8124) );
	xnor2_1 U8260( .A(n8128), .B(n10676), .Y(n8126) );
	a21oi_1 U8261( .A1(n6331), .A2(n8129), .B1(n6747), .Y(n8122) );
	o32ai_1 U8262( .A1(n8130), .A2(n6349), .A3(n6509), .B1(n6510), .B2(n6697), .Y(n5431) );
	inv_1 U8263( .A(n10313), .Y(n6697) );
	nand2_1 U8264( .A(n6509), .B(n6380), .Y(n6510) );
	nor2_1 U8265( .A(n10271), .B(n8131), .Y(n5430) );
	o21ai_0 U8266( .A1(n6241), .A2(n6023), .B1(n8132), .Y(n5429) );
	mux2i_1 U8267( .A0(n8133), .A1(n6520), .S(n8134), .Y(n8132) );
	nor2_1 U8268( .A(n10262), .B(n7916), .Y(n8134) );
	nor2_1 U8269( .A(n6289), .B(n5981), .Y(n8133) );
	o21ai_0 U8270( .A1(n6241), .A2(n8135), .B1(n8136), .Y(n5428) );
	mux2i_1 U8271( .A0(n8137), .A1(n6254), .S(n8138), .Y(n8136) );
	nor2_1 U8272( .A(n6870), .B(n8139), .Y(n8138) );
	nor2_1 U8273( .A(n6290), .B(n8140), .Y(n8137) );
	o211ai_1 U8274( .A1(n8141), .A2(n8142), .B1(n8143), .C1(n8144), .Y(n5427) );
	nand3_1 U8275( .A(n11810), .B(n8145), .C(n8146), .Y(n8143) );
	a21oi_1 U8276( .A1(n8147), .A2(n8148), .B1(n6437), .Y(n8141) );
	o32ai_1 U8277( .A1(n6310), .A2(n8149), .A3(n8150), .B1(n6199), .B2(n8151), .Y(n5426) );
	a21oi_1 U8278( .A1(n6551), .A2(n7766), .B1(n10912), .Y(n8150) );
	nor3_1 U8279( .A(n10431), .B(n11828), .C(n6554), .Y(n6551) );
	nor3_1 U8280( .A(n8152), .B(n6409), .C(n6554), .Y(n8149) );
	xnor2_1 U8281( .A(n10283), .B(n6555), .Y(n8152) );
	nand2_1 U8282( .A(n8153), .B(n19679), .Y(n6555) );
	o21ai_0 U8283( .A1(n6241), .A2(n8154), .B1(n8155), .Y(n5425) );
	mux2i_1 U8284( .A0(n8156), .A1(n6254), .S(n8157), .Y(n8155) );
	nor2_1 U8285( .A(n7229), .B(n7731), .Y(n8157) );
	nor2_1 U8286( .A(n6291), .B(n7607), .Y(n8156) );
	nor3_1 U8287( .A(n8158), .B(n6350), .C(n8159), .Y(n5424) );
	a21oi_1 U8288( .A1(n10852), .A2(n8160), .B1(n7257), .Y(n8159) );
	nor3_1 U8289( .A(n8161), .B(n6427), .C(n7259), .Y(n8158) );
	o21ai_0 U8290( .A1(n6241), .A2(n8162), .B1(n8163), .Y(n5423) );
	mux2i_1 U8291( .A0(n8164), .A1(n6254), .S(n8165), .Y(n8163) );
	nor2_1 U8292( .A(n7875), .B(n7485), .Y(n8165) );
	nor2_1 U8293( .A(n6293), .B(n5973), .Y(n8164) );
	o22ai_1 U8294( .A1(n6205), .A2(n8166), .B1(n8167), .B2(n8168), .Y(n5422) );
	a222oi_1 U8295( .A1(n4714), .A2(n8169), .B1(n8170), .B2(n6382), .C1(n8171), .C2(n6341), .Y(n8168) );
	o22ai_1 U8296( .A1(n7241), .A2(n7239), .B1(n8172), .B2(n8173), .Y(n5421) );
	a21oi_1 U8297( .A1(n7242), .A2(n7241), .B1(n6437), .Y(n8172) );
	inv_1 U8298( .A(n8174), .Y(n7242) );
	o21ai_0 U8299( .A1(n6241), .A2(n8175), .B1(n8176), .Y(n5420) );
	mux2i_1 U8300( .A0(n8177), .A1(n8178), .S(n8179), .Y(n8176) );
	nor2_1 U8301( .A(n10409), .B(n6364), .Y(n8178) );
	nor2_1 U8302( .A(n7544), .B(n7538), .Y(n8177) );
	inv_1 U8303( .A(n10409), .Y(n7538) );
	o32ai_1 U8304( .A1(n8180), .A2(n6349), .A3(n8181), .B1(n7308), .B2(n7312), .Y(n5419) );
	inv_1 U8305( .A(n10628), .Y(n7312) );
	o22ai_1 U8306( .A1(n6302), .A2(n8182), .B1(n6196), .B2(n5880), .Y(n5418) );
	mux2i_1 U8307( .A0(n8183), .A1(n8184), .S(n8185), .Y(n5417) );
	or2_0 U8308( .A(n8025), .B(n8186), .X(n8184) );
	a21oi_1 U8309( .A1(n8187), .A2(n8186), .B1(n6437), .Y(n8183) );
	o21ai_0 U8310( .A1(n6241), .A2(n6008), .B1(n8188), .Y(n5416) );
	mux2i_1 U8311( .A0(n8189), .A1(n6254), .S(n8190), .Y(n8188) );
	nor2_1 U8312( .A(n6858), .B(n8191), .Y(n8190) );
	nor2_1 U8313( .A(n6282), .B(n5974), .Y(n8189) );
	o32ai_1 U8314( .A1(n8192), .A2(n6349), .A3(n7757), .B1(n7758), .B2(n8193), .Y(n5415) );
	inv_1 U8315( .A(n10693), .Y(n8192) );
	o22ai_1 U8316( .A1(n6204), .A2(n8194), .B1(n8195), .B2(n7863), .Y(n5414) );
	xnor2_1 U8317( .A(n8196), .B(n10357), .Y(n8195) );
	o21ai_0 U8318( .A1(n6242), .A2(n7508), .B1(n8197), .Y(n5413) );
	mux2i_1 U8319( .A0(n8198), .A1(n8199), .S(n8200), .Y(n8197) );
	nor2_1 U8320( .A(n6362), .B(n8201), .Y(n8199) );
	and2_0 U8321( .A(n8201), .B(n7513), .X(n8198) );
	inv_1 U8322( .A(n10571), .Y(n7508) );
	o21ai_0 U8323( .A1(n6242), .A2(n7043), .B1(n8202), .Y(n5412) );
	a22oi_1 U8324( .A1(n8203), .A2(n6529), .B1(n11938), .B2(n6534), .Y(n8202) );
	nand3_1 U8325( .A(n10340), .B(n7043), .C(n7862), .Y(n6529) );
	o22ai_1 U8326( .A1(n6204), .A2(n8204), .B1(n8205), .B2(n6294), .Y(n5411) );
	nor3_1 U8327( .A(n8113), .B(n10438), .C(n6822), .Y(n8205) );
	o221ai_1 U8328( .A1(n7208), .A2(n8206), .B1(n6219), .B2(n8207), .C1(n8208), .Y(n5410) );
	inv_1 U8329( .A(n10502), .Y(n8207) );
	inv_1 U8330( .A(n10640), .Y(n8206) );
	o21ai_0 U8331( .A1(n6242), .A2(n8209), .B1(n8210), .Y(n5409) );
	mux2i_1 U8332( .A0(n8211), .A1(n8212), .S(n8213), .Y(n8210) );
	nor2_1 U8333( .A(n10400), .B(n6364), .Y(n8212) );
	nor2_1 U8334( .A(n8043), .B(n8048), .Y(n8211) );
	o21ai_0 U8335( .A1(n6242), .A2(n7698), .B1(n8214), .Y(n5408) );
	mux2i_1 U8336( .A0(n8215), .A1(n6254), .S(n8216), .Y(n8214) );
	nor2_1 U8337( .A(n6888), .B(n8023), .Y(n8216) );
	nor2_1 U8338( .A(n6279), .B(n5994), .Y(n8215) );
	inv_1 U8339( .A(n10780), .Y(n7698) );
	o22ai_1 U8340( .A1(n8217), .A2(n8218), .B1(n8219), .B2(n8220), .Y(n5407) );
	a21oi_1 U8341( .A1(n8221), .A2(n8217), .B1(n6437), .Y(n8219) );
	o221ai_1 U8342( .A1(n8222), .A2(n8223), .B1(n6302), .B2(n8224), .C1(n6400), .Y(n5406) );
	a21oi_1 U8343( .A1(n6378), .A2(n8225), .B1(n6437), .Y(n8222) );
	o221ai_1 U8344( .A1(n8226), .A2(n7239), .B1(n6219), .B2(n7238), .C1(n8227), .Y(n5405) );
	a21oi_1 U8345( .A1(n8228), .A2(n8229), .B1(n8230), .Y(n8227) );
	nor3_1 U8346( .A(n8174), .B(n8231), .C(n7241), .Y(n8230) );
	nor2_1 U8347( .A(n7824), .B(n6300), .Y(n8228) );
	o221ai_1 U8348( .A1(n6212), .A2(n6068), .B1(n10182), .B2(n6312), .C1(n8232), .Y(n5404) );
	o21ai_0 U8349( .A1(n6242), .A2(n6024), .B1(n8233), .Y(n5403) );
	mux2i_1 U8350( .A0(n8234), .A1(n6559), .S(n8235), .Y(n8233) );
	nor2_1 U8351( .A(n10247), .B(n7562), .Y(n8235) );
	inv_1 U8352( .A(n8236), .Y(n7562) );
	nor2_1 U8353( .A(n6284), .B(n5995), .Y(n8234) );
	o221ai_1 U8354( .A1(n8237), .A2(n5890), .B1(n6764), .B2(n8238), .C1(n8239), .Y(n5402) );
	inv_1 U8355( .A(n8240), .Y(n6764) );
	a21oi_1 U8356( .A1(n6771), .A2(n6374), .B1(n6437), .Y(n8237) );
	o21ai_0 U8357( .A1(n6242), .A2(n5868), .B1(n8241), .Y(n5401) );
	mux2_1 U8358( .A0(n6844), .A1(n7168), .S(n10694), .X(n8241) );
	nand2_1 U8359( .A(n8242), .B(n6333), .Y(n6844) );
	o21ai_0 U8360( .A1(n6242), .A2(n5996), .B1(n8243), .Y(n5400) );
	mux2i_1 U8361( .A0(n8244), .A1(n7345), .S(n8245), .Y(n8243) );
	nor2_1 U8362( .A(n10259), .B(n7845), .Y(n8245) );
	nor2_1 U8363( .A(n6284), .B(n5975), .Y(n8244) );
	o221ai_1 U8364( .A1(n7038), .A2(n7427), .B1(n6217), .B2(n7040), .C1(n8246), .Y(n5399) );
	or3_1 U8365( .A(n7036), .B(n6369), .C(n7845), .X(n8246) );
	nand2_1 U8366( .A(n10249), .B(n7522), .Y(n7845) );
	o21ai_0 U8367( .A1(n6242), .A2(n5938), .B1(n8247), .Y(n5398) );
	mux2i_1 U8368( .A0(n8248), .A1(n6254), .S(n8249), .Y(n8247) );
	nor2_1 U8369( .A(n8250), .B(n8251), .Y(n8249) );
	nor2_1 U8370( .A(n6280), .B(n7707), .Y(n8248) );
	o22ai_1 U8371( .A1(n8252), .A2(n8253), .B1(n8254), .B2(n6297), .Y(n5397) );
	a21oi_1 U8372( .A1(n11842), .A2(n5962), .B1(n8255), .Y(n8254) );
	a211oi_1 U8373( .A1(n11842), .A2(n7514), .B1(n10918), .C1(n10543), .Y(n8255) );
	inv_1 U8374( .A(n10918), .Y(n8253) );
	nor2_1 U8375( .A(n8256), .B(n6437), .Y(n8252) );
	o221ai_1 U8376( .A1(n7075), .A2(n7374), .B1(n6219), .B2(n7644), .C1(n7376), .Y(n5396) );
	nand3_1 U8377( .A(n7375), .B(n6375), .C(n10324), .Y(n7376) );
	inv_1 U8378( .A(n10324), .Y(n7644) );
	inv_1 U8379( .A(n10637), .Y(n7374) );
	or2_0 U8380( .A(n6312), .B(n7375), .X(n7075) );
	nor3_1 U8381( .A(n6588), .B(n7954), .C(n5889), .Y(n7375) );
	o22ai_1 U8382( .A1(n6294), .A2(n7315), .B1(n6196), .B2(n7798), .Y(n5395) );
	inv_1 U8383( .A(n10702), .Y(n7798) );
	inv_1 U8384( .A(n10476), .Y(n7315) );
	o32ai_1 U8385( .A1(n8257), .A2(n6349), .A3(n6934), .B1(n6202), .B2(n8053), .Y(n5394) );
	mux2i_1 U8386( .A0(n8258), .A1(n10191), .S(n8259), .Y(n8257) );
	a21oi_1 U8387( .A1(n8260), .A2(n8261), .B1(n8054), .Y(n8258) );
	and2_0 U8388( .A(n8262), .B(n7050), .X(n8054) );
	o21ai_0 U8389( .A1(n6242), .A2(n5926), .B1(n8263), .Y(n5393) );
	mux2i_1 U8390( .A0(n8264), .A1(n6254), .S(n8265), .Y(n8263) );
	nor2_1 U8391( .A(n7026), .B(n8266), .Y(n8265) );
	nor2_1 U8392( .A(n6281), .B(n8267), .Y(n8264) );
	o22ai_1 U8393( .A1(n6206), .A2(n8268), .B1(n8269), .B2(n8048), .Y(n5392) );
	xnor2_1 U8394( .A(n8270), .B(n11858), .Y(n8269) );
	o21ai_0 U8395( .A1(n6242), .A2(n5879), .B1(n8271), .Y(n5391) );
	mux2i_1 U8396( .A0(n8272), .A1(n6425), .S(n10684), .Y(n8271) );
	inv_1 U8397( .A(n8273), .Y(n6425) );
	nor2_1 U8398( .A(n6283), .B(n8274), .Y(n8272) );
	o21ai_0 U8399( .A1(n6242), .A2(n7593), .B1(n8275), .Y(n5390) );
	mux2i_1 U8400( .A0(n8276), .A1(n8277), .S(n8278), .Y(n8275) );
	nor2_1 U8401( .A(n10401), .B(n6364), .Y(n8277) );
	nor2_1 U8402( .A(n7108), .B(n7993), .Y(n8276) );
	o21ai_0 U8403( .A1(n6242), .A2(n6535), .B1(n8279), .Y(n5389) );
	mux2i_1 U8404( .A0(n8280), .A1(n8281), .S(n8282), .Y(n8279) );
	nor2_1 U8405( .A(n7861), .B(n8283), .Y(n8281) );
	o21ai_0 U8406( .A1(n6313), .A2(n8284), .B1(n6810), .Y(n8280) );
	o22ai_1 U8407( .A1(n7051), .A2(n5905), .B1(n8285), .B2(n8286), .Y(n8284) );
	o22ai_1 U8408( .A1(n6207), .A2(n8286), .B1(n8287), .B2(n8288), .Y(n5388) );
	mux2i_1 U8409( .A0(n8289), .A1(n7746), .S(n8290), .Y(n8288) );
	o21ai_0 U8410( .A1(n6242), .A2(n5976), .B1(n8291), .Y(n5387) );
	mux2i_1 U8411( .A0(n8292), .A1(n6254), .S(n8293), .Y(n8291) );
	nor2_1 U8412( .A(n6680), .B(n7386), .Y(n8293) );
	nor2_1 U8413( .A(n6284), .B(n5977), .Y(n8292) );
	o21ai_0 U8414( .A1(n6242), .A2(n8294), .B1(n8295), .Y(n5386) );
	mux2i_1 U8415( .A0(n8296), .A1(n8297), .S(n8298), .Y(n8295) );
	nor2_1 U8416( .A(n8299), .B(n8300), .Y(n8296) );
	o32ai_1 U8417( .A1(n6072), .A2(n6349), .A3(n8301), .B1(n8194), .B2(n8302), .Y(n5385) );
	o22ai_1 U8418( .A1(n6208), .A2(n8303), .B1(n6347), .B2(n8304), .Y(n5384) );
	o21ai_0 U8419( .A1(n6242), .A2(n5983), .B1(n8305), .Y(n5383) );
	mux2i_1 U8420( .A0(n8306), .A1(n7303), .S(n8307), .Y(n8305) );
	nor2_1 U8421( .A(n7742), .B(n7602), .Y(n8307) );
	inv_1 U8422( .A(g25259), .Y(n7602) );
	nor2_1 U8423( .A(n6292), .B(n8308), .Y(n8306) );
	o21ai_0 U8424( .A1(n6242), .A2(n8309), .B1(n8310), .Y(n5382) );
	mux2i_1 U8425( .A0(n8311), .A1(n8312), .S(n8313), .Y(n8310) );
	nor2_1 U8426( .A(n10531), .B(n6364), .Y(n8312) );
	nor2_1 U8427( .A(n7103), .B(n7108), .Y(n8311) );
	inv_1 U8428( .A(n10531), .Y(n7103) );
	o32ai_1 U8429( .A1(n6310), .A2(n8314), .A3(n8315), .B1(n6202), .B2(n6853), .Y(n5381) );
	a21oi_1 U8430( .A1(n6850), .A2(n7102), .B1(n10583), .Y(n8315) );
	inv_1 U8431( .A(n7578), .Y(n7102) );
	nor4_1 U8432( .A(n10241), .B(n7578), .C(n8316), .D(n7914), .Y(n8314) );
	o221ai_1 U8433( .A1(n8317), .A2(n6308), .B1(n6218), .B2(n6647), .C1(n8232), .Y(n5380) );
	xnor2_1 U8434( .A(n10328), .B(n8318), .Y(n8317) );
	o21ai_0 U8435( .A1(n6242), .A2(n8319), .B1(n8320), .Y(n5379) );
	mux2i_1 U8436( .A0(n8321), .A1(n8322), .S(n8323), .Y(n8320) );
	nor2_1 U8437( .A(n6362), .B(n8324), .Y(n8322) );
	and2_0 U8438( .A(n8324), .B(n7083), .X(n8321) );
	inv_1 U8439( .A(n8325), .Y(n5378) );
	a22oi_1 U8440( .A1(n6437), .A2(n11964), .B1(n8326), .B2(n6337), .Y(n8325) );
	o221ai_1 U8441( .A1(n8327), .A2(n5968), .B1(n6218), .B2(n8328), .C1(n8329), .Y(n5377) );
	nand3_1 U8442( .A(n6340), .B(n8330), .C(n8331), .Y(n8329) );
	o22ai_1 U8443( .A1(n6301), .A2(n8332), .B1(n6195), .B2(n8333), .Y(n5376) );
	o21ai_0 U8444( .A1(n6243), .A2(n8334), .B1(n8335), .Y(n5375) );
	mux2i_1 U8445( .A0(n8336), .A1(n6254), .S(n8337), .Y(n8335) );
	nor2_1 U8446( .A(n8069), .B(n7731), .Y(n8337) );
	nor2_1 U8447( .A(n6289), .B(n5978), .Y(n8336) );
	o22ai_1 U8448( .A1(n6208), .A2(n5949), .B1(n8338), .B2(n6295), .Y(n5374) );
	nor2_1 U8449( .A(n8339), .B(n8340), .Y(n8338) );
	xnor2_1 U8450( .A(n10245), .B(n8341), .Y(n8340) );
	inv_1 U8451( .A(n8342), .Y(n8339) );
	o22ai_1 U8452( .A1(n6208), .A2(n8343), .B1(n8344), .B2(n6295), .Y(n5373) );
	nor3_1 U8453( .A(n7317), .B(n11859), .C(n10437), .Y(n8344) );
	inv_1 U8454( .A(g44), .Y(n7317) );
	o221ai_1 U8455( .A1(n8345), .A2(n8218), .B1(n6217), .B2(n8217), .C1(n8346), .Y(n5372) );
	a21oi_1 U8456( .A1(n8347), .A2(n8348), .B1(n8349), .Y(n8346) );
	nor3_1 U8457( .A(n8350), .B(n8220), .C(n8351), .Y(n8349) );
	and2_0 U8458( .A(n8352), .B(n6344), .X(n8347) );
	o21ai_0 U8459( .A1(n6243), .A2(n8353), .B1(n8354), .Y(n5371) );
	mux2i_1 U8460( .A0(n8355), .A1(n8356), .S(n8173), .Y(n8354) );
	nor2_1 U8461( .A(n10289), .B(n8174), .Y(n8356) );
	nand3_1 U8462( .A(n8107), .B(n6375), .C(n8357), .Y(n8174) );
	nor2_1 U8463( .A(n8357), .B(n7239), .Y(n8355) );
	o21ai_0 U8464( .A1(n6243), .A2(n8358), .B1(n8359), .Y(n5370) );
	mux2i_1 U8465( .A0(n6701), .A1(n8360), .S(n8361), .Y(n8359) );
	nor2_1 U8466( .A(n8362), .B(n8363), .Y(n8360) );
	inv_1 U8467( .A(n6700), .Y(n8363) );
	o221ai_1 U8468( .A1(n8364), .A2(n6309), .B1(n6217), .B2(n8365), .C1(n6400), .Y(n5369) );
	xnor2_1 U8469( .A(n10338), .B(n8366), .Y(n8364) );
	o21ai_0 U8470( .A1(n6243), .A2(n8367), .B1(n8368), .Y(n5368) );
	mux2i_1 U8471( .A0(n8369), .A1(n8370), .S(n8371), .Y(n8368) );
	nor2_1 U8472( .A(n10307), .B(n6364), .Y(n8370) );
	nor2_1 U8473( .A(n7108), .B(n8372), .Y(n8369) );
	o32ai_1 U8474( .A1(n8373), .A2(n10917), .A3(n6313), .B1(n6201), .B2(n6398), .Y(n5367) );
	and2_0 U8475( .A(n6384), .B(g8358), .X(n5366) );
	o21ai_0 U8476( .A1(n7758), .A2(n6049), .B1(n8374), .Y(n5365) );
	mux2i_1 U8477( .A0(n8375), .A1(n8376), .S(n8193), .Y(n8374) );
	inv_1 U8478( .A(n10626), .Y(n8193) );
	nor3_1 U8479( .A(n8377), .B(n10693), .C(n6306), .Y(n8376) );
	nand2_1 U8480( .A(n6221), .B(n8378), .Y(n8375) );
	nand3_1 U8481( .A(n7566), .B(n6378), .C(n10693), .Y(n8378) );
	a21oi_1 U8482( .A1(n6197), .A2(n8379), .B1(n5909), .Y(n5364) );
	or2_0 U8483( .A(n8380), .B(n6369), .X(n8379) );
	nor3_1 U8484( .A(n8381), .B(n6351), .C(n8382), .Y(n5363) );
	a21oi_1 U8485( .A1(n10856), .A2(n8383), .B1(n7257), .Y(n8382) );
	nor3_1 U8486( .A(n8384), .B(n7259), .C(n8385), .Y(n8381) );
	o32ai_1 U8487( .A1(n6297), .A2(g9741), .A3(n8386), .B1(n6202), .B2(n8387), .Y(n5362) );
	a21oi_1 U8488( .A1(g9682), .A2(n8387), .B1(n10607), .Y(n8386) );
	inv_1 U8489( .A(n10606), .Y(n8387) );
	o22ai_1 U8490( .A1(n7905), .A2(n8388), .B1(n7907), .B2(n8389), .Y(n5361) );
	o21ai_0 U8491( .A1(n8390), .A2(n10597), .B1(n6342), .Y(n8389) );
	a21oi_1 U8492( .A1(n8391), .A2(n8392), .B1(n8393), .Y(n8390) );
	mux2i_1 U8493( .A0(n8394), .A1(n8395), .S(n5910), .Y(n8392) );
	mux2i_1 U8494( .A0(n8396), .A1(n8397), .S(n8398), .Y(n8391) );
	inv_1 U8495( .A(n7908), .Y(n7907) );
	nor2_1 U8496( .A(n8399), .B(n8400), .Y(n7908) );
	inv_1 U8497( .A(n10597), .Y(n7905) );
	o21ai_0 U8498( .A1(n6243), .A2(n6049), .B1(n8401), .Y(n5360) );
	mux2i_1 U8499( .A0(n7565), .A1(n8402), .S(n8403), .Y(n8401) );
	nor2_1 U8500( .A(n6289), .B(n8377), .Y(n8402) );
	inv_1 U8501( .A(n7566), .Y(n8377) );
	inv_1 U8502( .A(n7758), .Y(n7565) );
	nand2_1 U8503( .A(n7757), .B(n6380), .Y(n7758) );
	nor2_1 U8504( .A(n6934), .B(n7566), .Y(n7757) );
	o21ai_0 U8505( .A1(n6243), .A2(n8404), .B1(n8405), .Y(n5359) );
	mux2i_1 U8506( .A0(n8406), .A1(n8407), .S(n8408), .Y(n8405) );
	nor2_1 U8507( .A(n8409), .B(n8410), .Y(n8407) );
	inv_1 U8508( .A(n8411), .Y(n8410) );
	o32ai_1 U8509( .A1(n8412), .A2(n6349), .A3(n8181), .B1(n7159), .B2(n7308), .Y(n5358) );
	nand2_1 U8510( .A(n8181), .B(n6380), .Y(n7308) );
	inv_1 U8511( .A(n10731), .Y(n7159) );
	nor2_1 U8512( .A(n6934), .B(n7313), .Y(n8181) );
	nor3_1 U8513( .A(n8413), .B(n6351), .C(n8414), .Y(n5357) );
	a21oi_1 U8514( .A1(n10853), .A2(n6509), .B1(n7257), .Y(n8414) );
	nor2_1 U8515( .A(n6934), .B(g26801), .Y(n6509) );
	nor3_1 U8516( .A(n8130), .B(n7259), .C(g26801), .Y(n8413) );
	inv_1 U8517( .A(n10853), .Y(n8130) );
	o21ai_0 U8518( .A1(n6517), .A2(n6098), .B1(n8415), .Y(n5356) );
	mux2i_1 U8519( .A0(n8416), .A1(n8417), .S(n8418), .Y(n8415) );
	nor2_1 U8520( .A(n10319), .B(n6516), .Y(n8417) );
	nand2_1 U8521( .A(n8419), .B(n6334), .Y(n6516) );
	nand2_1 U8522( .A(n6220), .B(n8420), .Y(n8416) );
	o21ai_0 U8523( .A1(n5933), .A2(n8421), .B1(n8422), .Y(n5355) );
	inv_1 U8524( .A(n8423), .Y(n8422) );
	o21ai_0 U8525( .A1(n6802), .A2(n8424), .B1(n6342), .Y(n8421) );
	o221ai_1 U8526( .A1(n8425), .A2(n6308), .B1(n6217), .B2(n8014), .C1(n8426), .Y(n5354) );
	nand4_1 U8527( .A(n10477), .B(n8427), .C(n8428), .D(n8429), .Y(n8426) );
	nor2_1 U8528( .A(n6362), .B(n8430), .Y(n8428) );
	a21oi_1 U8529( .A1(n10247), .A2(g35), .B1(n10265), .Y(n8430) );
	a21oi_1 U8530( .A1(n8431), .A2(n10477), .B1(n8432), .Y(n8425) );
	a21oi_1 U8531( .A1(n8429), .A2(n8427), .B1(n8433), .Y(n8432) );
	a21oi_1 U8532( .A1(n6561), .A2(n8434), .B1(n7653), .Y(n8433) );
	inv_1 U8533( .A(n8431), .Y(n6561) );
	or2_0 U8534( .A(n8435), .B(n10688), .X(n8427) );
	o221ai_1 U8535( .A1(n8436), .A2(n5877), .B1(n6217), .B2(n8437), .C1(n8438), .Y(n5353) );
	nand3_1 U8536( .A(n6757), .B(n8439), .C(n6759), .Y(n8438) );
	xnor2_1 U8537( .A(n8440), .B(n10675), .Y(n8439) );
	a21oi_1 U8538( .A1(n6331), .A2(n8441), .B1(n7836), .Y(n8436) );
	o21ai_0 U8539( .A1(n6243), .A2(n5979), .B1(n8442), .Y(n5352) );
	mux2i_1 U8540( .A0(n8443), .A1(n6254), .S(n8444), .Y(n8442) );
	nor2_1 U8541( .A(n6905), .B(n7611), .Y(n8444) );
	nor2_1 U8542( .A(n6289), .B(n5980), .Y(n8443) );
	o21ai_0 U8543( .A1(n7530), .A2(n6050), .B1(n8445), .Y(n5351) );
	mux2i_1 U8544( .A0(n8446), .A1(n8447), .S(n8448), .Y(n8445) );
	nor3_1 U8545( .A(n7645), .B(n10696), .C(n6306), .Y(n8447) );
	inv_1 U8546( .A(n7022), .Y(n7645) );
	nand2_1 U8547( .A(n6222), .B(n8449), .Y(n8446) );
	nand3_1 U8548( .A(n7022), .B(n6375), .C(n10696), .Y(n8449) );
	mux2i_1 U8549( .A0(n8450), .A1(n8451), .S(n10506), .Y(n5350) );
	a21oi_1 U8550( .A1(n6451), .A2(n6379), .B1(n6437), .Y(n8451) );
	xor2_1 U8551( .A(n8452), .B(n11896), .X(n6451) );
	nand2_1 U8552( .A(n8453), .B(n6333), .Y(n8450) );
	o21ai_0 U8553( .A1(n6243), .A2(n8454), .B1(n8455), .Y(n5349) );
	mux2i_1 U8554( .A0(n8456), .A1(n8457), .S(n8458), .Y(n8455) );
	nor2_1 U8555( .A(n10398), .B(n6364), .Y(n8457) );
	nor2_1 U8556( .A(n7108), .B(n8459), .Y(n8456) );
	o21ai_0 U8557( .A1(n6243), .A2(n8460), .B1(n8461), .Y(n5348) );
	a22oi_1 U8558( .A1(n7136), .A2(n7654), .B1(n10736), .B2(n7138), .Y(n8461) );
	inv_1 U8559( .A(n10583), .Y(n7654) );
	and2_0 U8560( .A(n6384), .B(g8279), .X(n5347) );
	o21ai_0 U8561( .A1(n6243), .A2(n5981), .B1(n8462), .Y(n5346) );
	mux2i_1 U8562( .A0(n8463), .A1(n6520), .S(n8464), .Y(n8462) );
	nor2_1 U8563( .A(n6522), .B(n6573), .Y(n8464) );
	inv_1 U8564( .A(n6456), .Y(n6522) );
	nor2_1 U8565( .A(n10252), .B(n6579), .Y(n6456) );
	nor2_1 U8566( .A(n6289), .B(n8465), .Y(n8463) );
	o22ai_1 U8567( .A1(n6303), .A2(n8182), .B1(n6195), .B2(n5951), .Y(n5345) );
	inv_1 U8568( .A(g6749), .Y(n8182) );
	o22ai_1 U8569( .A1(n8466), .A2(n8467), .B1(n8468), .B2(n8469), .Y(n5344) );
	a21oi_1 U8570( .A1(n8470), .A2(n8471), .B1(n6437), .Y(n8468) );
	and2_0 U8571( .A(n8472), .B(n7339), .X(n8470) );
	inv_1 U8572( .A(n8473), .Y(n7339) );
	inv_1 U8573( .A(n10719), .Y(n8466) );
	o21ai_0 U8574( .A1(n8123), .A2(n8474), .B1(n8475), .Y(n5343) );
	mux2i_1 U8575( .A0(n8476), .A1(n8477), .S(n10545), .Y(n8475) );
	nand2_1 U8576( .A(n6221), .B(n8478), .Y(n8477) );
	nand3_1 U8577( .A(n8479), .B(n6380), .C(n7088), .Y(n8478) );
	nor2_1 U8578( .A(n6289), .B(n8479), .Y(n8476) );
	nand2_1 U8579( .A(n10676), .B(n8129), .Y(n8479) );
	inv_1 U8580( .A(n8125), .Y(n8129) );
	inv_1 U8581( .A(n10676), .Y(n8123) );
	o21ai_0 U8582( .A1(n6243), .A2(n7253), .B1(n8480), .Y(n5342) );
	inv_1 U8583( .A(n8481), .Y(n8480) );
	o22ai_1 U8584( .A1(n8482), .A2(n6501), .B1(n8483), .B2(n8484), .Y(n8481) );
	o22ai_1 U8585( .A1(n6208), .A2(n8485), .B1(n10924), .B2(n8486), .Y(n5341) );
	mux2i_1 U8586( .A0(n8487), .A1(n8488), .S(n10406), .Y(n5340) );
	a21oi_1 U8587( .A1(n10671), .A2(n6373), .B1(n6437), .Y(n8488) );
	nand2_1 U8588( .A(n6338), .B(n8489), .Y(n8487) );
	and2_0 U8589( .A(n6385), .B(g8719), .X(n5339) );
	nor2_1 U8590( .A(n6361), .B(n8490), .Y(n5338) );
	o221ai_1 U8591( .A1(n8491), .A2(n6309), .B1(n6216), .B2(n7111), .C1(n8492), .Y(n5337) );
	nand4_1 U8592( .A(n10479), .B(n8493), .C(n8494), .D(n8495), .Y(n8492) );
	nor2_1 U8593( .A(n6362), .B(n8496), .Y(n8494) );
	a21oi_1 U8594( .A1(n10239), .A2(g35), .B1(n10260), .Y(n8496) );
	a21oi_1 U8595( .A1(n10479), .A2(n7884), .B1(n8497), .Y(n8491) );
	a21oi_1 U8596( .A1(n8495), .A2(n8493), .B1(n8498), .Y(n8497) );
	a21oi_1 U8597( .A1(n8499), .A2(n8500), .B1(n8501), .Y(n8498) );
	or2_0 U8598( .A(n8502), .B(n10688), .X(n8493) );
	o221ai_1 U8599( .A1(n8503), .A2(n6706), .B1(n6216), .B2(n5964), .C1(n8504), .Y(n5336) );
	a21oi_1 U8600( .A1(n7662), .A2(n10301), .B1(n7716), .Y(n8504) );
	inv_1 U8601( .A(n7661), .Y(n6706) );
	o221ai_1 U8602( .A1(n8505), .A2(n5896), .B1(n7832), .B2(n6753), .C1(n7828), .Y(n5335) );
	inv_1 U8603( .A(n6758), .Y(n7828) );
	a21oi_1 U8604( .A1(n8506), .A2(n6381), .B1(n6437), .Y(n8505) );
	nor2_1 U8605( .A(n6599), .B(n8507), .Y(n5334) );
	nor2_1 U8606( .A(n6362), .B(n8508), .Y(n5333) );
	nor2_1 U8607( .A(n6362), .B(n8509), .Y(n5332) );
	o21ai_0 U8608( .A1(n6243), .A2(n8510), .B1(n8511), .Y(n5331) );
	mux2i_1 U8609( .A0(n8512), .A1(n8513), .S(n8209), .Y(n8511) );
	nor2_1 U8610( .A(n6362), .B(n8514), .Y(n8513) );
	and2_0 U8611( .A(n8514), .B(n7237), .X(n8512) );
	o21ai_0 U8612( .A1(n6243), .A2(n7424), .B1(n8515), .Y(n5330) );
	mux2i_1 U8613( .A0(n8516), .A1(n8517), .S(n8518), .Y(n8515) );
	nor2_1 U8614( .A(n8519), .B(n8520), .Y(n8517) );
	nor2_1 U8615( .A(n6289), .B(n8521), .Y(n8516) );
	o22ai_1 U8616( .A1(n8522), .A2(n8523), .B1(n8524), .B2(n6530), .Y(n5329) );
	nor2_1 U8617( .A(n7416), .B(n8525), .Y(n8524) );
	a21oi_1 U8618( .A1(n6331), .A2(n8526), .B1(n6534), .Y(n8522) );
	nor2_1 U8619( .A(n10275), .B(n8527), .Y(n5328) );
	o22ai_1 U8620( .A1(n8528), .A2(n8529), .B1(n8530), .B2(n8531), .Y(n5327) );
	o21ai_0 U8621( .A1(n8532), .A2(n8259), .B1(n6342), .Y(n8531) );
	o21ai_0 U8622( .A1(n8533), .A2(n8534), .B1(n8056), .Y(n8529) );
	mux2i_1 U8623( .A0(n8260), .A1(n8535), .S(n5912), .Y(n8534) );
	mux2i_1 U8624( .A0(n8536), .A1(n8261), .S(n8049), .Y(n8533) );
	inv_1 U8625( .A(n10413), .Y(n8049) );
	o22ai_1 U8626( .A1(n6207), .A2(n8537), .B1(n8538), .B2(n6295), .Y(n5326) );
	and4_1 U8627( .A(n8539), .B(n8540), .C(n8541), .D(n8542), .X(n8538) );
	o21ai_0 U8628( .A1(n6243), .A2(n6005), .B1(n8543), .Y(n5325) );
	mux2i_1 U8629( .A0(n8544), .A1(n6254), .S(n8545), .Y(n8543) );
	nor2_1 U8630( .A(n7353), .B(n6971), .Y(n8545) );
	nor2_1 U8631( .A(n6289), .B(n6687), .Y(n8544) );
	inv_1 U8632( .A(n10493), .Y(n6687) );
	o21ai_0 U8633( .A1(n8033), .A2(n8036), .B1(n8546), .Y(n5324) );
	mux2i_1 U8634( .A0(n8547), .A1(n8548), .S(n8549), .Y(n8546) );
	nor2_1 U8635( .A(n10505), .B(n8035), .Y(n8548) );
	nand2_1 U8636( .A(n6220), .B(n8550), .Y(n8547) );
	o21ai_0 U8637( .A1(n7154), .A2(n8551), .B1(n8552), .Y(n5323) );
	mux2i_1 U8638( .A0(n8553), .A1(n8554), .S(n10345), .Y(n8552) );
	nand2_1 U8639( .A(n6222), .B(n8555), .Y(n8554) );
	nand3_1 U8640( .A(n8556), .B(n6375), .C(n7220), .Y(n8555) );
	nor2_1 U8641( .A(n6288), .B(n8556), .Y(n8553) );
	nand2_1 U8642( .A(n10679), .B(n7160), .Y(n8556) );
	inv_1 U8643( .A(n7156), .Y(n7160) );
	inv_1 U8644( .A(n10679), .Y(n7154) );
	o221ai_1 U8645( .A1(n7485), .A2(n8557), .B1(n6212), .B2(n8558), .C1(n8559), .Y(n5322) );
	or3_1 U8646( .A(n6314), .B(n8560), .C(n7386), .X(n8559) );
	o21ai_0 U8647( .A1(n6243), .A2(n8561), .B1(n8562), .Y(n5321) );
	mux2i_1 U8648( .A0(n8563), .A1(n8564), .S(n8565), .Y(n8562) );
	nor2_1 U8649( .A(n6363), .B(n8566), .Y(n8564) );
	and2_0 U8650( .A(n8566), .B(n6344), .X(n8563) );
	nand3_1 U8651( .A(n10909), .B(n8567), .C(n8568), .Y(n8566) );
	inv_1 U8652( .A(n10909), .Y(n8561) );
	o21ai_0 U8653( .A1(n6243), .A2(n8140), .B1(n8569), .Y(n5320) );
	mux2i_1 U8654( .A0(n8570), .A1(n6254), .S(n8571), .Y(n8569) );
	nor2_1 U8655( .A(n6868), .B(n8139), .Y(n8571) );
	nand2_1 U8656( .A(n11943), .B(n6865), .Y(n6868) );
	nor2_1 U8657( .A(n6288), .B(n5940), .Y(n8570) );
	inv_1 U8658( .A(n10800), .Y(n8140) );
	o221ai_1 U8659( .A1(n6034), .A2(n8572), .B1(n8573), .B2(n8574), .C1(n8575), .Y(n5319) );
	a22oi_1 U8660( .A1(n7161), .A2(n10345), .B1(n10336), .B2(n6437), .Y(n8575) );
	inv_1 U8661( .A(n7158), .Y(n8574) );
	a221oi_1 U8662( .A1(n10724), .A2(n7219), .B1(n7156), .B2(n11804), .C1(n8576), .Y(n8573) );
	o32ai_1 U8663( .A1(n7218), .A2(n11915), .A3(n10336), .B1(n10175), .B2(n8577), .Y(n8576) );
	a22oi_1 U8664( .A1(n10336), .A2(n11778), .B1(n11805), .B2(n11915), .Y(n8577) );
	o21ai_0 U8665( .A1(n6243), .A2(n7934), .B1(n8578), .Y(n5318) );
	a22oi_1 U8666( .A1(n10459), .A2(n7369), .B1(g14201), .B2(n7370), .Y(n8578) );
	o22ai_1 U8667( .A1(n6207), .A2(n8579), .B1(n8580), .B2(n6296), .Y(n5317) );
	nor2_1 U8668( .A(n10516), .B(n6531), .Y(n8580) );
	inv_1 U8669( .A(g20899), .Y(n6531) );
	inv_1 U8670( .A(n10233), .Y(n8579) );
	o32ai_1 U8671( .A1(n8581), .A2(n10261), .A3(n7432), .B1(n7121), .B2(n7429), .Y(n5316) );
	nand2_1 U8672( .A(n7433), .B(n6334), .Y(n7429) );
	o21ai_0 U8673( .A1(n10240), .A2(n7461), .B1(n6342), .Y(n8581) );
	nor2_1 U8674( .A(n10251), .B(n7433), .Y(n7461) );
	o21ai_0 U8675( .A1(n6244), .A2(n6051), .B1(n8582), .Y(n5315) );
	mux2i_1 U8676( .A0(n8583), .A1(n8584), .S(n8585), .Y(n8582) );
	nor2_1 U8677( .A(n6288), .B(n7523), .Y(n8584) );
	o22ai_1 U8678( .A1(n6303), .A2(n8586), .B1(n6195), .B2(n8587), .Y(n5314) );
	o22ai_1 U8679( .A1(n6303), .A2(n8588), .B1(n6195), .B2(n8332), .Y(n5313) );
	inv_1 U8680( .A(n8589), .Y(n5312) );
	a221oi_1 U8681( .A1(n7918), .A2(n7136), .B1(n7138), .B2(n10845), .C1(n8590), .Y(n8589) );
	and2_0 U8682( .A(g20654), .B(n6437), .X(n8590) );
	inv_1 U8683( .A(n10582), .Y(n7918) );
	and2_0 U8684( .A(g6745), .B(n6344), .X(n5311) );
	o221ai_1 U8685( .A1(n7221), .A2(n8591), .B1(n6213), .B2(n6075), .C1(n8592), .Y(n5310) );
	or4_1 U8686( .A(n7887), .B(n6314), .C(n7893), .D(n8593), .X(n8592) );
	o22ai_1 U8687( .A1(n6207), .A2(n8594), .B1(n8595), .B2(n6296), .Y(n5309) );
	nor2_1 U8688( .A(n10622), .B(n8596), .Y(n8595) );
	inv_1 U8689( .A(n10577), .Y(n8594) );
	o21ai_0 U8690( .A1(n6244), .A2(n6979), .B1(n8597), .Y(n5308) );
	mux2i_1 U8691( .A0(n8598), .A1(n8599), .S(n8600), .Y(n8597) );
	nor2_1 U8692( .A(n6288), .B(n6977), .Y(n8599) );
	o21ai_0 U8693( .A1(n6244), .A2(n6042), .B1(n8601), .Y(n5307) );
	mux2i_1 U8694( .A0(n6689), .A1(n8602), .S(n8603), .Y(n8601) );
	nor2_1 U8695( .A(n6288), .B(n8604), .Y(n8602) );
	inv_1 U8696( .A(n7396), .Y(n6689) );
	o22ai_1 U8697( .A1(n6206), .A2(n6975), .B1(n8600), .B2(n6296), .Y(n5306) );
	o21ai_0 U8698( .A1(n6244), .A2(n8459), .B1(n8605), .Y(n5305) );
	mux2i_1 U8699( .A0(n8606), .A1(n8607), .S(n8608), .Y(n8605) );
	nor2_1 U8700( .A(n10392), .B(n6364), .Y(n8607) );
	nor2_1 U8701( .A(n7108), .B(n8609), .Y(n8606) );
	inv_1 U8702( .A(n10398), .Y(n8459) );
	o21ai_0 U8703( .A1(n6244), .A2(n8610), .B1(n8611), .Y(n5304) );
	mux2i_1 U8704( .A0(n8612), .A1(n6254), .S(n8613), .Y(n8611) );
	nor2_1 U8705( .A(n8614), .B(n7178), .Y(n8613) );
	nor2_1 U8706( .A(n6288), .B(n8615), .Y(n8612) );
	o22ai_1 U8707( .A1(n6207), .A2(n8616), .B1(n8617), .B2(n6296), .Y(n5303) );
	nor2_1 U8708( .A(n11818), .B(n8618), .Y(n8617) );
	inv_1 U8709( .A(n10622), .Y(n8616) );
	nor2_1 U8710( .A(n6362), .B(n8619), .Y(n5302) );
	o22ai_1 U8711( .A1(n6840), .A2(n8620), .B1(n6837), .B2(n8621), .Y(n5301) );
	o21ai_0 U8712( .A1(n6842), .A2(n8622), .B1(n6342), .Y(n8621) );
	inv_1 U8713( .A(n10935), .Y(n6837) );
	o21ai_0 U8714( .A1(n8623), .A2(n8624), .B1(n6700), .Y(n8620) );
	mux2i_1 U8715( .A0(n8625), .A1(n8626), .S(n5911), .Y(n8624) );
	mux2i_1 U8716( .A0(n8627), .A1(n8628), .S(n8358), .Y(n8623) );
	inv_1 U8717( .A(n10417), .Y(n8358) );
	o22ai_1 U8718( .A1(n6206), .A2(n8225), .B1(n8629), .B2(n6396), .Y(n5300) );
	nand2_1 U8719( .A(n10714), .B(n6333), .Y(n6396) );
	xnor2_1 U8720( .A(n8630), .B(n10244), .Y(n8629) );
	mux2i_1 U8721( .A0(n8631), .A1(n8632), .S(n10924), .Y(n5299) );
	a21oi_1 U8722( .A1(n8633), .A2(n8634), .B1(n6437), .Y(n8632) );
	nor2_1 U8723( .A(n11819), .B(n6364), .Y(n8633) );
	or2_0 U8724( .A(n6053), .B(n8486), .X(n8631) );
	nor2_1 U8725( .A(n6361), .B(n8635), .Y(n5298) );
	o21ai_0 U8726( .A1(n5878), .A2(n8636), .B1(n8637), .Y(n5297) );
	mux2i_1 U8727( .A0(n8638), .A1(n8639), .S(n10901), .Y(n8637) );
	nand2_1 U8728( .A(n6221), .B(n8640), .Y(n8639) );
	nand3_1 U8729( .A(n6386), .B(n8641), .C(n8642), .Y(n8640) );
	nor2_1 U8730( .A(n8643), .B(n8641), .Y(n8638) );
	o32ai_1 U8731( .A1(n6296), .A2(n10326), .A3(n8644), .B1(n6202), .B2(n7581), .Y(n5296) );
	inv_1 U8732( .A(n10703), .Y(n7581) );
	xnor2_1 U8733( .A(n11861), .B(n7896), .Y(n8644) );
	and3_1 U8734( .A(g12923), .B(n7898), .C(n10703), .X(n7896) );
	o21ai_0 U8735( .A1(n6244), .A2(n8645), .B1(n8646), .Y(n5295) );
	mux2i_1 U8736( .A0(n8647), .A1(n6255), .S(n8648), .Y(n8646) );
	nor2_1 U8737( .A(n6482), .B(n7015), .Y(n8648) );
	nor2_1 U8738( .A(n6288), .B(n8649), .Y(n8647) );
	o22ai_1 U8739( .A1(n6206), .A2(n7775), .B1(n8650), .B2(n6296), .Y(n5294) );
	a22oi_1 U8740( .A1(n10406), .A2(n8651), .B1(n10219), .B2(n10671), .Y(n8650) );
	o21ai_0 U8741( .A1(n7381), .A2(n8652), .B1(n10219), .Y(n8651) );
	a211oi_1 U8742( .A1(n6816), .A2(n8653), .B1(n8654), .C1(n10340), .Y(n8652) );
	inv_1 U8743( .A(n8655), .Y(n7381) );
	o21ai_0 U8744( .A1(n6244), .A2(n8308), .B1(n8656), .Y(n5293) );
	mux2i_1 U8745( .A0(n8657), .A1(n7303), .S(n8658), .Y(n8656) );
	nor2_1 U8746( .A(n10268), .B(n8659), .Y(n8658) );
	nor2_1 U8747( .A(n6288), .B(n5997), .Y(n8657) );
	inv_1 U8748( .A(n10930), .Y(n8308) );
	nor2_1 U8749( .A(n10272), .B(n8660), .Y(n5292) );
	o22ai_1 U8750( .A1(n6206), .A2(n8661), .B1(n8662), .B2(n6296), .Y(n5291) );
	nor3_1 U8751( .A(n8618), .B(n10716), .C(n8596), .Y(n8662) );
	or2_0 U8752( .A(n8663), .B(n8664), .X(n8596) );
	inv_1 U8753( .A(g91), .Y(n8618) );
	o32ai_1 U8754( .A1(n6295), .A2(g9817), .A3(n8665), .B1(n6201), .B2(n8666), .Y(n5290) );
	a21oi_1 U8755( .A1(g9743), .A2(n8666), .B1(n10605), .Y(n8665) );
	inv_1 U8756( .A(n10604), .Y(n8666) );
	a21oi_1 U8757( .A1(n6197), .A2(n8667), .B1(n5913), .Y(n5289) );
	or2_0 U8758( .A(n8668), .B(n6369), .X(n8667) );
	o21ai_0 U8759( .A1(n6244), .A2(n7808), .B1(n8669), .Y(n5288) );
	mux2i_1 U8760( .A0(n8670), .A1(n6255), .S(n8671), .Y(n8669) );
	nor2_1 U8761( .A(n6898), .B(n7669), .Y(n8671) );
	nor2_1 U8762( .A(n6288), .B(n6002), .Y(n8670) );
	inv_1 U8763( .A(n10747), .Y(n7808) );
	o21ai_0 U8764( .A1(n6244), .A2(n7187), .B1(n8672), .Y(n5287) );
	a22oi_1 U8765( .A1(n6719), .A2(n10836), .B1(n8385), .B2(n6249), .Y(n8672) );
	inv_1 U8766( .A(n8673), .Y(n6719) );
	inv_1 U8767( .A(n10500), .Y(n7187) );
	o21ai_0 U8768( .A1(n6244), .A2(n5888), .B1(n8674), .Y(n5286) );
	mux2i_1 U8769( .A0(n8675), .A1(n8676), .S(n8677), .Y(n8674) );
	nor2_1 U8770( .A(n6363), .B(n8678), .Y(n8676) );
	nor2_1 U8771( .A(n8679), .B(n7108), .Y(n8675) );
	inv_1 U8772( .A(n8678), .Y(n8679) );
	o21ai_0 U8773( .A1(n6244), .A2(n8680), .B1(n8681), .Y(n5285) );
	a22oi_1 U8774( .A1(n8110), .A2(n11773), .B1(n7653), .B2(n6559), .Y(n8681) );
	inv_1 U8775( .A(n7646), .Y(n8110) );
	o21ai_0 U8776( .A1(n6753), .A2(n8437), .B1(n8682), .Y(n5284) );
	mux2i_1 U8777( .A0(n8683), .A1(n8684), .S(n10344), .Y(n8682) );
	nand2_1 U8778( .A(n6222), .B(n8685), .Y(n8684) );
	nand3_1 U8779( .A(n8686), .B(n6381), .C(n8506), .Y(n8685) );
	nor2_1 U8780( .A(n6287), .B(n8686), .Y(n8683) );
	nand2_1 U8781( .A(n10675), .B(n8441), .Y(n8686) );
	inv_1 U8782( .A(n6759), .Y(n8441) );
	nor2_1 U8783( .A(n7832), .B(n11901), .Y(n6759) );
	inv_1 U8784( .A(n10675), .Y(n8437) );
	o32ai_1 U8785( .A1(n6310), .A2(n10364), .A3(g4467), .B1(n6202), .B2(n7870), .Y(n5283) );
	inv_1 U8786( .A(n10297), .Y(n7870) );
	o221ai_1 U8787( .A1(n7731), .A2(n8687), .B1(n6214), .B2(n8688), .C1(n8689), .Y(n5282) );
	or3_1 U8788( .A(n6314), .B(n8690), .C(n7611), .X(n8689) );
	nor2_1 U8789( .A(n8691), .B(n6063), .Y(n5281) );
	a221oi_1 U8790( .A1(n8256), .A2(n7514), .B1(n8692), .B2(n6377), .C1(n6437), .Y(n8691) );
	nor2_1 U8791( .A(n11791), .B(n10543), .Y(n8692) );
	inv_1 U8792( .A(n10464), .Y(n7514) );
	o22ai_1 U8793( .A1(n6299), .A2(n8333), .B1(n6195), .B2(n8693), .Y(n5280) );
	o221ai_1 U8794( .A1(n6795), .A2(n8694), .B1(n6214), .B2(n8695), .C1(n8696), .Y(n5279) );
	nand3_1 U8795( .A(n8697), .B(n5933), .C(n8423), .Y(n8696) );
	nor3_1 U8796( .A(n6306), .B(n10430), .C(n6802), .Y(n8423) );
	o21ai_0 U8797( .A1(n6802), .A2(n8697), .B1(n6342), .Y(n8694) );
	xnor2_1 U8798( .A(n8698), .B(n10285), .Y(n8697) );
	inv_1 U8799( .A(n8699), .Y(n6802) );
	inv_1 U8800( .A(n10907), .Y(n6795) );
	nor2_1 U8801( .A(n6287), .B(n8700), .Y(n5278) );
	mux2i_1 U8802( .A0(n8701), .A1(n10870), .S(n8654), .Y(n8700) );
	nand4_1 U8803( .A(g8719), .B(n10537), .C(n10921), .D(n6523), .Y(n8654) );
	nand2_1 U8804( .A(n6816), .B(n8653), .Y(n8701) );
	nand3_1 U8805( .A(n6815), .B(n7043), .C(n8702), .Y(n8653) );
	mux2i_1 U8806( .A0(n8703), .A1(n8704), .S(n7743), .Y(n8702) );
	o211ai_1 U8807( .A1(n7769), .A2(n8705), .B1(n8706), .C1(n6811), .Y(n8704) );
	nand2_1 U8808( .A(n8707), .B(n8708), .Y(n8703) );
	xnor2_1 U8809( .A(n5919), .B(n10354), .Y(n8707) );
	xnor2_1 U8810( .A(n10168), .B(n8709), .Y(n6816) );
	a21oi_1 U8811( .A1(n10859), .A2(n8710), .B1(n8711), .Y(n8709) );
	mux2i_1 U8812( .A0(n8712), .A1(n8713), .S(n7770), .Y(n8711) );
	nand2_1 U8813( .A(n10442), .B(n7743), .Y(n8713) );
	nand2_1 U8814( .A(n10734), .B(n10339), .Y(n8712) );
	xnor2_1 U8815( .A(n7770), .B(n10339), .Y(n8710) );
	o21ai_0 U8816( .A1(n6244), .A2(n8714), .B1(n8715), .Y(n5277) );
	mux2i_1 U8817( .A0(n8716), .A1(n8717), .S(n8718), .Y(n8715) );
	nor3_1 U8818( .A(n8719), .B(n10719), .C(n8473), .Y(n8717) );
	nor2_1 U8819( .A(n8720), .B(n8467), .Y(n8716) );
	inv_1 U8820( .A(n8719), .Y(n8720) );
	o221ai_1 U8821( .A1(n8721), .A2(n8722), .B1(n8723), .B2(n6225), .C1(n8724), .Y(n5276) );
	a21oi_1 U8822( .A1(n8725), .A2(n8726), .B1(n8727), .Y(n8724) );
	a21oi_1 U8823( .A1(n7279), .A2(n6389), .B1(n6309), .Y(n8727) );
	inv_1 U8824( .A(n7275), .Y(n6389) );
	nor2_1 U8825( .A(g7946), .B(n6364), .Y(n8725) );
	inv_1 U8826( .A(n61), .Y(n8721) );
	o21ai_0 U8827( .A1(n6948), .A2(n6951), .B1(n8728), .Y(n5275) );
	mux2i_1 U8828( .A0(n8729), .A1(n8730), .S(n8731), .Y(n8728) );
	nor2_1 U8829( .A(n10683), .B(n6950), .Y(n8730) );
	nand2_1 U8830( .A(n7946), .B(n6333), .Y(n6950) );
	nand2_1 U8831( .A(n6221), .B(n8732), .Y(n8729) );
	inv_1 U8832( .A(n10865), .Y(n6948) );
	o22ai_1 U8833( .A1(g23612), .A2(n6203), .B1(n8733), .B2(n6296), .Y(n5274) );
	nor2_1 U8834( .A(n10234), .B(n10663), .Y(n8733) );
	o21ai_0 U8835( .A1(n8734), .A2(n8735), .B1(n8736), .Y(n5273) );
	nand4_1 U8836( .A(n6339), .B(n8737), .C(n8738), .D(n8014), .Y(n8736) );
	o21ai_0 U8837( .A1(n8431), .A2(n10287), .B1(n8734), .Y(n8737) );
	o21ai_0 U8838( .A1(n6244), .A2(n5887), .B1(n8739), .Y(n5272) );
	mux2i_1 U8839( .A0(n8740), .A1(n8741), .S(n7051), .Y(n8739) );
	inv_1 U8840( .A(n10427), .Y(n7051) );
	and2_0 U8841( .A(n7058), .B(n7057), .X(n8741) );
	nor2_1 U8842( .A(n7058), .B(n7056), .Y(n8740) );
	nor2_1 U8843( .A(n5887), .B(n8742), .Y(n7058) );
	a21oi_1 U8844( .A1(n6198), .A2(n8743), .B1(n5914), .Y(n5271) );
	nand2_1 U8845( .A(n8744), .B(n6380), .Y(n8743) );
	o21ai_0 U8846( .A1(n6244), .A2(n8745), .B1(n8746), .Y(n5270) );
	mux2i_1 U8847( .A0(n8747), .A1(n6255), .S(n8748), .Y(n8746) );
	nor2_1 U8848( .A(n7016), .B(n7965), .Y(n8748) );
	nor2_1 U8849( .A(n6287), .B(n8749), .Y(n8747) );
	o22ai_1 U8850( .A1(n6303), .A2(n7799), .B1(n6194), .B2(n5872), .Y(n5269) );
	o221ai_1 U8851( .A1(n5895), .A2(n8551), .B1(n6214), .B2(n8077), .C1(n8750), .Y(n5268) );
	a21oi_1 U8852( .A1(n8751), .A2(n7158), .B1(n8752), .Y(n8750) );
	nor2_1 U8853( .A(n10336), .B(n7156), .Y(n8751) );
	nor2_1 U8854( .A(n7722), .B(n11915), .Y(n7156) );
	inv_1 U8855( .A(n10584), .Y(n8077) );
	o32ai_1 U8856( .A1(n6622), .A2(n6349), .A3(n8753), .B1(n7646), .B2(n7650), .Y(n5267) );
	inv_1 U8857( .A(n10623), .Y(n7650) );
	inv_1 U8858( .A(n10690), .Y(n6622) );
	o21ai_0 U8859( .A1(n6244), .A2(n8754), .B1(n8755), .Y(n5266) );
	mux2i_1 U8860( .A0(n8756), .A1(n8757), .S(n8758), .Y(n8755) );
	nor2_1 U8861( .A(n10408), .B(n6365), .Y(n8757) );
	nor2_1 U8862( .A(n8486), .B(n8759), .Y(n8756) );
	nor2_1 U8863( .A(n8760), .B(n8761), .Y(n5265) );
	nor2_1 U8864( .A(n6361), .B(n6554), .Y(n5264) );
	o21ai_0 U8865( .A1(n6244), .A2(n8762), .B1(n8763), .Y(n5263) );
	a22oi_1 U8866( .A1(n11821), .A2(n6603), .B1(n6602), .B2(n6605), .Y(n8763) );
	nand2_1 U8867( .A(n8764), .B(n8765), .Y(n6605) );
	mux2i_1 U8868( .A0(n8766), .A1(n8767), .S(n8768), .Y(n8765) );
	xnor2_1 U8869( .A(n8769), .B(g11349), .Y(n8768) );
	nand3_1 U8870( .A(n8770), .B(n8771), .C(n8772), .Y(n8767) );
	nand3_1 U8871( .A(n8773), .B(g16603), .C(n10500), .Y(n8772) );
	nand3_1 U8872( .A(g13895), .B(n8774), .C(n11823), .Y(n8771) );
	nand3_1 U8873( .A(n8775), .B(g16718), .C(n11856), .Y(n8770) );
	nand3_1 U8874( .A(n8776), .B(n8777), .C(n8778), .Y(n8766) );
	nand3_1 U8875( .A(n6607), .B(n11899), .C(g16718), .Y(n8778) );
	nand3_1 U8876( .A(n8774), .B(n10842), .C(g16603), .Y(n8777) );
	nand3_1 U8877( .A(g13895), .B(n8773), .C(n11900), .Y(n8776) );
	mux2_1 U8878( .A0(n8779), .A1(n8780), .S(n8769), .X(n8764) );
	a221oi_1 U8879( .A1(n8773), .A2(n8781), .B1(n6607), .B2(n8782), .C1(n8783), .Y(n8780) );
	o32ai_1 U8880( .A1(n5937), .A2(n7201), .A3(n8784), .B1(n8785), .B2(n7199), .Y(n8783) );
	a22oi_1 U8881( .A1(n10834), .A2(g16624), .B1(n10835), .B2(g16686), .Y(n8785) );
	o22ai_1 U8882( .A1(n6503), .A2(n8786), .B1(n8787), .B2(n7191), .Y(n8782) );
	o22ai_1 U8883( .A1(n8788), .A2(n6675), .B1(n6497), .B2(n8789), .Y(n8781) );
	inv_1 U8884( .A(n10830), .Y(n6497) );
	inv_1 U8885( .A(n10831), .Y(n6675) );
	inv_1 U8886( .A(n7200), .Y(n8773) );
	a221oi_1 U8887( .A1(n8775), .A2(n8790), .B1(n6607), .B2(n8791), .C1(n8792), .Y(n8779) );
	o32ai_1 U8888( .A1(n5935), .A2(n7200), .A3(n8784), .B1(n8793), .B2(n7201), .Y(n8792) );
	inv_1 U8889( .A(n8774), .Y(n7201) );
	nor2_1 U8890( .A(n11917), .B(n10327), .Y(n8774) );
	a22oi_1 U8891( .A1(g14421), .A2(n10840), .B1(n10228), .B2(n10841), .Y(n8793) );
	o22ai_1 U8892( .A1(n6872), .A2(n6997), .B1(n8794), .B2(n8762), .Y(n8791) );
	inv_1 U8893( .A(g16686), .Y(n6872) );
	o22ai_1 U8894( .A1(n8786), .A2(n7148), .B1(n6543), .B2(n8787), .Y(n8790) );
	inv_1 U8895( .A(n10838), .Y(n6543) );
	nor2_1 U8896( .A(n7202), .B(n6299), .Y(n6602) );
	nor2_1 U8897( .A(n6287), .B(n7196), .Y(n6603) );
	inv_1 U8898( .A(n7202), .Y(n7196) );
	inv_1 U8899( .A(n10836), .Y(n8762) );
	o21ai_0 U8900( .A1(n6245), .A2(n6873), .B1(n8795), .Y(n5262) );
	mux2_1 U8901( .A0(n6478), .A1(n6654), .S(n11889), .X(n8795) );
	nand2_1 U8902( .A(n6339), .B(n6471), .Y(n6654) );
	inv_1 U8903( .A(n6477), .Y(n6471) );
	nand2_1 U8904( .A(n6477), .B(n6333), .Y(n6478) );
	nor4_1 U8905( .A(n8769), .B(n8794), .C(n7198), .D(n7202), .Y(n6477) );
	o21ai_0 U8906( .A1(n6245), .A2(n7739), .B1(n8796), .Y(n5261) );
	a22oi_1 U8907( .A1(n8797), .A2(n8056), .B1(n8051), .B2(n10896), .Y(n8796) );
	xnor2_1 U8908( .A(n8798), .B(n8799), .Y(n8797) );
	nand2_1 U8909( .A(n10896), .B(n8800), .Y(n8798) );
	nand3_1 U8910( .A(g17722), .B(n8801), .C(n10373), .Y(n8800) );
	inv_1 U8911( .A(n10309), .Y(n7739) );
	o221ai_1 U8912( .A1(n8636), .A2(n8802), .B1(n6215), .B2(n6652), .C1(n8803), .Y(n5260) );
	inv_1 U8913( .A(n10504), .Y(n6652) );
	o32ai_1 U8914( .A1(n8804), .A2(n7141), .A3(n7412), .B1(n6367), .B2(n8805), .Y(n5259) );
	inv_1 U8915( .A(n10919), .Y(n8805) );
	inv_1 U8916( .A(n10929), .Y(n7141) );
	o21ai_0 U8917( .A1(n6313), .A2(n6419), .B1(n8806), .Y(n5258) );
	mux2i_1 U8918( .A0(n8807), .A1(n8808), .S(n10514), .Y(n8806) );
	o21ai_0 U8919( .A1(n6368), .A2(n8809), .B1(n6248), .Y(n8808) );
	mux2i_1 U8920( .A0(n8810), .A1(n8811), .S(n6773), .Y(n8809) );
	nor3_1 U8921( .A(n7515), .B(n8811), .C(n8812), .Y(n8810) );
	nor3_1 U8922( .A(n6727), .B(n8813), .C(n6773), .Y(n8807) );
	o21ai_0 U8923( .A1(n6245), .A2(n7439), .B1(n8814), .Y(n5257) );
	mux2i_1 U8924( .A0(n8815), .A1(n7286), .S(n8816), .Y(n8814) );
	nor3_1 U8925( .A(n7442), .B(n10362), .C(n6793), .Y(n8816) );
	nand3_1 U8926( .A(n8817), .B(n8818), .C(n8819), .Y(n7442) );
	nor3_1 U8927( .A(n10288), .B(n10356), .C(n10328), .Y(n8819) );
	nor2_1 U8928( .A(n5953), .B(n6298), .Y(n7286) );
	nor2_1 U8929( .A(n6287), .B(n6032), .Y(n8815) );
	inv_1 U8930( .A(n10858), .Y(n7439) );
	o21ai_0 U8931( .A1(n8036), .A2(n5946), .B1(n8820), .Y(n5256) );
	mux2i_1 U8932( .A0(n8821), .A1(n8822), .S(n10902), .Y(n8820) );
	nand2_1 U8933( .A(n6221), .B(n8823), .Y(n8822) );
	nand3_1 U8934( .A(n6385), .B(n7466), .C(n8824), .Y(n8823) );
	nor2_1 U8935( .A(n7466), .B(n8035), .Y(n8821) );
	nand2_1 U8936( .A(n8824), .B(n6334), .Y(n8035) );
	nor2_1 U8937( .A(n6362), .B(n8825), .Y(n5255) );
	o22ai_1 U8938( .A1(n6205), .A2(n8826), .B1(n8827), .B2(n8232), .Y(n5254) );
	nor4_1 U8939( .A(n8828), .B(n8818), .C(n8829), .D(n8830), .Y(n8827) );
	nand4_1 U8940( .A(n6793), .B(n8831), .C(n6647), .D(n6641), .Y(n8828) );
	inv_1 U8941( .A(n10362), .Y(n6641) );
	inv_1 U8942( .A(n10182), .Y(n6793) );
	inv_1 U8943( .A(n10592), .Y(n8826) );
	o211ai_1 U8944( .A1(n8832), .A2(n8833), .B1(n8834), .C1(n8144), .Y(n5253) );
	nand3_1 U8945( .A(n11905), .B(n8835), .C(n8146), .Y(n8834) );
	a21oi_1 U8946( .A1(n8836), .A2(n8147), .B1(n6437), .Y(n8832) );
	a21oi_1 U8947( .A1(n6198), .A2(n8837), .B1(n5912), .Y(n5252) );
	or2_0 U8948( .A(n7473), .B(n6369), .X(n8837) );
	nor2_1 U8949( .A(n8838), .B(n7474), .Y(n7473) );
	o32ai_1 U8950( .A1(n8434), .A2(n6349), .A3(n8753), .B1(n7646), .B2(n8680), .Y(n5251) );
	nand2_1 U8951( .A(n8753), .B(n6380), .Y(n7646) );
	nor2_1 U8952( .A(n6934), .B(n7653), .Y(n8753) );
	nor3_1 U8953( .A(n10247), .B(n10265), .C(n8431), .Y(n7653) );
	inv_1 U8954( .A(n10477), .Y(n8434) );
	o221ai_1 U8955( .A1(n6745), .A2(n8474), .B1(n6215), .B2(n5918), .C1(n8839), .Y(n5250) );
	a21oi_1 U8956( .A1(n8127), .A2(n10172), .B1(n8840), .Y(n8839) );
	o21ai_0 U8957( .A1(n6043), .A2(n8841), .B1(n8842), .Y(n5249) );
	mux2i_1 U8958( .A0(n8843), .A1(n8844), .S(n10898), .Y(n8842) );
	nand2_1 U8959( .A(n6221), .B(n8845), .Y(n8844) );
	nand3_1 U8960( .A(n6387), .B(n8846), .C(n8847), .Y(n8845) );
	nor2_1 U8961( .A(n8848), .B(n8846), .Y(n8843) );
	o22ai_1 U8962( .A1(n6304), .A2(n7264), .B1(n6194), .B2(n7394), .Y(n5248) );
	o22ai_1 U8963( .A1(n8849), .A2(n6462), .B1(n8850), .B2(n6879), .Y(n5247) );
	a21oi_1 U8964( .A1(n8851), .A2(n6462), .B1(n6460), .Y(n8850) );
	o21ai_0 U8965( .A1(n10668), .A2(n8852), .B1(n8853), .Y(n6460) );
	inv_1 U8966( .A(n10687), .Y(n6462) );
	a21oi_1 U8967( .A1(n6461), .A2(n6879), .B1(n6437), .Y(n8849) );
	and3_1 U8968( .A(n8854), .B(n10668), .C(n10920), .X(n6461) );
	o22ai_1 U8969( .A1(n6303), .A2(n8587), .B1(n6194), .B2(n8855), .Y(n5246) );
	inv_1 U8970( .A(n10878), .Y(n8855) );
	o221ai_1 U8971( .A1(n6454), .A2(n7914), .B1(n6215), .B2(n6077), .C1(n8856), .Y(n5245) );
	or4_1 U8972( .A(n6455), .B(n6313), .C(n6453), .D(n6579), .X(n8856) );
	nand2_1 U8973( .A(n6579), .B(n6333), .Y(n6454) );
	o21ai_0 U8974( .A1(n6245), .A2(n5935), .B1(n8857), .Y(n5244) );
	mux2i_1 U8975( .A0(n8858), .A1(n6255), .S(n8859), .Y(n8857) );
	nor2_1 U8976( .A(n6467), .B(n6570), .Y(n8859) );
	nor2_1 U8977( .A(n6287), .B(n6997), .Y(n8858) );
	inv_1 U8978( .A(n10837), .Y(n6997) );
	o22ai_1 U8979( .A1(n6205), .A2(n8489), .B1(n6305), .B2(n8860), .Y(n5243) );
	mux2i_1 U8980( .A0(n10406), .A1(n8489), .S(n10219), .Y(n8860) );
	o21ai_0 U8981( .A1(n8861), .A2(n6535), .B1(n8862), .Y(n5242) );
	mux2i_1 U8982( .A0(n6437), .A1(n8863), .S(n8285), .Y(n8862) );
	and4_1 U8983( .A(n7746), .B(n10521), .C(n11912), .D(n10916), .X(n8863) );
	inv_1 U8984( .A(n10340), .Y(n6535) );
	a21oi_1 U8985( .A1(n6332), .A2(n8864), .B1(n8289), .Y(n8861) );
	nand3_1 U8986( .A(n10308), .B(n10180), .C(n10372), .Y(n8864) );
	nor2_1 U8987( .A(n6362), .B(n7699), .Y(n5241) );
	inv_1 U8988( .A(g17678), .Y(n7699) );
	o21ai_0 U8989( .A1(n6245), .A2(n7235), .B1(n8865), .Y(n5240) );
	mux2i_1 U8990( .A0(n8866), .A1(n8867), .S(n8868), .Y(n8865) );
	nor2_1 U8991( .A(n10385), .B(n6365), .Y(n8867) );
	nor2_1 U8992( .A(n8048), .B(n8869), .Y(n8866) );
	o22ai_1 U8993( .A1(n6205), .A2(n8718), .B1(n8870), .B2(n8467), .Y(n5239) );
	xnor2_1 U8994( .A(n10515), .B(n8471), .Y(n8870) );
	nor2_1 U8995( .A(n8719), .B(n8718), .Y(n8471) );
	nand2_1 U8996( .A(n8871), .B(n10269), .Y(n8719) );
	o21ai_0 U8997( .A1(n6245), .A2(n5940), .B1(n8872), .Y(n5238) );
	mux2i_1 U8998( .A0(n8873), .A1(n6255), .S(n8874), .Y(n8872) );
	nor2_1 U8999( .A(n6492), .B(n8139), .Y(n8874) );
	nor2_1 U9000( .A(n6286), .B(n8875), .Y(n8873) );
	o221ai_1 U9001( .A1(n8876), .A2(n8877), .B1(n6215), .B2(n7121), .C1(n8878), .Y(tempn5237) );
	o21ai_0 U9002( .A1(n8879), .A2(n6746), .B1(n11865), .Y(n8878) );
	a21oi_1 U9003( .A1(n8880), .A2(n8881), .B1(n6309), .Y(n8879) );
	inv_1 U9004( .A(n10240), .Y(n7121) );
	a21oi_1 U9005( .A1(n8882), .A2(n7432), .B1(n8883), .Y(n8876) );
	nor4_1 U9006( .A(n10251), .B(n7039), .C(n8884), .D(n7460), .Y(n8883) );
	nor2_1 U9007( .A(n8884), .B(n8885), .Y(n7432) );
	a21oi_1 U9008( .A1(n10261), .A2(n7430), .B1(n6309), .Y(n8882) );
	and2_0 U9009( .A(n6345), .B(n10890), .X(n5236) );
	o22ai_1 U9010( .A1(n8886), .A2(n6630), .B1(n6632), .B2(n5950), .Y(n5235) );
	o221ai_1 U9011( .A1(n7880), .A2(n8887), .B1(n6216), .B2(n8888), .C1(n8889), .Y(n5234) );
	or3_1 U9012( .A(n6314), .B(n8167), .C(n8191), .X(n8889) );
	o221ai_1 U9013( .A1(n7768), .A2(n8890), .B1(n6216), .B2(n8891), .C1(n8892), .Y(n5233) );
	nand3_1 U9014( .A(n7772), .B(n6330), .C(n10178), .Y(n8892) );
	o32ai_1 U9015( .A1(n8161), .A2(n6348), .A3(n8160), .B1(n8273), .B2(n7670), .Y(n5232) );
	inv_1 U9016( .A(n10312), .Y(n7670) );
	inv_1 U9017( .A(n10852), .Y(n8161) );
	o32ai_1 U9018( .A1(n8893), .A2(n6348), .A3(n7529), .B1(n7530), .B2(n8448), .Y(n5231) );
	inv_1 U9019( .A(n10629), .Y(n8448) );
	nand2_1 U9020( .A(n7529), .B(n6381), .Y(n7530) );
	nor2_1 U9021( .A(n6934), .B(n7022), .Y(n7529) );
	inv_1 U9022( .A(n10696), .Y(n8893) );
	o21ai_0 U9023( .A1(n6245), .A2(n7935), .B1(n8894), .Y(n5230) );
	a22oi_1 U9024( .A1(n10302), .A2(n7369), .B1(g14096), .B2(n7370), .Y(n8894) );
	o22ai_1 U9025( .A1(n8895), .A2(n8896), .B1(n8897), .B2(n8898), .Y(n5229) );
	o21ai_0 U9026( .A1(n8899), .A2(n10598), .B1(n6342), .Y(n8898) );
	a21oi_1 U9027( .A1(n8900), .A2(n8901), .B1(n8902), .Y(n8899) );
	mux2i_1 U9028( .A0(n8903), .A1(n8904), .S(n8404), .Y(n8901) );
	inv_1 U9029( .A(n10415), .Y(n8404) );
	mux2i_1 U9030( .A0(n8905), .A1(n8906), .S(n5913), .Y(n8900) );
	inv_1 U9031( .A(n8406), .Y(n8895) );
	o221ai_1 U9032( .A1(n7305), .A2(n7486), .B1(n6216), .B2(n7487), .C1(n8907), .Y(n5228) );
	nand3_1 U9033( .A(n7489), .B(n6383), .C(n8908), .Y(n8907) );
	nand2_1 U9034( .A(n7599), .B(n8909), .Y(n7489) );
	nand2_1 U9035( .A(n7742), .B(n6333), .Y(n7486) );
	o21ai_0 U9036( .A1(n6245), .A2(n6468), .B1(n8910), .Y(n5227) );
	mux2i_1 U9037( .A0(n8911), .A1(n6255), .S(n8912), .Y(n8910) );
	nor2_1 U9038( .A(n6286), .B(n7249), .Y(n8911) );
	inv_1 U9039( .A(n10834), .Y(n7249) );
	inv_1 U9040( .A(n10842), .Y(n6468) );
	nor3_1 U9041( .A(n8913), .B(n6351), .C(n8914), .Y(n5226) );
	a21oi_1 U9042( .A1(n10849), .A2(n7395), .B1(n7257), .Y(n8914) );
	nor3_1 U9043( .A(n7738), .B(n7259), .C(n6690), .Y(n8913) );
	inv_1 U9044( .A(n10849), .Y(n7738) );
	o21ai_0 U9045( .A1(n6245), .A2(n8465), .B1(n8915), .Y(n5225) );
	mux2i_1 U9046( .A0(n8916), .A1(n6520), .S(n8917), .Y(n8915) );
	nor2_1 U9047( .A(n10241), .B(n7916), .Y(n8917) );
	nand2_1 U9048( .A(n10252), .B(n6582), .Y(n7916) );
	nor2_1 U9049( .A(n6286), .B(n6000), .Y(n8916) );
	inv_1 U9050( .A(n10723), .Y(n8465) );
	o21ai_0 U9051( .A1(n6245), .A2(n7191), .B1(n8918), .Y(n5224) );
	mux2i_1 U9052( .A0(n8919), .A1(n6255), .S(n8920), .Y(n8918) );
	nor2_1 U9053( .A(n6501), .B(n7186), .Y(n8920) );
	nand2_1 U9054( .A(n10295), .B(n7254), .Y(n6501) );
	nor2_1 U9055( .A(n6286), .B(n6018), .Y(n8919) );
	inv_1 U9056( .A(n10832), .Y(n7191) );
	o21ai_0 U9057( .A1(n6245), .A2(n8921), .B1(n8922), .Y(n5223) );
	mux2i_1 U9058( .A0(n8923), .A1(n6255), .S(n8924), .Y(n8922) );
	nor2_1 U9059( .A(n6789), .B(n8139), .Y(n8924) );
	nor2_1 U9060( .A(n6286), .B(n8135), .Y(n8923) );
	o32ai_1 U9061( .A1(n8500), .A2(n6348), .A3(n8925), .B1(n8926), .B2(n8128), .Y(n5222) );
	inv_1 U9062( .A(n10479), .Y(n8500) );
	nor2_1 U9063( .A(n5874), .B(n8761), .Y(n5221) );
	o21ai_0 U9064( .A1(n6245), .A2(n8083), .B1(n8927), .Y(n5220) );
	mux2i_1 U9065( .A0(n8928), .A1(n6255), .S(n8929), .Y(n8927) );
	nor2_1 U9066( .A(n7496), .B(n7880), .Y(n8929) );
	nor2_1 U9067( .A(n6286), .B(n8930), .Y(n8928) );
	inv_1 U9068( .A(n10752), .Y(n8083) );
	o21ai_0 U9069( .A1(n6245), .A2(n8931), .B1(n8932), .Y(n5219) );
	mux2i_1 U9070( .A0(n8933), .A1(n6255), .S(n8934), .Y(n8932) );
	nor2_1 U9071( .A(n7072), .B(n7965), .Y(n8934) );
	nor2_1 U9072( .A(n6286), .B(n5930), .Y(n8933) );
	o221ai_1 U9073( .A1(n8841), .A2(n8935), .B1(n6216), .B2(n6863), .C1(n8936), .Y(n5218) );
	inv_1 U9074( .A(n10503), .Y(n6863) );
	o21ai_0 U9075( .A1(n6245), .A2(n8937), .B1(n8938), .Y(n5217) );
	mux2i_1 U9076( .A0(n8939), .A1(n6255), .S(n8940), .Y(n8938) );
	nor2_1 U9077( .A(n7071), .B(n8941), .Y(n8940) );
	nor2_1 U9078( .A(n6286), .B(n5982), .Y(n8939) );
	o21ai_0 U9079( .A1(n6245), .A2(n8942), .B1(n8943), .Y(n5216) );
	mux2i_1 U9080( .A0(n8944), .A1(n6255), .S(n8945), .Y(n8943) );
	nor2_1 U9081( .A(n8023), .B(n8250), .Y(n8945) );
	nor2_1 U9082( .A(n6286), .B(n7708), .Y(n8944) );
	o21ai_0 U9083( .A1(n6245), .A2(n6011), .B1(n8946), .Y(n5215) );
	mux2i_1 U9084( .A0(n8947), .A1(n6256), .S(n8948), .Y(n8946) );
	nor2_1 U9085( .A(n7321), .B(n8949), .Y(n8948) );
	nor2_1 U9086( .A(n6286), .B(n8950), .Y(n8947) );
	o21ai_0 U9087( .A1(n6245), .A2(n8951), .B1(n8952), .Y(n5214) );
	mux2i_1 U9088( .A0(n8953), .A1(n7064), .S(n8954), .Y(n8952) );
	nor2_1 U9089( .A(n10239), .B(n7066), .Y(n8954) );
	nand2_1 U9090( .A(n10250), .B(n8499), .Y(n7066) );
	inv_1 U9091( .A(n7884), .Y(n8499) );
	nor2_1 U9092( .A(n6285), .B(n6001), .Y(n8953) );
	o221ai_1 U9093( .A1(n5894), .A2(n8955), .B1(n6216), .B2(n7552), .C1(n8956), .Y(n5213) );
	a21oi_1 U9094( .A1(n8957), .A2(n7626), .B1(n8958), .Y(n8956) );
	nor2_1 U9095( .A(n10331), .B(n7628), .Y(n8957) );
	inv_1 U9096( .A(n10579), .Y(n7552) );
	o221ai_1 U9097( .A1(n6530), .A2(n8959), .B1(n8960), .B2(n8302), .C1(n8961), .Y(n5212) );
	nand3_1 U9098( .A(n8962), .B(n6377), .C(n10550), .Y(n8961) );
	o221ai_1 U9099( .A1(n7895), .A2(n8591), .B1(n6216), .B2(n7221), .C1(n8963), .Y(n5211) );
	or3_1 U9100( .A(n7893), .B(n6369), .C(n6432), .X(n8963) );
	nand2_1 U9101( .A(n10253), .B(n8964), .Y(n6432) );
	inv_1 U9102( .A(n10253), .Y(n7221) );
	nor2_1 U9103( .A(n6362), .B(n8965), .Y(n5210) );
	o21ai_0 U9104( .A1(n6246), .A2(n5936), .B1(n8966), .Y(n5209) );
	mux2i_1 U9105( .A0(n8967), .A1(n6256), .S(n8968), .Y(n8966) );
	nor2_1 U9106( .A(n6971), .B(n7332), .Y(n8968) );
	nor2_1 U9107( .A(n6285), .B(n7989), .Y(n8967) );
	o22ai_1 U9108( .A1(n6204), .A2(n5961), .B1(n7275), .B2(n8969), .Y(n5208) );
	mux2i_1 U9109( .A0(n8970), .A1(n8971), .S(n7390), .Y(n8969) );
	inv_1 U9110( .A(n7276), .Y(n7390) );
	nor4_1 U9111( .A(n5961), .B(n7279), .C(n7281), .D(n7280), .Y(n7276) );
	nor2_1 U9112( .A(n6285), .B(n7391), .Y(n8971) );
	inv_1 U9113( .A(n10893), .Y(n7391) );
	nor2_1 U9114( .A(n10893), .B(n6365), .Y(n8970) );
	nor4_1 U9115( .A(n7392), .B(n7281), .C(n8972), .D(n7393), .Y(n7275) );
	a21oi_1 U9116( .A1(n7787), .A2(n7788), .B1(n8973), .Y(n7393) );
	nor3_1 U9117( .A(n7128), .B(n7401), .C(n5908), .Y(n7788) );
	nor2_1 U9118( .A(n7277), .B(n8974), .Y(n8972) );
	inv_1 U9119( .A(n7280), .Y(n7392) );
	nor3_1 U9120( .A(n8975), .B(n10874), .C(n6484), .Y(n7280) );
	inv_1 U9121( .A(n10468), .Y(n6484) );
	nor2_1 U9122( .A(n6362), .B(n8976), .Y(n5207) );
	o21ai_0 U9123( .A1(n6246), .A2(n7326), .B1(n8977), .Y(n5206) );
	mux2i_1 U9124( .A0(n8978), .A1(n6256), .S(n8979), .Y(n8977) );
	nor2_1 U9125( .A(n6899), .B(n7331), .Y(n8979) );
	nand3_1 U9126( .A(n8980), .B(n5898), .C(n7407), .Y(n7331) );
	nor2_1 U9127( .A(n6285), .B(n6894), .Y(n8978) );
	inv_1 U9128( .A(n10743), .Y(n7326) );
	o211ai_1 U9129( .A1(n8981), .A2(n8982), .B1(n8983), .C1(n6839), .Y(n5205) );
	nand3_1 U9130( .A(n6841), .B(n8984), .C(n11967), .Y(n8983) );
	inv_1 U9131( .A(n8985), .Y(n8984) );
	inv_1 U9132( .A(n10599), .Y(n8982) );
	a21oi_1 U9133( .A1(n8985), .A2(n6843), .B1(n6437), .Y(n8981) );
	o22ai_1 U9134( .A1(n6304), .A2(n6659), .B1(n6194), .B2(n8986), .Y(n5204) );
	o21ai_0 U9135( .A1(n6246), .A2(n5944), .B1(n8300), .Y(n5203) );
	o22ai_1 U9136( .A1(n6073), .A2(n6599), .B1(n8987), .B2(n8988), .Y(n5202) );
	inv_1 U9137( .A(n10932), .Y(n8988) );
	a21oi_1 U9138( .A1(n6598), .A2(n8989), .B1(n6437), .Y(n8987) );
	and2_0 U9139( .A(n6384), .B(g9743), .X(n5201) );
	o21ai_0 U9140( .A1(n6246), .A2(n8615), .B1(n8990), .Y(n5200) );
	mux2i_1 U9141( .A0(n8991), .A1(n6256), .S(n8992), .Y(n8990) );
	nor2_1 U9142( .A(n7570), .B(n6789), .Y(n8992) );
	nor2_1 U9143( .A(n6285), .B(n7957), .Y(n8991) );
	o22ai_1 U9144( .A1(n6810), .A2(n7770), .B1(n7743), .B2(n7546), .Y(n5199) );
	inv_1 U9145( .A(n10339), .Y(n7743) );
	inv_1 U9146( .A(n10355), .Y(n7770) );
	o22ai_1 U9147( .A1(n6206), .A2(n8993), .B1(n8994), .B2(n6869), .Y(n5198) );
	a211oi_1 U9148( .A1(n10351), .A2(n8614), .B1(n8995), .C1(n7781), .Y(n8994) );
	nor2_1 U9149( .A(n8614), .B(n6491), .Y(n7781) );
	nand2_1 U9150( .A(n10204), .B(n8921), .Y(n6491) );
	o21ai_0 U9151( .A1(n6246), .A2(n8996), .B1(n8997), .Y(n5197) );
	o21ai_0 U9152( .A1(n11826), .A2(n7043), .B1(n7237), .Y(n8997) );
	inv_1 U9153( .A(n10587), .Y(n8996) );
	o21ai_0 U9154( .A1(n6246), .A2(n8998), .B1(n8999), .Y(n5196) );
	mux2i_1 U9155( .A0(n9000), .A1(n9001), .S(n8695), .Y(n8999) );
	inv_1 U9156( .A(n10257), .Y(n8695) );
	nor2_1 U9157( .A(n6362), .B(n9002), .Y(n9001) );
	and2_0 U9158( .A(n9002), .B(n6344), .X(n9000) );
	nand3_1 U9159( .A(n8568), .B(n8726), .C(n10908), .Y(n9002) );
	inv_1 U9160( .A(n10908), .Y(n8998) );
	o221ai_1 U9161( .A1(n9003), .A2(n9004), .B1(n6215), .B2(n8734), .C1(n9005), .Y(n5195) );
	o21ai_0 U9162( .A1(n9006), .A2(n6746), .B1(n11862), .Y(n9005) );
	a21oi_1 U9163( .A1(n9007), .A2(n9008), .B1(n6309), .Y(n9006) );
	nand2_1 U9164( .A(n9007), .B(n9008), .Y(n9004) );
	mux2i_1 U9165( .A0(n7601), .A1(n7600), .S(n6562), .Y(n9003) );
	nor2_1 U9166( .A(n6285), .B(n8885), .Y(n7601) );
	a21oi_1 U9167( .A1(n7041), .A2(n9009), .B1(n6309), .Y(n5194) );
	o22ai_1 U9168( .A1(n8525), .A2(n8302), .B1(n9010), .B2(n8526), .Y(n5193) );
	o21ai_0 U9169( .A1(n6246), .A2(n8075), .B1(n9011), .Y(n5192) );
	mux2i_1 U9170( .A0(n9012), .A1(n6256), .S(n9013), .Y(n9011) );
	nor2_1 U9171( .A(n6994), .B(n8074), .Y(n9013) );
	nor2_1 U9172( .A(n6285), .B(n6676), .Y(n9012) );
	inv_1 U9173( .A(n10815), .Y(n6676) );
	o21ai_0 U9174( .A1(n6246), .A2(n5946), .B1(n9014), .Y(n5191) );
	mux2i_1 U9175( .A0(n6662), .A1(n9015), .S(n9016), .Y(n9014) );
	nor2_1 U9176( .A(n6285), .B(n9017), .Y(n9015) );
	inv_1 U9177( .A(n7465), .Y(n6662) );
	o21ai_0 U9178( .A1(n6246), .A2(n7354), .B1(n9018), .Y(n5190) );
	mux2i_1 U9179( .A0(n9019), .A1(n6256), .S(n9020), .Y(n9018) );
	nor2_1 U9180( .A(n7353), .B(n6898), .Y(n9020) );
	nor2_1 U9181( .A(n6285), .B(n6004), .Y(n9019) );
	o22ai_1 U9182( .A1(n6204), .A2(n9021), .B1(n8560), .B2(n9022), .Y(n5189) );
	a222oi_1 U9183( .A1(n4697), .A2(n6994), .B1(n9023), .B2(n6382), .C1(n9024), .C2(n6341), .Y(n9022) );
	o21ai_0 U9184( .A1(n6246), .A2(n8980), .B1(n9025), .Y(n5188) );
	inv_1 U9185( .A(n9026), .Y(n9025) );
	o22ai_1 U9186( .A1(n6972), .A2(n6898), .B1(n7506), .B2(n7667), .Y(n9026) );
	nand2_1 U9187( .A(n10270), .B(n5898), .Y(n6898) );
	inv_1 U9188( .A(n7409), .Y(n6972) );
	a21oi_1 U9189( .A1(n9027), .A2(n8817), .B1(n6368), .Y(n7409) );
	o221ai_1 U9190( .A1(n9028), .A2(n5863), .B1(n6215), .B2(n6938), .C1(n9029), .Y(n5187) );
	nand3_1 U9191( .A(n7663), .B(n9030), .C(n7662), .Y(n9029) );
	xnor2_1 U9192( .A(n6989), .B(n10681), .Y(n9030) );
	inv_1 U9193( .A(n10681), .Y(n6938) );
	a21oi_1 U9194( .A1(n6332), .A2(n6944), .B1(n7661), .Y(n9028) );
	inv_1 U9195( .A(n7663), .Y(n6944) );
	nor2_1 U9196( .A(n6707), .B(n11953), .Y(n7663) );
	o21ai_0 U9197( .A1(n6246), .A2(n6735), .B1(n9031), .Y(n5186) );
	mux2i_1 U9198( .A0(n9032), .A1(n9033), .S(n9034), .Y(n9031) );
	nor2_1 U9199( .A(n6361), .B(n9035), .Y(n9033) );
	nor2_1 U9200( .A(n9036), .B(n6734), .Y(n9032) );
	inv_1 U9201( .A(n9035), .Y(n9036) );
	inv_1 U9202( .A(n10564), .Y(n6735) );
	o221ai_1 U9203( .A1(n9037), .A2(n5867), .B1(n10331), .B2(n9038), .C1(n9039), .Y(n5185) );
	mux2i_1 U9204( .A0(n9040), .A1(n9041), .S(n9042), .Y(n9039) );
	nor4_1 U9205( .A(n7633), .B(n7632), .C(n6744), .D(n9043), .Y(n9041) );
	nand2_1 U9206( .A(n6223), .B(n9038), .Y(n9040) );
	a211oi_1 U9207( .A1(n6330), .A2(n9043), .B1(n7625), .C1(n6746), .Y(n9037) );
	o21ai_0 U9208( .A1(n5932), .A2(n9044), .B1(n9045), .Y(n5184) );
	inv_1 U9209( .A(n6969), .Y(n9045) );
	nor3_1 U9210( .A(n6306), .B(n10431), .C(n6970), .Y(n6969) );
	o21ai_0 U9211( .A1(n6970), .A2(n7571), .B1(n6342), .Y(n9044) );
	inv_1 U9212( .A(n7572), .Y(n6970) );
	o21ai_0 U9213( .A1(n6246), .A2(n9046), .B1(n9047), .Y(n5183) );
	mux2i_1 U9214( .A0(n9048), .A1(n6256), .S(n9049), .Y(n9047) );
	nor2_1 U9215( .A(n6627), .B(n8082), .Y(n9049) );
	nor2_1 U9216( .A(n6285), .B(n7876), .Y(n9048) );
	inv_1 U9217( .A(n10762), .Y(n7876) );
	o32ai_1 U9218( .A1(n5934), .A2(n9050), .A3(n6312), .B1(n9051), .B2(n7401), .Y(n5182) );
	nor2_1 U9219( .A(n9052), .B(n6437), .Y(n9051) );
	nor4_1 U9220( .A(n11829), .B(n6367), .C(n7402), .D(n6438), .Y(n9052) );
	o22ai_1 U9221( .A1(n6203), .A2(n9053), .B1(n6347), .B2(n9054), .Y(n5181) );
	o22ai_1 U9222( .A1(n6204), .A2(n8186), .B1(n9055), .B2(n8025), .Y(n5180) );
	a211oi_1 U9223( .A1(n10350), .A2(n8185), .B1(n9056), .C1(n9057), .Y(n9055) );
	o22ai_1 U9224( .A1(n9058), .A2(n8833), .B1(n8835), .B2(n9059), .Y(n5179) );
	o21ai_0 U9225( .A1(n9060), .A2(n10595), .B1(n6341), .Y(n9059) );
	a21oi_1 U9226( .A1(n9061), .A2(n9062), .B1(n9063), .Y(n9060) );
	mux2i_1 U9227( .A0(n9064), .A1(n9065), .S(n6829), .Y(n9062) );
	inv_1 U9228( .A(n10419), .Y(n6829) );
	mux2i_1 U9229( .A0(n9066), .A1(n9067), .S(n5917), .Y(n9061) );
	inv_1 U9230( .A(n8836), .Y(n8835) );
	nor2_1 U9231( .A(n9068), .B(n8231), .Y(n8836) );
	inv_1 U9232( .A(n10595), .Y(n8833) );
	inv_1 U9233( .A(n6831), .Y(n9058) );
	o22ai_1 U9234( .A1(n6631), .A2(n6630), .B1(n9069), .B2(n6632), .Y(n5178) );
	inv_1 U9235( .A(n10358), .Y(n6631) );
	o21ai_0 U9236( .A1(n6246), .A2(n5943), .B1(n9070), .Y(n5177) );
	mux2_1 U9237( .A0(n9071), .A1(n6960), .S(n10692), .X(n9070) );
	o32ai_1 U9238( .A1(n6310), .A2(n9072), .A3(n9073), .B1(n6201), .B2(n7840), .Y(n5176) );
	a21oi_1 U9239( .A1(n9074), .A2(n6771), .B1(n10582), .Y(n9073) );
	nor4_1 U9240( .A(n10240), .B(n9075), .C(n7430), .D(n9076), .Y(n9072) );
	o21ai_0 U9241( .A1(n8955), .A2(n9077), .B1(n9078), .Y(n5175) );
	mux2i_1 U9242( .A0(n9079), .A1(n9080), .S(n10553), .Y(n9078) );
	nand2_1 U9243( .A(n6223), .B(n9081), .Y(n9080) );
	nand3_1 U9244( .A(n9082), .B(n6379), .C(n9083), .Y(n9081) );
	nor2_1 U9245( .A(n6285), .B(n9082), .Y(n9079) );
	nand2_1 U9246( .A(n10674), .B(n9084), .Y(n9082) );
	o221ai_1 U9247( .A1(n9085), .A2(n9086), .B1(n6215), .B2(n9087), .C1(n9088), .Y(n5174) );
	o21ai_0 U9248( .A1(n9089), .A2(n6746), .B1(n11867), .Y(n9088) );
	inv_1 U9249( .A(n9090), .Y(n9089) );
	o21ai_0 U9250( .A1(n9086), .A2(n9091), .B1(n6342), .Y(n9090) );
	a21oi_1 U9251( .A1(n9092), .A2(n9093), .B1(n9094), .Y(n9085) );
	nor4_1 U9252( .A(n10254), .B(n7039), .C(n9091), .D(n7449), .Y(n9094) );
	a21oi_1 U9253( .A1(n10264), .A2(n7956), .B1(n6309), .Y(n9092) );
	o21ai_0 U9254( .A1(n6246), .A2(n9095), .B1(n9096), .Y(n5173) );
	mux2i_1 U9255( .A0(n9097), .A1(n7303), .S(n9098), .Y(n9096) );
	nor2_1 U9256( .A(n10266), .B(n8659), .Y(n9098) );
	inv_1 U9257( .A(n8908), .Y(n8659) );
	nor2_1 U9258( .A(n7487), .B(n7742), .Y(n8908) );
	nor2_1 U9259( .A(n6284), .B(n5983), .Y(n9097) );
	o221ai_1 U9260( .A1(n7632), .A2(n8955), .B1(n6214), .B2(n5867), .C1(n9099), .Y(n5172) );
	a21oi_1 U9261( .A1(n7626), .A2(n10299), .B1(n8958), .Y(n9099) );
	inv_1 U9262( .A(n10331), .Y(n7632) );
	o21ai_0 U9263( .A1(n6246), .A2(n9100), .B1(n9101), .Y(n5171) );
	mux2i_1 U9264( .A0(n9102), .A1(n9103), .S(n9104), .Y(n9101) );
	nor2_1 U9265( .A(n10532), .B(n6364), .Y(n9103) );
	nor2_1 U9266( .A(n8309), .B(n7108), .Y(n9102) );
	inv_1 U9267( .A(n10532), .Y(n8309) );
	nor3_1 U9268( .A(n9105), .B(n6351), .C(n9106), .Y(n5170) );
	a21oi_1 U9269( .A1(n10855), .A2(n7464), .B1(n7257), .Y(n9106) );
	nor3_1 U9270( .A(n7463), .B(n7259), .C(n6663), .Y(n9105) );
	inv_1 U9271( .A(n10855), .Y(n7463) );
	o221ai_1 U9272( .A1(n7809), .A2(n7813), .B1(n6214), .B2(n8403), .C1(n7815), .Y(n5169) );
	nand3_1 U9273( .A(n9107), .B(n6376), .C(n10321), .Y(n7815) );
	inv_1 U9274( .A(n10321), .Y(n8403) );
	inv_1 U9275( .A(n10634), .Y(n7813) );
	o21ai_0 U9276( .A1(n6247), .A2(n9108), .B1(n9109), .Y(n5168) );
	mux2i_1 U9277( .A0(n9110), .A1(n9111), .S(n5914), .Y(n9109) );
	nor2_1 U9278( .A(n6361), .B(n9112), .Y(n9111) );
	nor2_1 U9279( .A(n8744), .B(n6734), .Y(n9110) );
	inv_1 U9280( .A(n9112), .Y(n8744) );
	nand2_1 U9281( .A(n10539), .B(n9113), .Y(n9112) );
	o221ai_1 U9282( .A1(n6587), .A2(n5889), .B1(n6214), .B2(n7137), .C1(n9114), .Y(n5167) );
	a21oi_1 U9283( .A1(n9115), .A2(n6590), .B1(n6591), .Y(n9114) );
	nor2_1 U9284( .A(n7954), .B(n6300), .Y(n6590) );
	nor2_1 U9285( .A(n10337), .B(n7360), .Y(n9115) );
	nor2_1 U9286( .A(n7793), .B(n11958), .Y(n7360) );
	inv_1 U9287( .A(n10585), .Y(n7137) );
	inv_1 U9288( .A(n7358), .Y(n6587) );
	o211ai_1 U9289( .A1(n6203), .A2(n9116), .B1(n9117), .C1(n9118), .Y(n5166) );
	nand3_1 U9290( .A(n9119), .B(n6648), .C(n9120), .Y(n9118) );
	nor2_1 U9291( .A(n7207), .B(n6366), .Y(n6648) );
	nand3_1 U9292( .A(n10342), .B(n9121), .C(n6794), .Y(n9117) );
	o21ai_0 U9293( .A1(n6246), .A2(n5921), .B1(n9122), .Y(n5165) );
	mux2i_1 U9294( .A0(n9123), .A1(n6256), .S(n9124), .Y(n9122) );
	nor2_1 U9295( .A(n6808), .B(n6995), .Y(n9124) );
	nor2_1 U9296( .A(n6284), .B(n6990), .Y(n9123) );
	nor2_1 U9297( .A(n6361), .B(n9125), .Y(n5164) );
	o22ai_1 U9298( .A1(n6204), .A2(n8641), .B1(n6297), .B2(n9126), .Y(n5163) );
	mux2i_1 U9299( .A0(n9127), .A1(n10901), .S(n9128), .Y(n9126) );
	xnor2_1 U9300( .A(n9129), .B(n8330), .Y(n9127) );
	nand2_1 U9301( .A(n9130), .B(n9131), .Y(n8330) );
	mux2i_1 U9302( .A0(n9132), .A1(n9133), .S(n9134), .Y(n9131) );
	xnor2_1 U9303( .A(n9135), .B(g11418), .Y(n9134) );
	nand3_1 U9304( .A(n9136), .B(n9137), .C(n9138), .Y(n9133) );
	nand3_1 U9305( .A(g16775), .B(n11800), .C(n9139), .Y(n9138) );
	nand3_1 U9306( .A(g16659), .B(n9140), .C(n10498), .Y(n9137) );
	nand3_1 U9307( .A(g13966), .B(n11811), .C(n9141), .Y(n9136) );
	nand3_1 U9308( .A(n9142), .B(n9143), .C(n9144), .Y(n9132) );
	nand3_1 U9309( .A(n9145), .B(n11873), .C(g16775), .Y(n9144) );
	nand3_1 U9310( .A(n9140), .B(n11874), .C(g13966), .Y(n9143) );
	nand3_1 U9311( .A(n9141), .B(n10816), .C(g16659), .Y(n9142) );
	mux2_1 U9312( .A0(n9146), .A1(n9147), .S(n9135), .X(n9130) );
	a221oi_1 U9313( .A1(n9139), .A2(n9148), .B1(n9145), .B2(n9149), .C1(n9150), .Y(n9147) );
	o32ai_1 U9314( .A1(n9151), .A2(n5921), .A3(n9152), .B1(n9153), .B2(n9154), .Y(n9150) );
	a22oi_1 U9315( .A1(g14518), .A2(n10804), .B1(n10226), .B2(n10805), .Y(n9153) );
	o22ai_1 U9316( .A1(n7382), .A2(n9155), .B1(n8162), .B2(n9156), .Y(n9149) );
	inv_1 U9317( .A(n10807), .Y(n7382) );
	o22ai_1 U9318( .A1(n6990), .A2(n7917), .B1(n9157), .B2(n9158), .Y(n9148) );
	inv_1 U9319( .A(n10809), .Y(n6990) );
	a221oi_1 U9320( .A1(n9139), .A2(n9159), .B1(n9145), .B2(n9160), .C1(n9161), .Y(n9146) );
	o32ai_1 U9321( .A1(n9151), .A2(n5923), .A3(n9154), .B1(n9162), .B2(n9152), .Y(n9161) );
	inv_1 U9322( .A(n9141), .Y(n9152) );
	a22oi_1 U9323( .A1(n10814), .A2(g14518), .B1(n10226), .B2(n10815), .Y(n9162) );
	o22ai_1 U9324( .A1(n7917), .A2(n8075), .B1(n9157), .B2(n8328), .Y(n9160) );
	inv_1 U9325( .A(n10810), .Y(n8328) );
	inv_1 U9326( .A(n10811), .Y(n8075) );
	inv_1 U9327( .A(g16748), .Y(n7917) );
	o22ai_1 U9328( .A1(n9155), .A2(n9163), .B1(n6682), .B2(n9156), .Y(n9159) );
	inv_1 U9329( .A(n10812), .Y(n6682) );
	nand2_1 U9330( .A(n10901), .B(n9164), .Y(n9129) );
	nand3_1 U9331( .A(n10377), .B(n9145), .C(g16693), .Y(n9164) );
	o22ai_1 U9332( .A1(n6810), .A2(n8708), .B1(n7546), .B2(n6085), .Y(n5162) );
	o32ai_1 U9333( .A1(n6310), .A2(n10415), .A3(n8668), .B1(n6201), .B2(n9165), .Y(n5161) );
	nor2_1 U9334( .A(n9165), .B(n9166), .Y(n8668) );
	o22ai_1 U9335( .A1(n6810), .A2(n7744), .B1(n7546), .B2(n7984), .Y(n5160) );
	inv_1 U9336( .A(n10882), .Y(n7984) );
	inv_1 U9337( .A(n10734), .Y(n7744) );
	o21ai_0 U9338( .A1(n6247), .A2(n7938), .B1(n9167), .Y(n5159) );
	a22oi_1 U9339( .A1(n10187), .A2(n7369), .B1(g14147), .B2(n7370), .Y(n9167) );
	o32ai_1 U9340( .A1(n6310), .A2(g9615), .A3(n9168), .B1(n6201), .B2(n9169), .Y(n5158) );
	a21oi_1 U9341( .A1(g9555), .A2(n9169), .B1(n10612), .Y(n9168) );
	inv_1 U9342( .A(n10611), .Y(n9169) );
	o22ai_1 U9343( .A1(n6204), .A2(n6833), .B1(n9170), .B2(n9171), .Y(n5157) );
	o21ai_0 U9344( .A1(n9065), .A2(n9172), .B1(n6382), .Y(n9171) );
	a21oi_1 U9345( .A1(n9173), .A2(n9174), .B1(n6934), .Y(n9172) );
	mux2i_1 U9346( .A0(n6834), .A1(n10196), .S(n9063), .Y(n9170) );
	nand2_1 U9347( .A(n9175), .B(n8262), .Y(n6834) );
	o21ai_0 U9348( .A1(n6246), .A2(n9176), .B1(n9177), .Y(n5156) );
	a22oi_1 U9349( .A1(n11831), .A2(n6831), .B1(n6835), .B2(n9178), .Y(n9177) );
	o21ai_0 U9350( .A1(n6247), .A2(n9179), .B1(n9180), .Y(n5155) );
	a22oi_1 U9351( .A1(n7136), .A2(n6754), .B1(n10843), .B2(n7138), .Y(n9180) );
	inv_1 U9352( .A(n10580), .Y(n6754) );
	o22ai_1 U9353( .A1(n7768), .A2(n8891), .B1(n8705), .B2(n9181), .Y(n5154) );
	inv_1 U9354( .A(n10433), .Y(n8891) );
	o22ai_1 U9355( .A1(n6204), .A2(n9182), .B1(n9183), .B2(n6297), .Y(n5153) );
	a21oi_1 U9356( .A1(n9184), .A2(n9185), .B1(n9186), .Y(n9183) );
	nor4_1 U9357( .A(n10879), .B(n10526), .C(n10185), .D(g26885), .Y(n9186) );
	nand2_1 U9358( .A(n9187), .B(n7411), .Y(n9185) );
	inv_1 U9359( .A(g26885), .Y(n7411) );
	mux2i_1 U9360( .A0(n10185), .A1(n10526), .S(n6977), .Y(n9187) );
	inv_1 U9361( .A(n10549), .Y(n6977) );
	inv_1 U9362( .A(n8600), .Y(n9184) );
	inv_1 U9363( .A(n10879), .Y(n9182) );
	o22ai_1 U9364( .A1(n6205), .A2(n6496), .B1(n9188), .B2(n6298), .Y(n5152) );
	nor4_1 U9365( .A(n10655), .B(n10447), .C(n10444), .D(n7043), .Y(n9188) );
	o21ai_0 U9366( .A1(n6247), .A2(n8267), .B1(n9189), .Y(n5151) );
	mux2i_1 U9367( .A0(n9190), .A1(n6256), .S(n9191), .Y(n9189) );
	nor2_1 U9368( .A(n7228), .B(n8266), .Y(n9191) );
	nor2_1 U9369( .A(n6284), .B(n6901), .Y(n9190) );
	o32ai_1 U9370( .A1(n5905), .A2(n8287), .A3(n9192), .B1(n9193), .B2(n8290), .Y(n5150) );
	a21oi_1 U9371( .A1(n9194), .A2(n7057), .B1(n6437), .Y(n9193) );
	nor2_1 U9372( .A(n8287), .B(n6366), .Y(n7057) );
	nor2_1 U9373( .A(n11913), .B(n9195), .Y(n9194) );
	a21oi_1 U9374( .A1(n6332), .A2(n8290), .B1(n8289), .Y(n9192) );
	inv_1 U9375( .A(n10521), .Y(n8290) );
	o32ai_1 U9376( .A1(n9196), .A2(n6348), .A3(n8282), .B1(n6200), .B2(n5948), .Y(n5149) );
	mux2i_1 U9377( .A0(n9197), .A1(n9198), .S(n8286), .Y(n9196) );
	nor2_1 U9378( .A(n8283), .B(n5948), .Y(n9198) );
	a21oi_1 U9379( .A1(n11940), .A2(n9199), .B1(n6934), .Y(n9197) );
	mux2i_1 U9380( .A0(n9200), .A1(n9201), .S(n6674), .Y(n5148) );
	or2_0 U9381( .A(n8484), .B(n9202), .X(n9201) );
	a21oi_1 U9382( .A1(n9203), .A2(n9202), .B1(n6437), .Y(n9200) );
	inv_1 U9383( .A(n9204), .Y(n5147) );
	a21oi_1 U9384( .A1(n6616), .A2(n11931), .B1(n9205), .Y(n9204) );
	mux2_1 U9385( .A0(n9206), .A1(n9207), .S(n10636), .X(n9205) );
	nand2_1 U9386( .A(n6222), .B(n6618), .Y(n9207) );
	nand3_1 U9387( .A(n9208), .B(n6382), .C(n10323), .Y(n6618) );
	nor2_1 U9388( .A(n10323), .B(n8572), .Y(n9206) );
	o22ai_1 U9389( .A1(n6206), .A2(n9209), .B1(n8690), .B2(n9210), .Y(n5146) );
	a222oi_1 U9390( .A1(n4696), .A2(n7228), .B1(n9211), .B2(n6382), .C1(n9212), .C2(n6341), .Y(n9210) );
	o22ai_1 U9391( .A1(n6204), .A2(n9213), .B1(n9214), .B2(n9215), .Y(n5145) );
	o21ai_0 U9392( .A1(n9139), .A2(n9216), .B1(n6382), .Y(n9215) );
	a21oi_1 U9393( .A1(n8331), .A2(n9154), .B1(n6934), .Y(n9216) );
	inv_1 U9394( .A(n9140), .Y(n9154) );
	mux2i_1 U9395( .A0(n9217), .A1(n10195), .S(n9128), .Y(n9214) );
	nor2_1 U9396( .A(n6360), .B(n9218), .Y(n5144) );
	and2_0 U9397( .A(n6384), .B(g8416), .X(n5143) );
	o21ai_0 U9398( .A1(n6247), .A2(n7545), .B1(n9219), .Y(n5142) );
	a22oi_1 U9399( .A1(n10178), .A2(n7746), .B1(n11761), .B2(n8289), .Y(n9219) );
	nor2_1 U9400( .A(n6361), .B(n9220), .Y(n5141) );
	o211ai_1 U9401( .A1(n6203), .A2(n8829), .B1(n8232), .C1(n9221), .Y(n5140) );
	mux2i_1 U9402( .A0(n9222), .A1(n9223), .S(n9224), .Y(n9221) );
	nor2_1 U9403( .A(n6360), .B(n9225), .Y(n9223) );
	and2_0 U9404( .A(n9225), .B(n6344), .X(n9222) );
	nor2_1 U9405( .A(n6284), .B(n8094), .Y(n5139) );
	inv_1 U9406( .A(n10167), .Y(n8094) );
	o21ai_0 U9407( .A1(n6247), .A2(n8677), .B1(n9226), .Y(n5138) );
	mux2i_1 U9408( .A0(n9227), .A1(n9228), .S(n9229), .Y(n9226) );
	nor2_1 U9409( .A(n10533), .B(n6365), .Y(n9228) );
	nor2_1 U9410( .A(n9100), .B(n7108), .Y(n9227) );
	inv_1 U9411( .A(n10533), .Y(n9100) );
	o221ai_1 U9412( .A1(n8014), .A2(n8735), .B1(n6213), .B2(n9230), .C1(n9231), .Y(n5137) );
	nand3_1 U9413( .A(n8738), .B(n6376), .C(n8236), .Y(n9231) );
	nor2_1 U9414( .A(n9230), .B(n8431), .Y(n8236) );
	o21ai_0 U9415( .A1(n6247), .A2(n5998), .B1(n9232), .Y(n5136) );
	mux2i_1 U9416( .A0(n9233), .A1(n6430), .S(n9234), .Y(n9232) );
	nor2_1 U9417( .A(n7895), .B(n7983), .Y(n9234) );
	inv_1 U9418( .A(n9235), .Y(n7983) );
	nor2_1 U9419( .A(n6281), .B(n7985), .Y(n9233) );
	inv_1 U9420( .A(n10724), .Y(n7985) );
	o21ai_0 U9421( .A1(n6247), .A2(n6420), .B1(n9236), .Y(n5135) );
	mux2i_1 U9422( .A0(n9237), .A1(n9238), .S(n6410), .Y(n9236) );
	nand2_1 U9423( .A(n6774), .B(n9239), .Y(n9238) );
	nand3_1 U9424( .A(n10177), .B(n6371), .C(n6779), .Y(n9239) );
	inv_1 U9425( .A(n6421), .Y(n6779) );
	nand3_1 U9426( .A(n6340), .B(n6420), .C(n6778), .Y(n6774) );
	nor2_1 U9427( .A(n9240), .B(n6727), .Y(n9237) );
	mux2i_1 U9428( .A0(n6421), .A1(n6419), .S(n6420), .Y(n9240) );
	inv_1 U9429( .A(n6778), .Y(n6419) );
	nor3_1 U9430( .A(n10360), .B(n10514), .C(n7265), .Y(n6778) );
	nand3_1 U9431( .A(n8811), .B(n10360), .C(n10514), .Y(n6421) );
	o221ai_1 U9432( .A1(n7956), .A2(n9241), .B1(n6213), .B2(n6076), .C1(n9242), .Y(n5134) );
	or4_1 U9433( .A(n9087), .B(n6314), .C(n9093), .D(n9243), .X(n9242) );
	o21ai_0 U9434( .A1(n6960), .A2(n6095), .B1(n9244), .Y(n5133) );
	mux2i_1 U9435( .A0(n9245), .A1(n9246), .S(n10633), .Y(n9244) );
	nand2_1 U9436( .A(n6223), .B(n6963), .Y(n9246) );
	nand3_1 U9437( .A(n9247), .B(n6376), .C(n10320), .Y(n6963) );
	nor2_1 U9438( .A(n10320), .B(n9071), .Y(n9245) );
	or2_0 U9439( .A(n6314), .B(n9247), .X(n6960) );
	nor2_1 U9440( .A(n6284), .B(n9248), .Y(n5132) );
	o21ai_0 U9441( .A1(n6247), .A2(n5999), .B1(n9249), .Y(n5131) );
	mux2i_1 U9442( .A0(n9250), .A1(n6256), .S(n9251), .Y(n9249) );
	nor2_1 U9443( .A(n6492), .B(n7570), .Y(n9251) );
	nor2_1 U9444( .A(n6284), .B(n6639), .Y(n9250) );
	inv_1 U9445( .A(n10497), .Y(n6639) );
	o21ai_0 U9446( .A1(n6247), .A2(n9252), .B1(n9253), .Y(n5130) );
	a22oi_1 U9447( .A1(n10463), .A2(n7369), .B1(g14217), .B2(n7370), .Y(n9253) );
	inv_1 U9448( .A(n10459), .Y(n9252) );
	o21ai_0 U9449( .A1(n6247), .A2(n9254), .B1(n9255), .Y(n5129) );
	mux2i_1 U9450( .A0(n9256), .A1(n6256), .S(n9257), .Y(n9255) );
	nor2_1 U9451( .A(n6858), .B(n8082), .Y(n9257) );
	nor2_1 U9452( .A(n6283), .B(n9258), .Y(n9256) );
	o21ai_0 U9453( .A1(n6247), .A2(n9259), .B1(n9260), .Y(n5128) );
	a22oi_1 U9454( .A1(n11832), .A2(n9261), .B1(n9262), .B2(n9263), .Y(n9260) );
	o22ai_1 U9455( .A1(n6305), .A2(n9264), .B1(n9265), .B2(n7144), .Y(n5127) );
	inv_1 U9456( .A(n10933), .Y(n7144) );
	a21oi_1 U9457( .A1(n9266), .A2(n9267), .B1(n6437), .Y(n9265) );
	inv_1 U9458( .A(n8804), .Y(n9267) );
	nor2_1 U9459( .A(n6360), .B(n9268), .Y(n9266) );
	o21ai_0 U9460( .A1(n6982), .A2(n6051), .B1(n9269), .Y(n5126) );
	mux2i_1 U9461( .A0(n9270), .A1(n9271), .S(n6983), .Y(n9269) );
	inv_1 U9462( .A(n10624), .Y(n6983) );
	nor3_1 U9463( .A(n7523), .B(n10691), .C(n6306), .Y(n9271) );
	inv_1 U9464( .A(n9272), .Y(n7523) );
	nand2_1 U9465( .A(n6224), .B(n9273), .Y(n9270) );
	nand3_1 U9466( .A(n10691), .B(n6376), .C(n9272), .Y(n9273) );
	o32ai_1 U9467( .A1(n6310), .A2(n9274), .A3(n9275), .B1(n6200), .B2(n7630), .Y(n5125) );
	inv_1 U9468( .A(n10486), .Y(n7630) );
	a21oi_1 U9469( .A1(n7627), .A2(n9083), .B1(n10579), .Y(n9275) );
	nor4_1 U9470( .A(n10247), .B(n7633), .C(n9230), .D(n9276), .Y(n9274) );
	o22ai_1 U9471( .A1(n6204), .A2(n5907), .B1(n6298), .B2(n9277), .Y(n5124) );
	mux2i_1 U9472( .A0(n9278), .A1(n10423), .S(n7425), .Y(n9277) );
	nor2_1 U9473( .A(n10423), .B(n7424), .Y(n9278) );
	o21ai_0 U9474( .A1(n6247), .A2(n9279), .B1(n9280), .Y(n5123) );
	a22oi_1 U9475( .A1(n9281), .A2(n10758), .B1(n9282), .B2(n6249), .Y(n9280) );
	o21ai_0 U9476( .A1(n6247), .A2(n9283), .B1(n9284), .Y(n5122) );
	mux2i_1 U9477( .A0(n9285), .A1(n6256), .S(n9286), .Y(n9284) );
	nor2_1 U9478( .A(n7880), .B(n9287), .Y(n9286) );
	nor2_1 U9479( .A(n6283), .B(n6012), .Y(n9285) );
	o22ai_1 U9480( .A1(n6305), .A2(n9288), .B1(n9289), .B2(n9290), .Y(n5121) );
	inv_1 U9481( .A(n10519), .Y(n9290) );
	a21oi_1 U9482( .A1(n9291), .A2(n6380), .B1(n6437), .Y(n9289) );
	o21ai_0 U9483( .A1(n6247), .A2(n9292), .B1(n9293), .Y(n5120) );
	mux2i_1 U9484( .A0(n9294), .A1(n6256), .S(n9295), .Y(n9293) );
	nor2_1 U9485( .A(n7485), .B(n8074), .Y(n9295) );
	nand2_1 U9486( .A(n10275), .B(n5901), .Y(n7485) );
	nor2_1 U9487( .A(n6283), .B(n9163), .Y(n9294) );
	o32ai_1 U9488( .A1(n6310), .A2(g8398), .A3(n9296), .B1(n6200), .B2(n9297), .Y(n5119) );
	a21oi_1 U9489( .A1(g8344), .A2(n9297), .B1(n10616), .Y(n9296) );
	inv_1 U9490( .A(n10615), .Y(n9297) );
	o21ai_0 U9491( .A1(n6248), .A2(n7709), .B1(n9298), .Y(n5118) );
	mux2i_1 U9492( .A0(n9299), .A1(n6257), .S(n9300), .Y(n9298) );
	nor2_1 U9493( .A(n8023), .B(n8099), .Y(n9300) );
	nor2_1 U9494( .A(n6283), .B(n6014), .Y(n9299) );
	inv_1 U9495( .A(n10786), .Y(n7709) );
	o32ai_1 U9496( .A1(n8557), .A2(n10157), .A3(n6808), .B1(n6200), .B2(n5901), .Y(n5117) );
	inv_1 U9497( .A(n9301), .Y(n8557) );
	o221ai_1 U9498( .A1(n9302), .A2(n9303), .B1(n6212), .B2(n6455), .C1(n9304), .Y(n5116) );
	o21ai_0 U9499( .A1(n9305), .A2(n6746), .B1(n11869), .Y(n9304) );
	inv_1 U9500( .A(n9306), .Y(n9305) );
	o21ai_0 U9501( .A1(n9303), .A2(n9307), .B1(n6341), .Y(n9306) );
	a21oi_1 U9502( .A1(n9308), .A2(n6453), .B1(n9309), .Y(n9302) );
	nor4_1 U9503( .A(n10252), .B(n9307), .C(n6573), .D(n7039), .Y(n9309) );
	inv_1 U9504( .A(n7600), .Y(n7039) );
	nor2_1 U9505( .A(n6973), .B(n10165), .Y(n7600) );
	nor2_1 U9506( .A(n8885), .B(n9307), .Y(n6453) );
	a21oi_1 U9507( .A1(n10262), .A2(n7914), .B1(n6305), .Y(n9308) );
	inv_1 U9508( .A(n10252), .Y(n7914) );
	o21ai_0 U9509( .A1(n6247), .A2(n5924), .B1(n9310), .Y(n5115) );
	mux2i_1 U9510( .A0(n9311), .A1(n6257), .S(n9312), .Y(n9310) );
	nor2_1 U9511( .A(n7026), .B(n7229), .Y(n9312) );
	nor2_1 U9512( .A(n6283), .B(n7224), .Y(n9311) );
	inv_1 U9513( .A(n10770), .Y(n7224) );
	o21ai_0 U9514( .A1(n6248), .A2(n7536), .B1(n9313), .Y(n5114) );
	a22oi_1 U9515( .A1(n7136), .A2(n9314), .B1(n10844), .B2(n7138), .Y(n9313) );
	a21oi_1 U9516( .A1(n10235), .A2(n9315), .B1(n6303), .Y(n7138) );
	nor3_1 U9517( .A(n9315), .B(n9316), .C(n6306), .Y(n7136) );
	inv_1 U9518( .A(n10845), .Y(n7536) );
	o21ai_0 U9519( .A1(n6247), .A2(n5984), .B1(n9317), .Y(n5113) );
	mux2i_1 U9520( .A0(n9318), .A1(n7064), .S(n9319), .Y(n9317) );
	nor2_1 U9521( .A(n7111), .B(n9320), .Y(n9319) );
	nor2_1 U9522( .A(n6282), .B(n8951), .Y(n9318) );
	inv_1 U9523( .A(n10721), .Y(n8951) );
	o22ai_1 U9524( .A1(n9021), .A2(n8527), .B1(n9321), .B2(n6994), .Y(n5112) );
	a21oi_1 U9525( .A1(n9301), .A2(n9021), .B1(n6437), .Y(n9321) );
	nor2_1 U9526( .A(n8560), .B(n6366), .Y(n9301) );
	or3_1 U9527( .A(n8560), .B(n10157), .C(n6309), .X(n8527) );
	nor3_1 U9528( .A(n9322), .B(n9323), .C(n9116), .Y(n8560) );
	o21ai_0 U9529( .A1(n6248), .A2(n6000), .B1(n9324), .Y(n5111) );
	mux2i_1 U9530( .A0(n9325), .A1(n6520), .S(n9326), .Y(n9324) );
	nor3_1 U9531( .A(n6573), .B(n6579), .C(n6455), .Y(n9326) );
	inv_1 U9532( .A(n10241), .Y(n6455) );
	nor2_1 U9533( .A(n6282), .B(n6853), .Y(n9325) );
	inv_1 U9534( .A(n10490), .Y(n6853) );
	o21ai_0 U9535( .A1(n6248), .A2(n6003), .B1(n9327), .Y(n5110) );
	mux2i_1 U9536( .A0(n9328), .A1(n6257), .S(n9329), .Y(n9327) );
	nor2_1 U9537( .A(n6971), .B(n7669), .Y(n9329) );
	nor2_1 U9538( .A(n6282), .B(n7322), .Y(n9328) );
	inv_1 U9539( .A(n10751), .Y(n7322) );
	o21ai_0 U9540( .A1(n6248), .A2(n8846), .B1(n9330), .Y(n5109) );
	a22oi_1 U9541( .A1(n9331), .A2(n8411), .B1(n10898), .B2(n8406), .Y(n9330) );
	xnor2_1 U9542( .A(n9332), .B(n9333), .Y(n9331) );
	nand2_1 U9543( .A(n10898), .B(n9334), .Y(n9332) );
	nand3_1 U9544( .A(n10375), .B(n8903), .C(g17646), .Y(n9334) );
	o221ai_1 U9545( .A1(n9335), .A2(n5873), .B1(n10334), .B2(n8239), .C1(n9336), .Y(n5108) );
	mux2i_1 U9546( .A0(n9337), .A1(n9338), .S(n8238), .Y(n9336) );
	nor4_1 U9547( .A(n6744), .B(n9075), .C(n9339), .D(n7584), .Y(n9338) );
	nand2_1 U9548( .A(n6224), .B(n8239), .Y(n9337) );
	inv_1 U9549( .A(n7587), .Y(n8239) );
	nor3_1 U9550( .A(n9075), .B(n7657), .C(n9339), .Y(n7587) );
	a211oi_1 U9551( .A1(n6330), .A2(n9339), .B1(n6746), .C1(n8240), .Y(n9335) );
	o22ai_1 U9552( .A1(n6205), .A2(n6597), .B1(n9340), .B2(n6599), .Y(n5107) );
	xnor2_1 U9553( .A(n10932), .B(n8989), .Y(n9340) );
	inv_1 U9554( .A(n10189), .Y(n6597) );
	and2_0 U9555( .A(n6384), .B(g9497), .X(n5106) );
	o21ai_0 U9556( .A1(n6248), .A2(n6001), .B1(n9341), .Y(n5105) );
	mux2i_1 U9557( .A0(n9342), .A1(n7064), .S(n9343), .Y(n9341) );
	nor3_1 U9558( .A(n7883), .B(n7884), .C(n7111), .Y(n9343) );
	inv_1 U9559( .A(n10260), .Y(n7111) );
	nor2_1 U9560( .A(n6282), .B(n7086), .Y(n9342) );
	o21ai_0 U9561( .A1(n7179), .A2(n7182), .B1(n9344), .Y(n5104) );
	mux2i_1 U9562( .A0(n9345), .A1(n9346), .S(n10643), .Y(n9344) );
	nand2_1 U9563( .A(n6225), .B(n9347), .Y(n9346) );
	nor2_1 U9564( .A(n10685), .B(n7181), .Y(n9345) );
	nand2_1 U9565( .A(n7502), .B(n6335), .Y(n7181) );
	o221ai_1 U9566( .A1(n9348), .A2(n6304), .B1(n6217), .B2(n7895), .C1(n9349), .Y(n5103) );
	nand4_1 U9567( .A(n10482), .B(n9350), .C(n9351), .D(n9352), .Y(n9349) );
	nor2_1 U9568( .A(n6360), .B(n9353), .Y(n9351) );
	a21oi_1 U9569( .A1(n10242), .A2(g35), .B1(n10263), .Y(n9353) );
	a21oi_1 U9570( .A1(n8593), .A2(n10482), .B1(n9354), .Y(n9348) );
	a21oi_1 U9571( .A1(n9352), .A2(n9350), .B1(n9355), .Y(n9354) );
	a21oi_1 U9572( .A1(n8964), .A2(n8412), .B1(n7313), .Y(n9355) );
	nor3_1 U9573( .A(n10242), .B(n10263), .C(n8593), .Y(n7313) );
	inv_1 U9574( .A(n10482), .Y(n8412) );
	nand2_1 U9575( .A(n10689), .B(n9356), .Y(n9350) );
	o21ai_0 U9576( .A1(n6248), .A2(n8042), .B1(n9357), .Y(n5102) );
	mux2i_1 U9577( .A0(n9358), .A1(n9359), .S(n8175), .Y(n9357) );
	nor2_1 U9578( .A(n6359), .B(n9360), .Y(n9359) );
	and2_0 U9579( .A(n9360), .B(n7513), .X(n9358) );
	inv_1 U9580( .A(n10565), .Y(n8042) );
	o22ai_1 U9581( .A1(n6205), .A2(n7076), .B1(n9361), .B2(n6296), .Y(n5101) );
	nor2_1 U9582( .A(n10591), .B(n9362), .Y(n9361) );
	o22ai_1 U9583( .A1(n6205), .A2(n9363), .B1(n9364), .B2(n8218), .Y(n5100) );
	xnor2_1 U9584( .A(n9365), .B(n9366), .Y(n9364) );
	inv_1 U9585( .A(n10601), .Y(n9363) );
	o211ai_1 U9586( .A1(n6203), .A2(n8060), .B1(n6400), .C1(n9367), .Y(n5099) );
	mux2i_1 U9587( .A0(n9368), .A1(n9369), .S(n7796), .Y(n9367) );
	inv_1 U9588( .A(n10435), .Y(n7796) );
	and2_0 U9589( .A(n6385), .B(n9370), .X(n9369) );
	nor2_1 U9590( .A(n9370), .B(n6301), .Y(n9368) );
	nor2_1 U9591( .A(n8061), .B(n8060), .Y(n9370) );
	inv_1 U9592( .A(n10424), .Y(n8060) );
	o32ai_1 U9593( .A1(n9371), .A2(n6348), .A3(n6934), .B1(n6201), .B2(n8361), .Y(n5098) );
	mux2i_1 U9594( .A0(n9372), .A1(n10188), .S(n8622), .Y(n9371) );
	a21oi_1 U9595( .A1(n8625), .A2(n8628), .B1(n8362), .Y(n9372) );
	and2_0 U9596( .A(n9373), .B(n7050), .X(n8362) );
	nor2_1 U9597( .A(n6360), .B(n8373), .Y(n5097) );
	inv_1 U9598( .A(g24265), .Y(n8373) );
	o22ai_1 U9599( .A1(n8302), .A2(n8526), .B1(n9010), .B2(n8960), .Y(n5096) );
	and2_0 U9600( .A(n6248), .B(n9374), .X(n9010) );
	nand3_1 U9601( .A(n8959), .B(n6376), .C(n9375), .Y(n9374) );
	inv_1 U9602( .A(n10300), .Y(n8526) );
	inv_1 U9603( .A(n6534), .Y(n8302) );
	nor2_1 U9604( .A(n8962), .B(n6367), .Y(n6534) );
	inv_1 U9605( .A(n8301), .Y(n8962) );
	nor2_1 U9606( .A(n6934), .B(n9375), .Y(n8301) );
	o21ai_0 U9607( .A1(n6237), .A2(n5863), .B1(n9376), .Y(n5095) );
	mux2_1 U9608( .A0(n6446), .A1(n6441), .S(n10697), .X(n9376) );
	or2_0 U9609( .A(n6314), .B(n7133), .X(n6441) );
	nand2_1 U9610( .A(n7133), .B(n6334), .Y(n6446) );
	nor3_1 U9611( .A(n8503), .B(n9377), .C(n5891), .Y(n7133) );
	o22ai_1 U9612( .A1(n6305), .A2(n9378), .B1(n6193), .B2(n8093), .Y(n5094) );
	o21ai_0 U9613( .A1(n6046), .A2(n8926), .B1(n9379), .Y(n5093) );
	mux2i_1 U9614( .A0(n9380), .A1(n9381), .S(n9382), .Y(n9379) );
	nor3_1 U9615( .A(n7803), .B(n10692), .C(n6306), .Y(n9381) );
	inv_1 U9616( .A(n8501), .Y(n7803) );
	nand2_1 U9617( .A(n6222), .B(n9383), .Y(n9380) );
	nand3_1 U9618( .A(n8501), .B(n6372), .C(n10692), .Y(n9383) );
	o22ai_1 U9619( .A1(n6205), .A2(n6694), .B1(n6301), .B2(n9384), .Y(n5092) );
	mux2i_1 U9620( .A0(n9385), .A1(n11917), .S(n7202), .Y(n9384) );
	nand2_1 U9621( .A(n10230), .B(n9386), .Y(n7202) );
	nand3_1 U9622( .A(n11916), .B(n9387), .C(n9388), .Y(n9386) );
	a21oi_1 U9623( .A1(n7199), .A2(n7200), .B1(n6695), .Y(n9385) );
	and2_0 U9624( .A(n7050), .B(n9389), .X(n6695) );
	and3_1 U9625( .A(n9390), .B(n6880), .C(n11769), .X(n7050) );
	nand2_1 U9626( .A(n11917), .B(n6694), .Y(n7200) );
	inv_1 U9627( .A(n8775), .Y(n7199) );
	nor2_1 U9628( .A(n6694), .B(n11917), .Y(n8775) );
	inv_1 U9629( .A(n10327), .Y(n6694) );
	o32ai_1 U9630( .A1(n9391), .A2(n6348), .A3(n6981), .B1(n6982), .B2(n8440), .Y(n5091) );
	inv_1 U9631( .A(n10478), .Y(n9391) );
	o21ai_0 U9632( .A1(n8636), .A2(n9392), .B1(n9393), .Y(n5090) );
	mux2i_1 U9633( .A0(n9394), .A1(n9395), .S(n8802), .Y(n9393) );
	inv_1 U9634( .A(n10644), .Y(n8802) );
	nor2_1 U9635( .A(n10504), .B(n8643), .Y(n9395) );
	nand2_1 U9636( .A(n6225), .B(n8803), .Y(n9394) );
	nand3_1 U9637( .A(n10504), .B(n6376), .C(n8642), .Y(n8803) );
	nor2_1 U9638( .A(n9396), .B(n6301), .Y(n5089) );
	and3_1 U9639( .A(n10297), .B(n7999), .C(g4467), .X(n9396) );
	o22ai_1 U9640( .A1(n6305), .A2(n6508), .B1(n6193), .B2(n9397), .Y(n5088) );
	inv_1 U9641( .A(n10660), .Y(n9397) );
	o221ai_1 U9642( .A1(n9398), .A2(n6309), .B1(n6217), .B2(n7449), .C1(n9399), .Y(n5087) );
	nand4_1 U9643( .A(n10483), .B(n9400), .C(n9401), .D(n9402), .Y(n9399) );
	nor2_1 U9644( .A(n6359), .B(n9403), .Y(n9401) );
	a21oi_1 U9645( .A1(n10243), .A2(g35), .B1(n10264), .Y(n9403) );
	a21oi_1 U9646( .A1(n9243), .A2(n10483), .B1(n9404), .Y(n9398) );
	a21oi_1 U9647( .A1(n9402), .A2(n9400), .B1(n9405), .Y(n9404) );
	a21oi_1 U9648( .A1(n9406), .A2(n7528), .B1(n7022), .Y(n9405) );
	nor3_1 U9649( .A(n10243), .B(n10264), .C(n9243), .Y(n7022) );
	inv_1 U9650( .A(n10483), .Y(n7528) );
	nand2_1 U9651( .A(n9407), .B(n6586), .Y(n9400) );
	nor2_1 U9652( .A(n6359), .B(n7206), .Y(n5086) );
	inv_1 U9653( .A(g25689), .Y(n7206) );
	o221ai_1 U9654( .A1(n6951), .A2(n8731), .B1(n6217), .B2(n8603), .C1(n8732), .Y(n5085) );
	nand3_1 U9655( .A(n7946), .B(n6376), .C(n10683), .Y(n8732) );
	inv_1 U9656( .A(n10683), .Y(n8603) );
	inv_1 U9657( .A(n10639), .Y(n8731) );
	or2_0 U9658( .A(n6314), .B(n7946), .X(n6951) );
	nor4_1 U9659( .A(n7474), .B(n9408), .C(n8536), .D(n8259), .Y(n7946) );
	o221ai_1 U9660( .A1(n9409), .A2(n6725), .B1(n6299), .B2(n9410), .C1(n9411), .Y(n5084) );
	nand3_1 U9661( .A(n6416), .B(n10536), .C(n9412), .Y(n9411) );
	mux2i_1 U9662( .A0(n10151), .A1(n10183), .S(n6725), .Y(n9412) );
	a21oi_1 U9663( .A1(n9413), .A2(n10151), .B1(n6437), .Y(n9409) );
	nor2_1 U9664( .A(n10536), .B(n6366), .Y(n9413) );
	o21ai_0 U9665( .A1(n6233), .A2(n8200), .B1(n9414), .Y(n5083) );
	mux2i_1 U9666( .A0(n9415), .A1(n9416), .S(n9417), .Y(n9414) );
	nor2_1 U9667( .A(n10567), .B(n6365), .Y(n9416) );
	nor2_1 U9668( .A(n7544), .B(n8037), .Y(n9415) );
	inv_1 U9669( .A(n10567), .Y(n8037) );
	o32ai_1 U9670( .A1(n9418), .A2(n6347), .A3(n6934), .B1(n6200), .B2(n8408), .Y(n5082) );
	mux2i_1 U9671( .A0(n9419), .A1(n10193), .S(n8902), .Y(n9418) );
	a21oi_1 U9672( .A1(n9420), .A2(n9421), .B1(n8409), .Y(n9419) );
	and2_0 U9673( .A(n9373), .B(n9175), .X(n8409) );
	o221ai_1 U9674( .A1(n6306), .A2(n9422), .B1(n6216), .B2(n6397), .C1(n6400), .Y(n5081) );
	nand2_1 U9675( .A(n6339), .B(n6398), .Y(n6400) );
	inv_1 U9676( .A(n10714), .Y(n6398) );
	nand2_1 U9677( .A(n9423), .B(n8061), .Y(n9422) );
	inv_1 U9678( .A(n8062), .Y(n8061) );
	nor2_1 U9679( .A(n9424), .B(n6638), .Y(n8062) );
	o21ai_0 U9680( .A1(n6395), .A2(n6397), .B1(n5882), .Y(n9423) );
	nand2_1 U9681( .A(n7635), .B(n10235), .Y(n6395) );
	nor2_1 U9682( .A(n6637), .B(n6638), .Y(n7635) );
	nand2_1 U9683( .A(n10338), .B(n8366), .Y(n6638) );
	nor2_1 U9684( .A(n8365), .B(n9425), .Y(n8366) );
	o32ai_1 U9685( .A1(n6311), .A2(n9426), .A3(n9427), .B1(n6200), .B2(n7348), .Y(n5080) );
	inv_1 U9686( .A(n10487), .Y(n7348) );
	a21oi_1 U9687( .A1(n7926), .A2(n8506), .B1(n10580), .Y(n9427) );
	nor4_1 U9688( .A(n10238), .B(n7833), .C(n7040), .D(n9428), .Y(n9426) );
	o32ai_1 U9689( .A1(n6311), .A2(n9429), .A3(n9430), .B1(n6200), .B2(n9431), .Y(n5079) );
	a21oi_1 U9690( .A1(n9432), .A2(n8726), .B1(n10908), .Y(n9430) );
	nor3_1 U9691( .A(n9433), .B(n7922), .C(n7472), .Y(n9429) );
	xnor2_1 U9692( .A(n10257), .B(n8698), .Y(n9433) );
	o32ai_1 U9693( .A1(n6312), .A2(n10418), .A3(n9434), .B1(n6199), .B2(n9135), .Y(n5078) );
	o32ai_1 U9694( .A1(n5970), .A2(n9435), .A3(n6312), .B1(n9436), .B2(n8518), .Y(n5077) );
	nor2_1 U9695( .A(n9437), .B(n6437), .Y(n9436) );
	nor4_1 U9696( .A(n11834), .B(n6368), .C(n8519), .D(n9438), .Y(n9437) );
	o21ai_0 U9697( .A1(n6233), .A2(n8029), .B1(n9439), .Y(n5076) );
	mux2i_1 U9698( .A0(n9440), .A1(n6257), .S(n9441), .Y(n9439) );
	nor2_1 U9699( .A(n7332), .B(n7506), .Y(n9441) );
	nand2_1 U9700( .A(n7410), .B(n7327), .Y(n7332) );
	inv_1 U9701( .A(n10202), .Y(n7410) );
	nor2_1 U9702( .A(n6281), .B(n5936), .Y(n9440) );
	inv_1 U9703( .A(n10748), .Y(n8029) );
	nor2_1 U9704( .A(n6359), .B(n9442), .Y(n5075) );
	o21ai_0 U9705( .A1(n6233), .A2(n5985), .B1(n9443), .Y(n5074) );
	mux2i_1 U9706( .A0(n9444), .A1(n6257), .S(n9445), .Y(n9443) );
	nor2_1 U9707( .A(n7875), .B(n6808), .Y(n9445) );
	nand2_1 U9708( .A(n11968), .B(n10275), .Y(n6808) );
	nor2_1 U9709( .A(n6281), .B(n9446), .Y(n9444) );
	o22ai_1 U9710( .A1(n6206), .A2(n9447), .B1(n9448), .B2(n6297), .Y(n5073) );
	nor2_1 U9711( .A(n9449), .B(n10429), .Y(n9448) );
	nor4_1 U9712( .A(g56), .B(g54), .C(g53), .D(n9450), .Y(n9449) );
	inv_1 U9713( .A(n10575), .Y(n9447) );
	o21ai_0 U9714( .A1(n6233), .A2(n9366), .B1(n9451), .Y(n5072) );
	mux2i_1 U9715( .A0(n9452), .A1(n9453), .S(n9454), .Y(n9451) );
	nor2_1 U9716( .A(n10290), .B(n8350), .Y(n9453) );
	nor2_1 U9717( .A(n9455), .B(n8218), .Y(n9452) );
	o22ai_1 U9718( .A1(n6206), .A2(n8818), .B1(n9456), .B2(n6646), .Y(n5071) );
	inv_1 U9719( .A(n6794), .Y(n6646) );
	nor2_1 U9720( .A(n7207), .B(n6300), .Y(n6794) );
	xnor2_1 U9721( .A(n10163), .B(n9120), .Y(n9456) );
	nor3_1 U9722( .A(n7667), .B(n10270), .C(n10153), .Y(n5070) );
	inv_1 U9723( .A(n7408), .Y(n7667) );
	a21oi_1 U9724( .A1(n9027), .A2(n8817), .B1(n6309), .Y(n7408) );
	o21ai_0 U9725( .A1(n6233), .A2(n9034), .B1(n9457), .Y(n5069) );
	mux2i_1 U9726( .A0(n9458), .A1(n9459), .S(n9460), .Y(n9457) );
	nor2_1 U9727( .A(n10561), .B(n6366), .Y(n9459) );
	nor2_1 U9728( .A(n6734), .B(n9461), .Y(n9458) );
	and2_0 U9729( .A(n6385), .B(g8475), .X(n5068) );
	nor3_1 U9730( .A(n6869), .B(n10274), .C(n10159), .Y(n5067) );
	inv_1 U9731( .A(n9462), .Y(n6869) );
	o221ai_1 U9732( .A1(n9071), .A2(n6030), .B1(n9463), .B2(n9464), .C1(n9465), .Y(n5066) );
	a22oi_1 U9733( .A1(n10545), .A2(n6747), .B1(n10333), .B2(n6437), .Y(n9465) );
	inv_1 U9734( .A(n8127), .Y(n9464) );
	a221oi_1 U9735( .A1(n10721), .A2(n7087), .B1(n8125), .B2(n11852), .C1(n9466), .Y(n9463) );
	o32ai_1 U9736( .A1(n7086), .A2(n11877), .A3(n10333), .B1(n10172), .B2(n9467), .Y(n9466) );
	a22oi_1 U9737( .A1(n11784), .A2(n10333), .B1(n11825), .B2(n11877), .Y(n9467) );
	inv_1 U9738( .A(n10488), .Y(n7086) );
	nand2_1 U9739( .A(n9247), .B(n6334), .Y(n9071) );
	nor3_1 U9740( .A(n6745), .B(n6742), .C(n5892), .Y(n9247) );
	inv_1 U9741( .A(n10333), .Y(n6745) );
	o21ai_0 U9742( .A1(n6233), .A2(n9468), .B1(n9469), .Y(n5065) );
	mux2i_1 U9743( .A0(n9470), .A1(n9471), .S(n9431), .Y(n9469) );
	nor2_1 U9744( .A(n6359), .B(n9472), .Y(n9471) );
	and2_0 U9745( .A(n9472), .B(n6344), .X(n9470) );
	nand3_1 U9746( .A(n8568), .B(n8974), .C(n10906), .Y(n9472) );
	nor3_1 U9747( .A(n7922), .B(n10440), .C(n6801), .Y(n8568) );
	inv_1 U9748( .A(n10906), .Y(n9468) );
	o221ai_1 U9749( .A1(n9230), .A2(n8735), .B1(n6217), .B2(n5881), .C1(n9473), .Y(n5064) );
	nand3_1 U9750( .A(n6340), .B(n8738), .C(n9474), .Y(n9473) );
	nand2_1 U9751( .A(n9008), .B(n8909), .Y(n8738) );
	inv_1 U9752( .A(n8885), .Y(n8909) );
	nand2_1 U9753( .A(n8431), .B(n6334), .Y(n8735) );
	inv_1 U9754( .A(n10287), .Y(n9230) );
	o21ai_0 U9755( .A1(n6233), .A2(n6044), .B1(n9475), .Y(n5063) );
	mux2i_1 U9756( .A0(n9476), .A1(n9281), .S(n10502), .Y(n9475) );
	inv_1 U9757( .A(n9477), .Y(n9281) );
	nor2_1 U9758( .A(n6281), .B(n9478), .Y(n9476) );
	o22ai_1 U9759( .A1(n6207), .A2(n9479), .B1(n9480), .B2(n6298), .Y(n5062) );
	nor3_1 U9760( .A(n9481), .B(n10216), .C(n9362), .Y(n9480) );
	o21ai_0 U9761( .A1(n6233), .A2(n9482), .B1(n9483), .Y(n5061) );
	mux2i_1 U9762( .A0(n9484), .A1(n6257), .S(n9485), .Y(n9483) );
	nor2_1 U9763( .A(n7731), .B(n8266), .Y(n9485) );
	nand2_1 U9764( .A(n10272), .B(n5902), .Y(n7731) );
	nor2_1 U9765( .A(n6281), .B(n9486), .Y(n9484) );
	o21ai_0 U9766( .A1(n6233), .A2(n7881), .B1(n9487), .Y(n5060) );
	mux2i_1 U9767( .A0(n9488), .A1(n6257), .S(n9489), .Y(n9487) );
	nor2_1 U9768( .A(n6627), .B(n8191), .Y(n9489) );
	nor2_1 U9769( .A(n6280), .B(n5927), .Y(n9488) );
	o32ai_1 U9770( .A1(n6312), .A2(g9680), .A3(n9490), .B1(n6200), .B2(n9491), .Y(n5059) );
	a21oi_1 U9771( .A1(g9617), .A2(n9491), .B1(n10609), .Y(n9490) );
	inv_1 U9772( .A(n10608), .Y(n9491) );
	o21ai_0 U9773( .A1(n6233), .A2(n9492), .B1(n7544), .Y(n5058) );
	o32ai_1 U9774( .A1(n8687), .A2(n10155), .A3(n7026), .B1(n6199), .B2(n5902), .Y(n5057) );
	inv_1 U9775( .A(n9493), .Y(n8687) );
	o21ai_0 U9776( .A1(n6234), .A2(n9494), .B1(n9495), .Y(n5056) );
	mux2i_1 U9777( .A0(n9496), .A1(n6257), .S(n9497), .Y(n9495) );
	nor2_1 U9778( .A(n6668), .B(n8023), .Y(n9497) );
	nand2_1 U9779( .A(n10273), .B(n5899), .Y(n8023) );
	nor2_1 U9780( .A(n6280), .B(n6664), .Y(n9496) );
	inv_1 U9781( .A(n10781), .Y(n6664) );
	o21ai_0 U9782( .A1(n6234), .A2(n7782), .B1(n9498), .Y(n5055) );
	mux2i_1 U9783( .A0(n9499), .A1(n6257), .S(n9500), .Y(n9498) );
	nor2_1 U9784( .A(n6789), .B(n7178), .Y(n9500) );
	nand3_1 U9785( .A(n6865), .B(n5903), .C(n8614), .Y(n6789) );
	inv_1 U9786( .A(n10274), .Y(n6865) );
	nor2_1 U9787( .A(n6280), .B(n9501), .Y(n9499) );
	inv_1 U9788( .A(n10795), .Y(n7782) );
	o32ai_1 U9789( .A1(n6058), .A2(n6347), .A3(n8160), .B1(n8273), .B2(n9502), .Y(n5054) );
	o221ai_1 U9790( .A1(n5892), .A2(n8474), .B1(n6218), .B2(n9314), .C1(n9503), .Y(n5053) );
	a21oi_1 U9791( .A1(n9504), .A2(n8127), .B1(n8840), .Y(n9503) );
	nor2_1 U9792( .A(n6742), .B(n6299), .Y(n8127) );
	nor2_1 U9793( .A(n10333), .B(n8125), .Y(n9504) );
	nor2_1 U9794( .A(n6741), .B(n11877), .Y(n8125) );
	inv_1 U9795( .A(n10581), .Y(n9314) );
	o21ai_0 U9796( .A1(n6234), .A2(n7270), .B1(n9505), .Y(n5052) );
	mux2i_1 U9797( .A0(n9506), .A1(n9507), .S(n10514), .Y(n9505) );
	nor3_1 U9798( .A(n6727), .B(n8811), .C(n8813), .Y(n9507) );
	inv_1 U9799( .A(n6416), .Y(n6727) );
	nor3_1 U9800( .A(n7515), .B(n8812), .C(n6307), .Y(n6416) );
	and4_1 U9801( .A(n9508), .B(n10177), .C(n10151), .D(n6414), .X(n7515) );
	mux2i_1 U9802( .A0(n6410), .A1(n6773), .S(g84), .Y(n9508) );
	inv_1 U9803( .A(n10360), .Y(n6773) );
	inv_1 U9804( .A(n10359), .Y(n6410) );
	o22ai_1 U9805( .A1(n6305), .A2(n7265), .B1(n6347), .B2(n9509), .Y(n9506) );
	inv_1 U9806( .A(n8811), .Y(n9509) );
	nor2_1 U9807( .A(n7270), .B(n7271), .Y(n8811) );
	inv_1 U9808( .A(n7273), .Y(n7271) );
	nor3_1 U9809( .A(n6725), .B(n9510), .C(n7266), .Y(n7273) );
	inv_1 U9810( .A(n10536), .Y(n7266) );
	inv_1 U9811( .A(n10298), .Y(n6725) );
	inv_1 U9812( .A(n8813), .Y(n7265) );
	nor2_1 U9813( .A(n9410), .B(n10558), .Y(n8813) );
	inv_1 U9814( .A(n7272), .Y(n9410) );
	nor3_1 U9815( .A(n10298), .B(n10536), .C(n6721), .Y(n7272) );
	inv_1 U9816( .A(n10183), .Y(n6721) );
	inv_1 U9817( .A(n10558), .Y(n7270) );
	o22ai_1 U9818( .A1(n9209), .A2(n8660), .B1(n9511), .B2(n7228), .Y(n5051) );
	a21oi_1 U9819( .A1(n9493), .A2(n9209), .B1(n6437), .Y(n9511) );
	nor2_1 U9820( .A(n8690), .B(n6367), .Y(n9493) );
	or3_1 U9821( .A(n8690), .B(n10155), .C(n6308), .X(n8660) );
	nor3_1 U9822( .A(n9322), .B(n10163), .C(n9512), .Y(n8690) );
	nand3_1 U9823( .A(n6760), .B(n9513), .C(n9514), .Y(n5050) );
	nand2_1 U9824( .A(g4501), .B(n6763), .Y(n9514) );
	o22ai_1 U9825( .A1(n6305), .A2(n9515), .B1(n6193), .B2(n5967), .Y(n5049) );
	o21ai_0 U9826( .A1(n6234), .A2(n6092), .B1(n9516), .Y(n5048) );
	a22oi_1 U9827( .A1(n10458), .A2(n7369), .B1(g14189), .B2(n7370), .Y(n9516) );
	nor2_1 U9828( .A(n6358), .B(n9517), .Y(n5047) );
	o21ai_0 U9829( .A1(n6234), .A2(n5922), .B1(n9518), .Y(n5046) );
	mux2i_1 U9830( .A0(n9519), .A1(n6257), .S(n9520), .Y(n9518) );
	nor2_1 U9831( .A(n6899), .B(n6971), .Y(n9520) );
	nand2_1 U9832( .A(n11942), .B(n10270), .Y(n6971) );
	inv_1 U9833( .A(n7668), .Y(n6899) );
	nor2_1 U9834( .A(n7327), .B(n10202), .Y(n7668) );
	nor2_1 U9835( .A(n6280), .B(n7846), .Y(n9519) );
	inv_1 U9836( .A(n10744), .Y(n7846) );
	and2_0 U9837( .A(n6384), .B(g9682), .X(n5045) );
	o21ai_0 U9838( .A1(n6234), .A2(n6610), .B1(n9521), .Y(n5044) );
	mux2i_1 U9839( .A0(n9522), .A1(n9523), .S(n6823), .Y(n9521) );
	nor2_1 U9840( .A(n6358), .B(n9524), .Y(n9523) );
	and2_0 U9841( .A(n9524), .B(n6344), .X(n9522) );
	o221ai_1 U9842( .A1(n9525), .A2(n6308), .B1(n6218), .B2(n7460), .C1(n9526), .Y(n5043) );
	nand4_1 U9843( .A(n10480), .B(n9527), .C(n9528), .D(n9529), .Y(n9526) );
	nor2_1 U9844( .A(n6358), .B(n9530), .Y(n9528) );
	a21oi_1 U9845( .A1(n10240), .A2(g35), .B1(n10261), .Y(n9530) );
	inv_1 U9846( .A(n10261), .Y(n7460) );
	a21oi_1 U9847( .A1(n10480), .A2(n7433), .B1(n9531), .Y(n9525) );
	a21oi_1 U9848( .A1(n9529), .A2(n9527), .B1(n9532), .Y(n9531) );
	a21oi_1 U9849( .A1(n9533), .A2(n7756), .B1(n7566), .Y(n9532) );
	nor3_1 U9850( .A(n10240), .B(n10261), .C(n7433), .Y(n7566) );
	inv_1 U9851( .A(n10480), .Y(n7756) );
	or2_0 U9852( .A(n9534), .B(n9535), .X(n9527) );
	nor2_1 U9853( .A(n6353), .B(n9536), .Y(n5042) );
	o21ai_0 U9854( .A1(n6234), .A2(n7148), .B1(n9537), .Y(n5041) );
	mux2i_1 U9855( .A0(n9538), .A1(n6257), .S(n9539), .Y(n9537) );
	nor2_1 U9856( .A(n6570), .B(n8483), .Y(n9539) );
	nand2_1 U9857( .A(n9202), .B(n6566), .Y(n6570) );
	nor2_1 U9858( .A(n6280), .B(n5935), .Y(n9538) );
	inv_1 U9859( .A(n10839), .Y(n7148) );
	o21ai_0 U9860( .A1(n6234), .A2(n9540), .B1(n9541), .Y(n5040) );
	mux2i_1 U9861( .A0(n9542), .A1(n9543), .S(n9544), .Y(n9541) );
	nor2_1 U9862( .A(n6279), .B(n9545), .Y(n9543) );
	nor2_1 U9863( .A(n10304), .B(n8520), .Y(n9542) );
	o32ai_1 U9864( .A1(n6311), .A2(g9497), .A3(n9546), .B1(n6199), .B2(n9547), .Y(n5039) );
	a21oi_1 U9865( .A1(g9553), .A2(n9547), .B1(n10183), .Y(n9546) );
	inv_1 U9866( .A(n10613), .Y(n9547) );
	o22ai_1 U9867( .A1(n6207), .A2(n9548), .B1(n9549), .B2(n6298), .Y(n5038) );
	nor3_1 U9868( .A(n9550), .B(n10451), .C(n9551), .Y(n9549) );
	o22ai_1 U9869( .A1(n6207), .A2(n7736), .B1(n6277), .B2(n9552), .Y(n5037) );
	mux2i_1 U9870( .A0(n9553), .A1(n9554), .S(n7556), .Y(n9552) );
	inv_1 U9871( .A(n10446), .Y(n7556) );
	nor2_1 U9872( .A(n10405), .B(n9553), .Y(n9554) );
	o21ai_0 U9873( .A1(n6234), .A2(n9555), .B1(n9556), .Y(n5036) );
	a22oi_1 U9874( .A1(n10218), .A2(n7369), .B1(g14125), .B2(n7370), .Y(n9556) );
	inv_1 U9875( .A(n10302), .Y(n9555) );
	o21ai_0 U9876( .A1(n8841), .A2(n9557), .B1(n9558), .Y(n5035) );
	mux2i_1 U9877( .A0(n9559), .A1(n9560), .S(n8935), .Y(n9558) );
	inv_1 U9878( .A(n10641), .Y(n8935) );
	nor2_1 U9879( .A(n10503), .B(n8848), .Y(n9560) );
	nand2_1 U9880( .A(n6224), .B(n8936), .Y(n9559) );
	nand3_1 U9881( .A(n10503), .B(n6377), .C(n8847), .Y(n8936) );
	o21ai_0 U9882( .A1(n6234), .A2(n8759), .B1(n9561), .Y(n5034) );
	mux2i_1 U9883( .A0(n9562), .A1(n9563), .S(n7725), .Y(n9561) );
	nor2_1 U9884( .A(n6351), .B(n9564), .Y(n9563) );
	nor2_1 U9885( .A(n9565), .B(n8486), .Y(n9562) );
	inv_1 U9886( .A(n9564), .Y(n9565) );
	inv_1 U9887( .A(n10408), .Y(n8759) );
	o22ai_1 U9888( .A1(n6208), .A2(n9566), .B1(n9567), .B2(n8467), .Y(n5033) );
	xnor2_1 U9889( .A(n9568), .B(n9569), .Y(n9567) );
	o32ai_1 U9890( .A1(n6059), .A2(n6347), .A3(n8383), .B1(n8673), .B2(n9570), .Y(n5032) );
	nor2_1 U9891( .A(n6352), .B(n9571), .Y(n5031) );
	o21ai_0 U9892( .A1(n6234), .A2(n8525), .B1(n9572), .Y(n5030) );
	nand3_1 U9893( .A(n8959), .B(n9573), .C(n9574), .Y(n9572) );
	o32ai_1 U9894( .A1(n9575), .A2(n9576), .A3(n6530), .B1(n6302), .B2(n7414), .Y(n9574) );
	inv_1 U9895( .A(n8203), .Y(n6530) );
	nor2_1 U9896( .A(n9577), .B(n6299), .Y(n8203) );
	inv_1 U9897( .A(n9578), .Y(n9576) );
	nand3_1 U9898( .A(n9579), .B(n9375), .C(n10371), .Y(n9573) );
	inv_1 U9899( .A(n7416), .Y(n8959) );
	o221ai_1 U9900( .A1(n9580), .A2(n6308), .B1(n6218), .B2(n9322), .C1(n8232), .Y(n5029) );
	xnor2_1 U9901( .A(n10288), .B(n9581), .Y(n9580) );
	inv_1 U9902( .A(n9582), .Y(n5028) );
	a21oi_1 U9903( .A1(n6437), .A2(g20049), .B1(n37), .Y(n9582) );
	inv_1 U9904( .A(n9583), .Y(n5027) );
	a22oi_1 U9905( .A1(n6437), .A2(n11892), .B1(n9584), .B2(n6337), .Y(n9583) );
	a21oi_1 U9906( .A1(n6197), .A2(n9585), .B1(n5916), .Y(n5026) );
	or2_0 U9907( .A(n9434), .B(n6369), .X(n9585) );
	nor2_1 U9908( .A(n9586), .B(n9135), .Y(n9434) );
	o21ai_0 U9909( .A1(n6234), .A2(n9587), .B1(n9588), .Y(n5025) );
	a22oi_1 U9910( .A1(n10178), .A2(n7369), .B1(g14167), .B2(n7370), .Y(n9588) );
	nor4_1 U9911( .A(n8489), .B(n6302), .C(n10219), .D(n10406), .Y(n7370) );
	and2_0 U9912( .A(n6345), .B(n9589), .X(n7369) );
	or3_1 U9913( .A(n10219), .B(n10406), .C(n8489), .X(n9589) );
	inv_1 U9914( .A(n10187), .Y(n9587) );
	o21ai_0 U9915( .A1(n6234), .A2(n6002), .B1(n9590), .Y(n5024) );
	mux2i_1 U9916( .A0(n9591), .A1(n6257), .S(n9592), .Y(n9590) );
	nor2_1 U9917( .A(n7669), .B(n7506), .Y(n9592) );
	nand2_1 U9918( .A(n10202), .B(n7327), .Y(n7669) );
	nor2_1 U9919( .A(n6279), .B(n6003), .Y(n9591) );
	o21ai_0 U9920( .A1(n6234), .A2(n9593), .B1(n8300), .Y(n5023) );
	o221ai_1 U9921( .A1(n9594), .A2(n5964), .B1(n10292), .B2(n6708), .C1(n9595), .Y(n5022) );
	mux2i_1 U9922( .A0(n9596), .A1(n9597), .S(n6707), .Y(n9595) );
	nor4_1 U9923( .A(n9377), .B(n8503), .C(n9598), .D(n6744), .Y(n9597) );
	inv_1 U9924( .A(n10292), .Y(n8503) );
	nand2_1 U9925( .A(n6222), .B(n6708), .Y(n9596) );
	inv_1 U9926( .A(n7716), .Y(n6708) );
	nor3_1 U9927( .A(n7657), .B(n9377), .C(n9598), .Y(n7716) );
	a211oi_1 U9928( .A1(n6329), .A2(n9598), .B1(n6746), .C1(n7661), .Y(n9594) );
	nor2_1 U9929( .A(n6279), .B(n6709), .Y(n7661) );
	inv_1 U9930( .A(n9377), .Y(n6709) );
	o221ai_1 U9931( .A1(n8036), .A2(n8549), .B1(n6220), .B2(n9016), .C1(n8550), .Y(n5021) );
	nand3_1 U9932( .A(n8824), .B(n6377), .C(n10505), .Y(n8550) );
	inv_1 U9933( .A(n9599), .Y(n8824) );
	inv_1 U9934( .A(n10505), .Y(n9016) );
	inv_1 U9935( .A(n10645), .Y(n8549) );
	nand2_1 U9936( .A(n6338), .B(n9599), .Y(n8036) );
	nand4_1 U9937( .A(g16656), .B(n9064), .C(n10378), .D(n9173), .Y(n9599) );
	o21ai_0 U9938( .A1(n6234), .A2(n9600), .B1(n9601), .Y(n5020) );
	mux2i_1 U9939( .A0(n9602), .A1(n6257), .S(n9603), .Y(n9601) );
	nor2_1 U9940( .A(n6681), .B(n8074), .Y(n9603) );
	nor2_1 U9941( .A(n6278), .B(n9292), .Y(n9602) );
	inv_1 U9942( .A(n10814), .Y(n9292) );
	o21ai_0 U9943( .A1(n6234), .A2(n8372), .B1(n9604), .Y(n5019) );
	mux2i_1 U9944( .A0(n9605), .A1(n9606), .S(n9607), .Y(n9604) );
	nor2_1 U9945( .A(n6351), .B(n9608), .Y(n9606) );
	nor2_1 U9946( .A(n9609), .B(n7108), .Y(n9605) );
	inv_1 U9947( .A(n9608), .Y(n9609) );
	nand2_1 U9948( .A(n10307), .B(n8371), .Y(n9608) );
	and2_0 U9949( .A(n9610), .B(n10383), .X(n8371) );
	o21ai_0 U9950( .A1(n6234), .A2(n6629), .B1(n9611), .Y(n5018) );
	mux2i_1 U9951( .A0(n9612), .A1(n6258), .S(n9613), .Y(n9611) );
	nor2_1 U9952( .A(n6627), .B(n8169), .Y(n9613) );
	nand2_1 U9953( .A(n8166), .B(n9046), .Y(n6627) );
	nor2_1 U9954( .A(n6279), .B(n9254), .Y(n9612) );
	inv_1 U9955( .A(n10763), .Y(n9254) );
	o21ai_0 U9956( .A1(n6235), .A2(n5986), .B1(n9614), .Y(n5017) );
	mux2i_1 U9957( .A0(n9615), .A1(n6258), .S(n9616), .Y(n9614) );
	nor2_1 U9958( .A(n8069), .B(n7026), .Y(n9616) );
	nand2_1 U9959( .A(n11956), .B(n10272), .Y(n7026) );
	nor2_1 U9960( .A(n6279), .B(n9617), .Y(n9615) );
	o21ai_0 U9961( .A1(n6235), .A2(n9618), .B1(n9619), .Y(n5016) );
	mux2i_1 U9962( .A0(n9620), .A1(n6258), .S(n9621), .Y(n9619) );
	nor2_1 U9963( .A(n7903), .B(n8250), .Y(n9621) );
	nor2_1 U9964( .A(n6279), .B(n8942), .Y(n9620) );
	inv_1 U9965( .A(n10788), .Y(n8942) );
	o21ai_0 U9966( .A1(n7396), .A2(n6089), .B1(n9622), .Y(n5015) );
	mux2i_1 U9967( .A0(n9623), .A1(n9624), .S(n7397), .Y(n9622) );
	inv_1 U9968( .A(n10647), .Y(n7397) );
	nor3_1 U9969( .A(n8604), .B(n11878), .C(n6307), .Y(n9624) );
	inv_1 U9970( .A(n6690), .Y(n8604) );
	nand2_1 U9971( .A(n6223), .B(n9625), .Y(n9623) );
	nand3_1 U9972( .A(n6690), .B(n6376), .C(n11878), .Y(n9625) );
	nand2_1 U9973( .A(n7395), .B(n6379), .Y(n7396) );
	nor2_1 U9974( .A(n6934), .B(n6690), .Y(n7395) );
	o21ai_0 U9975( .A1(n6235), .A2(n9626), .B1(n9627), .Y(n5014) );
	mux2i_1 U9976( .A0(n9628), .A1(n9629), .S(n9630), .Y(n9627) );
	nor2_1 U9977( .A(n10399), .B(n6367), .Y(n9629) );
	nor2_1 U9978( .A(n9631), .B(n8048), .Y(n9628) );
	and2_0 U9979( .A(n6385), .B(g10122), .X(n5013) );
	o21ai_0 U9980( .A1(n6235), .A2(n9632), .B1(n9633), .Y(n5012) );
	a22oi_1 U9981( .A1(n10187), .A2(n7746), .B1(n11763), .B2(n8289), .Y(n9633) );
	o22ai_1 U9982( .A1(n6208), .A2(n9634), .B1(n9635), .B2(n6296), .Y(n5011) );
	nor2_1 U9983( .A(g1277), .B(n10454), .Y(n9635) );
	inv_1 U9984( .A(n10590), .Y(n9634) );
	o21ai_0 U9985( .A1(n6047), .A2(n7605), .B1(n9636), .Y(n5010) );
	mux2i_1 U9986( .A0(n9637), .A1(n9638), .S(n7606), .Y(n9636) );
	inv_1 U9987( .A(n10627), .Y(n7606) );
	nor3_1 U9988( .A(n7005), .B(n10694), .C(n6306), .Y(n9638) );
	inv_1 U9989( .A(n6584), .Y(n7005) );
	nand2_1 U9990( .A(n6223), .B(n9639), .Y(n9637) );
	nand3_1 U9991( .A(n6584), .B(n6377), .C(n10694), .Y(n9639) );
	o21ai_0 U9992( .A1(n6235), .A2(n7017), .B1(n9640), .Y(n5009) );
	mux2i_1 U9993( .A0(n9641), .A1(n6258), .S(n9642), .Y(n9640) );
	nor2_1 U9994( .A(n7015), .B(n8941), .Y(n9642) );
	nor2_1 U9995( .A(n6279), .B(n7747), .Y(n9641) );
	and2_0 U9996( .A(n6385), .B(g8839), .X(n5008) );
	o221ai_1 U9997( .A1(n9643), .A2(n9644), .B1(n6220), .B2(n9645), .C1(n9646), .Y(n5007) );
	nand3_1 U9998( .A(n6340), .B(n9647), .C(n11837), .Y(n9646) );
	o21ai_0 U9999( .A1(n6917), .A2(n8460), .B1(n6919), .Y(n9644) );
	inv_1 U10000( .A(n9648), .Y(n6919) );
	inv_1 U10001( .A(n10846), .Y(n8460) );
	o21ai_0 U10002( .A1(n6235), .A2(n9461), .B1(n9649), .Y(n5006) );
	mux2i_1 U10003( .A0(n9650), .A1(n9651), .S(n9113), .Y(n9649) );
	and2_0 U10004( .A(n10561), .B(n9460), .X(n9113) );
	nor2_1 U10005( .A(n9034), .B(n9035), .Y(n9460) );
	nand2_1 U10006( .A(n10564), .B(n6733), .Y(n9035) );
	and3_1 U10007( .A(n7727), .B(n11954), .C(n9652), .X(n6733) );
	inv_1 U10008( .A(n10563), .Y(n9034) );
	nor2_1 U10009( .A(n10539), .B(n6367), .Y(n9651) );
	nor2_1 U10010( .A(n6734), .B(n9108), .Y(n9650) );
	inv_1 U10011( .A(n10539), .Y(n9108) );
	nand2_1 U10012( .A(n9652), .B(n6334), .Y(n6734) );
	and3_1 U10013( .A(n9653), .B(n9654), .C(n10267), .X(n9652) );
	o21ai_0 U10014( .A1(n10433), .A2(n8706), .B1(n7727), .Y(n9653) );
	inv_1 U10015( .A(n9655), .Y(n7727) );
	inv_1 U10016( .A(n10561), .Y(n9461) );
	o21ai_0 U10017( .A1(n7128), .A2(n6248), .B1(n9656), .Y(n5005) );
	mux2i_1 U10018( .A0(n9657), .A1(n9658), .S(n6439), .Y(n9656) );
	o21ai_0 U10019( .A1(n10559), .A2(n6438), .B1(n7131), .Y(n6439) );
	inv_1 U10020( .A(n7129), .Y(n7131) );
	o21ai_0 U10021( .A1(n11829), .A2(n6438), .B1(n9050), .Y(n7129) );
	a21oi_1 U10022( .A1(n7401), .A2(n6440), .B1(n7402), .Y(n9050) );
	inv_1 U10023( .A(n10386), .Y(n7401) );
	nor2_1 U10024( .A(n6279), .B(n6435), .Y(n9658) );
	nor2_1 U10025( .A(n10303), .B(n7130), .Y(n9657) );
	nand2_1 U10026( .A(n6440), .B(n6335), .Y(n7130) );
	inv_1 U10027( .A(n6438), .Y(n6440) );
	nand3_1 U10028( .A(n7790), .B(n6713), .C(n9659), .Y(n6438) );
	mux2i_1 U10029( .A0(n9660), .A1(n9661), .S(n6711), .Y(n9659) );
	and2_0 U10030( .A(n7787), .B(n7791), .X(n9660) );
	nor2_1 U10031( .A(n5934), .B(n6435), .Y(n7791) );
	inv_1 U10032( .A(n10303), .Y(n6435) );
	inv_1 U10033( .A(n10556), .Y(n6713) );
	nand2_1 U10034( .A(n11891), .B(n9661), .Y(n7790) );
	inv_1 U10035( .A(n10559), .Y(n7128) );
	o21ai_0 U10036( .A1(n6235), .A2(n6859), .B1(n9662), .Y(n5004) );
	mux2i_1 U10037( .A0(n9663), .A1(n6258), .S(n8170), .Y(n9662) );
	nor2_1 U10038( .A(n8169), .B(n6858), .Y(n8170) );
	nor2_1 U10039( .A(n6279), .B(n8078), .Y(n9663) );
	inv_1 U10040( .A(n10764), .Y(n6859) );
	o211ai_1 U10041( .A1(n9664), .A2(n8530), .B1(n9665), .C1(n8144), .Y(n5003) );
	nand3_1 U10042( .A(n11910), .B(n8528), .C(n8146), .Y(n9665) );
	inv_1 U10043( .A(n10934), .Y(n8530) );
	a21oi_1 U10044( .A1(n8532), .A2(n8147), .B1(n6437), .Y(n9664) );
	o21ai_0 U10045( .A1(n6235), .A2(n9158), .B1(n9666), .Y(n5002) );
	mux2i_1 U10046( .A0(n9667), .A1(n6258), .S(n9668), .Y(n9666) );
	nor2_1 U10047( .A(n6681), .B(n6995), .Y(n9668) );
	inv_1 U10048( .A(n9024), .Y(n6995) );
	nor2_1 U10049( .A(n9600), .B(n10208), .Y(n9024) );
	nor2_1 U10050( .A(n6280), .B(n7947), .Y(n9667) );
	inv_1 U10051( .A(n10804), .Y(n7947) );
	o22ai_1 U10052( .A1(n6305), .A2(n5906), .B1(n6193), .B2(n7404), .Y(n5001) );
	o21ai_0 U10053( .A1(n8273), .A2(n9669), .B1(n9670), .Y(n5000) );
	mux2i_1 U10054( .A0(n9671), .A1(n9672), .S(n9502), .Y(n9670) );
	inv_1 U10055( .A(n10650), .Y(n9502) );
	nor3_1 U10056( .A(n8274), .B(n11880), .C(n6307), .Y(n9672) );
	inv_1 U10057( .A(n6427), .Y(n8274) );
	nand2_1 U10058( .A(n6223), .B(n9673), .Y(n9671) );
	nand3_1 U10059( .A(n6427), .B(n6377), .C(n11880), .Y(n9673) );
	inv_1 U10060( .A(n10610), .Y(n9669) );
	nand2_1 U10061( .A(n8160), .B(n6379), .Y(n8273) );
	nor2_1 U10062( .A(n6934), .B(n6427), .Y(n8160) );
	o21ai_0 U10063( .A1(n6235), .A2(n9674), .B1(n9675), .Y(n50) );
	a22oi_1 U10064( .A1(n11766), .A2(n8051), .B1(n8056), .B2(n8799), .Y(n9675) );
	nand2_1 U10065( .A(n9676), .B(n9677), .Y(n8799) );
	mux2i_1 U10066( .A0(n9678), .A1(n9679), .S(n9680), .Y(n9677) );
	xnor2_1 U10067( .A(n7474), .B(g12470), .Y(n9680) );
	nand3_1 U10068( .A(n9681), .B(n9682), .C(n9683), .Y(n9679) );
	nand3_1 U10069( .A(g17688), .B(n10493), .C(n9684), .Y(n9683) );
	nand3_1 U10070( .A(n9685), .B(g17778), .C(n11841), .Y(n9682) );
	nand3_1 U10071( .A(n9686), .B(g14828), .C(n11827), .Y(n9681) );
	nand3_1 U10072( .A(n9687), .B(n9688), .C(n9689), .Y(n9678) );
	nand3_1 U10073( .A(g17778), .B(n8801), .C(n11870), .Y(n9689) );
	nand3_1 U10074( .A(g17688), .B(n10751), .C(n9686), .Y(n9688) );
	nand3_1 U10075( .A(n9684), .B(g14828), .C(n11871), .Y(n9687) );
	mux2_1 U10076( .A0(n9690), .A1(n9691), .S(n7474), .X(n9676) );
	a221oi_1 U10077( .A1(n9684), .A2(n9692), .B1(n8801), .B2(n9693), .C1(n9694), .Y(n9691) );
	o32ai_1 U10078( .A1(n9695), .A2(n5922), .A3(n8535), .B1(n9696), .B2(n8261), .Y(n9694) );
	a22oi_1 U10079( .A1(n10743), .A2(g17722), .B1(g17764), .B2(n10744), .Y( n9696) );
	inv_1 U10080( .A(n9686), .Y(n8535) );
	o22ai_1 U10081( .A1(n6900), .A2(n9697), .B1(n7354), .B2(n9698), .Y(n9693) );
	inv_1 U10082( .A(n10741), .Y(n7354) );
	inv_1 U10083( .A(n10742), .Y(n6900) );
	o22ai_1 U10084( .A1(n7349), .A2(n9699), .B1(n6894), .B2(n9700), .Y(n9692) );
	inv_1 U10085( .A(n10739), .Y(n6894) );
	inv_1 U10086( .A(n10740), .Y(n7349) );
	inv_1 U10087( .A(n8260), .Y(n9684) );
	a221oi_1 U10088( .A1(n9686), .A2(n9701), .B1(n8801), .B2(n9702), .C1(n9703), .Y(n9690) );
	o32ai_1 U10089( .A1(n5936), .A2(n8260), .A3(n9695), .B1(n9704), .B2(n8261), .Y(n9703) );
	inv_1 U10090( .A(n9685), .Y(n8261) );
	nor2_1 U10091( .A(n8053), .B(n10191), .Y(n9685) );
	a22oi_1 U10092( .A1(n10747), .A2(g12470), .B1(g17871), .B2(n10748), .Y( n9704) );
	nand2_1 U10093( .A(n10191), .B(n8053), .Y(n8260) );
	inv_1 U10094( .A(n10365), .Y(n8053) );
	o22ai_1 U10095( .A1(n7850), .A2(n7989), .B1(n9674), .B2(n9408), .Y(n9702) );
	inv_1 U10096( .A(n10746), .Y(n7989) );
	inv_1 U10097( .A(g17764), .Y(n7850) );
	inv_1 U10098( .A(n8536), .Y(n8801) );
	o22ai_1 U10099( .A1(n7804), .A2(n9699), .B1(n7333), .B2(n9700), .Y(n9701) );
	inv_1 U10100( .A(n10749), .Y(n7333) );
	inv_1 U10101( .A(n10750), .Y(n7804) );
	nor2_1 U10102( .A(n10365), .B(n10191), .Y(n9686) );
	nor2_1 U10103( .A(n8259), .B(n6300), .Y(n8056) );
	nor2_1 U10104( .A(n6280), .B(n9705), .Y(n8051) );
	inv_1 U10105( .A(n8259), .Y(n9705) );
	o21ai_0 U10106( .A1(n9706), .A2(n9707), .B1(n11906), .Y(n8259) );
	nand2_1 U10107( .A(n11910), .B(n9708), .Y(n9707) );
	inv_1 U10108( .A(n10745), .Y(n9674) );
	o21ai_0 U10109( .A1(n6235), .A2(n8649), .B1(n9709), .Y(n4999) );
	mux2i_1 U10110( .A0(n9710), .A1(n6258), .S(n9711), .Y(n9709) );
	nor2_1 U10111( .A(n7071), .B(n7016), .Y(n9711) );
	nor2_1 U10112( .A(n6280), .B(n8937), .Y(n9710) );
	o21ai_0 U10113( .A1(n6235), .A2(n7707), .B1(n9712), .Y(n4998) );
	mux2i_1 U10114( .A0(n9713), .A1(n6258), .S(n9714), .Y(n9712) );
	nor2_1 U10115( .A(n8185), .B(n8250), .Y(n9714) );
	nor2_1 U10116( .A(n6281), .B(n8095), .Y(n9713) );
	inv_1 U10117( .A(n10789), .Y(n8095) );
	inv_1 U10118( .A(n10785), .Y(n7707) );
	o21ai_0 U10119( .A1(n6235), .A2(n6009), .B1(n9715), .Y(n4997) );
	mux2i_1 U10120( .A0(n9716), .A1(n7021), .S(n9717), .Y(n9715) );
	nor3_1 U10121( .A(n9087), .B(n9243), .C(n7449), .Y(n9717) );
	nor2_1 U10122( .A(n6281), .B(n7362), .Y(n9716) );
	inv_1 U10123( .A(n10492), .Y(n7362) );
	nor3_1 U10124( .A(n9718), .B(n6350), .C(n9719), .Y(n4996) );
	o21ai_0 U10125( .A1(n6235), .A2(n7081), .B1(n9720), .Y(n4995) );
	mux2i_1 U10126( .A0(n9721), .A1(n9722), .S(n9723), .Y(n9720) );
	nor2_1 U10127( .A(n10568), .B(n6366), .Y(n9722) );
	nor2_1 U10128( .A(n8300), .B(n9724), .Y(n9721) );
	o221ai_1 U10129( .A1(n9643), .A2(n9725), .B1(n6220), .B2(n9726), .C1(n9727), .Y(n4994) );
	nand3_1 U10130( .A(n6341), .B(n9647), .C(n11840), .Y(n9727) );
	nand2_1 U10131( .A(n9728), .B(n8365), .Y(n9647) );
	o21ai_0 U10132( .A1(n6917), .A2(n7550), .B1(n9729), .Y(n9725) );
	inv_1 U10133( .A(n10843), .Y(n7550) );
	inv_1 U10134( .A(n9730), .Y(n9643) );
	o221ai_1 U10135( .A1(n9731), .A2(n5864), .B1(n6220), .B2(n6765), .C1(n9732), .Y(n4993) );
	nand3_1 U10136( .A(n7586), .B(n9733), .C(n7921), .Y(n9732) );
	xnor2_1 U10137( .A(n7563), .B(n10677), .Y(n9733) );
	inv_1 U10138( .A(n10729), .Y(n7563) );
	inv_1 U10139( .A(n10677), .Y(n6765) );
	a21oi_1 U10140( .A1(n6332), .A2(n6772), .B1(n8240), .Y(n9731) );
	inv_1 U10141( .A(n7921), .Y(n6772) );
	o32ai_1 U10142( .A1(n9734), .A2(n6347), .A3(n9735), .B1(n7213), .B2(n9477), .Y(n4992) );
	and2_0 U10143( .A(n6385), .B(g8344), .X(n4991) );
	o21ai_0 U10144( .A1(n6235), .A2(n6013), .B1(n9736), .Y(n4990) );
	mux2i_1 U10145( .A0(n9737), .A1(n6258), .S(n9738), .Y(n9736) );
	nor2_1 U10146( .A(n6628), .B(n9287), .Y(n9738) );
	nor2_1 U10147( .A(n6281), .B(n9279), .Y(n9737) );
	inv_1 U10148( .A(n10494), .Y(n9279) );
	o221ai_1 U10149( .A1(n9739), .A2(n5892), .B1(n6741), .B2(n8474), .C1(n6737), .Y(n4989) );
	inv_1 U10150( .A(n8840), .Y(n6737) );
	nor3_1 U10151( .A(n6742), .B(n7657), .C(n6743), .Y(n8840) );
	inv_1 U10152( .A(n6747), .Y(n8474) );
	nor2_1 U10153( .A(n6282), .B(n7088), .Y(n6747) );
	a21oi_1 U10154( .A1(n7088), .A2(n6381), .B1(n6437), .Y(n9739) );
	inv_1 U10155( .A(n6742), .Y(n7088) );
	o211ai_1 U10156( .A1(n9740), .A2(n7533), .B1(n10152), .C1(n9741), .Y(n6742) );
	o21ai_0 U10157( .A1(n6235), .A2(n9742), .B1(n9743), .Y(n4988) );
	mux2i_1 U10158( .A0(n9744), .A1(n9745), .S(n8151), .Y(n9743) );
	nor2_1 U10159( .A(n6351), .B(n9746), .Y(n9745) );
	and2_0 U10160( .A(n9746), .B(n6344), .X(n9744) );
	nand3_1 U10161( .A(n7767), .B(n6911), .C(n10910), .Y(n9746) );
	inv_1 U10162( .A(n10910), .Y(n9742) );
	mux2i_1 U10163( .A0(n9747), .A1(n6225), .S(n10593), .Y(n4987) );
	o21ai_0 U10164( .A1(n10210), .A2(n10603), .B1(n6343), .Y(n9747) );
	o221ai_1 U10165( .A1(n9748), .A2(n6308), .B1(n6220), .B2(n7305), .C1(n9749), .Y(n4986) );
	nand4_1 U10166( .A(n10484), .B(n9750), .C(n9751), .D(n9752), .Y(n9749) );
	nor2_1 U10167( .A(n6351), .B(n9753), .Y(n9751) );
	a21oi_1 U10168( .A1(n10268), .A2(g35), .B1(n10266), .Y(n9753) );
	a21oi_1 U10169( .A1(n7742), .A2(n10484), .B1(n9754), .Y(n9748) );
	a21oi_1 U10170( .A1(n9752), .A2(n9750), .B1(n9755), .Y(n9754) );
	inv_1 U10171( .A(n9756), .Y(n9755) );
	o21ai_0 U10172( .A1(n7742), .A2(n10484), .B1(n6957), .Y(n9756) );
	or2_0 U10173( .A(n6586), .B(n9757), .X(n9750) );
	o22ai_1 U10174( .A1(n7768), .A2(n8705), .B1(n7769), .B2(n9181), .Y(n4985) );
	o21ai_0 U10175( .A1(n6235), .A2(n6004), .B1(n9758), .Y(n4984) );
	mux2i_1 U10176( .A0(n9759), .A1(n6258), .S(n9760), .Y(n9758) );
	nor2_1 U10177( .A(n7353), .B(n7506), .Y(n9760) );
	nand2_1 U10178( .A(n11942), .B(n8980), .Y(n7506) );
	inv_1 U10179( .A(n10270), .Y(n8980) );
	nor2_1 U10180( .A(n6283), .B(n6005), .Y(n9759) );
	nor2_1 U10181( .A(n6352), .B(n9761), .Y(n4983) );
	o32ai_1 U10182( .A1(n8251), .A2(n10156), .A3(n8024), .B1(n6199), .B2(n5899), .Y(n4982) );
	inv_1 U10183( .A(n8187), .Y(n8024) );
	a21oi_1 U10184( .A1(n9762), .A2(n9119), .B1(n6368), .Y(n8187) );
	a21oi_1 U10185( .A1(n6197), .A2(n9763), .B1(n5962), .Y(n4981) );
	nand2_1 U10186( .A(n10464), .B(n6379), .Y(n9763) );
	o21ai_0 U10187( .A1(n9477), .A2(n6099), .B1(n9764), .Y(n4980) );
	mux2i_1 U10188( .A0(n9765), .A1(n9766), .S(n9767), .Y(n9764) );
	nor3_1 U10189( .A(n9478), .B(n11881), .C(n6307), .Y(n9766) );
	nand2_1 U10190( .A(n6222), .B(n9768), .Y(n9765) );
	nand3_1 U10191( .A(n11881), .B(n6377), .C(n9282), .Y(n9768) );
	o21ai_0 U10192( .A1(n6235), .A2(n9769), .B1(n9770), .Y(n4979) );
	mux2i_1 U10193( .A0(n9771), .A1(n9772), .S(n9213), .Y(n9770) );
	and3_1 U10194( .A(n8331), .B(n9217), .C(n6346), .X(n9772) );
	nand2_1 U10195( .A(n9175), .B(n9389), .Y(n9217) );
	o221ai_1 U10196( .A1(n7531), .A2(n9773), .B1(n6213), .B2(n5886), .C1(n9774), .Y(n4978) );
	nand3_1 U10197( .A(n10523), .B(n6377), .C(n6916), .Y(n9774) );
	a21oi_1 U10198( .A1(n9316), .A2(n9775), .B1(n6934), .Y(n6916) );
	o21ai_0 U10199( .A1(n6917), .A2(n9179), .B1(n9775), .Y(n9773) );
	inv_1 U10200( .A(n10844), .Y(n9179) );
	nor2_1 U10201( .A(n9776), .B(n6301), .Y(n4977) );
	a21oi_1 U10202( .A1(n10557), .A2(n7425), .B1(n9777), .Y(n9776) );
	mux2i_1 U10203( .A0(n9778), .A1(n9779), .S(n7424), .Y(n9777) );
	nand3_1 U10204( .A(n9780), .B(n8521), .C(n9781), .Y(n9779) );
	inv_1 U10205( .A(n8519), .Y(n8521) );
	nand2_1 U10206( .A(n7974), .B(n9782), .Y(n9778) );
	nor2_1 U10207( .A(n9783), .B(n8519), .Y(n7974) );
	o22ai_1 U10208( .A1(n6206), .A2(n5960), .B1(n6314), .B2(n9784), .Y(n4976) );
	nor2_1 U10209( .A(n6351), .B(n9785), .Y(n4975) );
	o21ai_0 U10210( .A1(n6236), .A2(n9724), .B1(n9786), .Y(n4974) );
	mux2i_1 U10211( .A0(n9787), .A1(n9788), .S(n9789), .Y(n9786) );
	nor2_1 U10212( .A(n10566), .B(n6367), .Y(n9788) );
	nor2_1 U10213( .A(n8300), .B(n8319), .Y(n9787) );
	inv_1 U10214( .A(n10566), .Y(n8319) );
	inv_1 U10215( .A(n10568), .Y(n9724) );
	o22ai_1 U10216( .A1(n6208), .A2(n5905), .B1(n9790), .B2(n7056), .Y(n4973) );
	or2_0 U10217( .A(n6314), .B(n8287), .X(n7056) );
	a21oi_1 U10218( .A1(n8286), .A2(n10180), .B1(n8285), .Y(n8287) );
	inv_1 U10219( .A(n10372), .Y(n8286) );
	xnor2_1 U10220( .A(n8742), .B(n5887), .Y(n9790) );
	nand3_1 U10221( .A(n10521), .B(n6819), .C(n11913), .Y(n8742) );
	o22ai_1 U10222( .A1(n6209), .A2(n6069), .B1(n8101), .B2(n9791), .Y(n4972) );
	mux2i_1 U10223( .A0(n9792), .A1(n9793), .S(n7094), .Y(n9791) );
	nand4_1 U10224( .A(n11807), .B(n6911), .C(g7916), .D(n7096), .Y(n7094) );
	nor2_1 U10225( .A(n6284), .B(n7095), .Y(n9793) );
	inv_1 U10226( .A(n10894), .Y(n7095) );
	nor2_1 U10227( .A(n10894), .B(n6365), .Y(n9792) );
	nor2_1 U10228( .A(n6284), .B(n8693), .Y(n4971) );
	o32ai_1 U10229( .A1(n6060), .A2(n6347), .A3(n9735), .B1(n9477), .B2(n9767), .Y(n4970) );
	inv_1 U10230( .A(n10648), .Y(n9767) );
	nand2_1 U10231( .A(n9735), .B(n6380), .Y(n9477) );
	o21ai_0 U10232( .A1(n6236), .A2(n9392), .B1(n9794), .Y(n4969) );
	mux2_1 U10233( .A0(n8643), .A1(n8636), .S(n11911), .X(n9794) );
	nand2_1 U10234( .A(n6338), .B(n9795), .Y(n8636) );
	nand2_1 U10235( .A(n8642), .B(n6335), .Y(n8643) );
	inv_1 U10236( .A(n9795), .Y(n8642) );
	nand4_1 U10237( .A(n8331), .B(g16693), .C(n10377), .D(n9145), .Y(n9795) );
	o21ai_0 U10238( .A1(n6236), .A2(n8440), .B1(n9796), .Y(n4968) );
	a22oi_1 U10239( .A1(n9272), .A2(n7345), .B1(n11764), .B2(n8583), .Y(n9796) );
	inv_1 U10240( .A(n6982), .Y(n8583) );
	nand2_1 U10241( .A(n6981), .B(n6379), .Y(n6982) );
	nor2_1 U10242( .A(n6934), .B(n9272), .Y(n6981) );
	and2_0 U10243( .A(n9797), .B(n6344), .X(n7345) );
	mux2i_1 U10244( .A0(n9798), .A1(n9492), .S(n7525), .Y(n9797) );
	and2_0 U10245( .A(n7527), .B(n7526), .X(n9798) );
	nor3_1 U10246( .A(n10238), .B(n10259), .C(n7347), .Y(n9272) );
	inv_1 U10247( .A(n10727), .Y(n8440) );
	o32ai_1 U10248( .A1(n9799), .A2(n10264), .A3(n9093), .B1(n9087), .B2(n9241), .Y(n4967) );
	o21ai_0 U10249( .A1(n10243), .A2(n9800), .B1(n6343), .Y(n9799) );
	o22ai_1 U10250( .A1(n6210), .A2(n9202), .B1(n9801), .B2(n8484), .Y(n4966) );
	a211oi_1 U10251( .A1(n10352), .A2(n6674), .B1(n9802), .C1(n8912), .Y(n9801) );
	nor2_1 U10252( .A(n6674), .B(n6466), .Y(n8912) );
	inv_1 U10253( .A(n10201), .Y(n9202) );
	mux2i_1 U10254( .A0(n9803), .A1(n9804), .S(n10198), .Y(n4965) );
	a21oi_1 U10255( .A1(n6598), .A2(n6592), .B1(n6437), .Y(n9804) );
	and3_1 U10256( .A(n8352), .B(n6370), .C(n9365), .X(n6598) );
	or2_0 U10257( .A(n6599), .B(n6592), .X(n9803) );
	nand3_1 U10258( .A(n9365), .B(n8352), .C(n6331), .Y(n6599) );
	o21ai_0 U10259( .A1(n6236), .A2(n9805), .B1(n9806), .Y(n4964) );
	mux2i_1 U10260( .A0(n9807), .A1(n6258), .S(n9808), .Y(n9806) );
	nor2_1 U10261( .A(n6906), .B(n8266), .Y(n9808) );
	nor2_1 U10262( .A(n6292), .B(n9482), .Y(n9807) );
	o221ai_1 U10263( .A1(n7427), .A2(n7040), .B1(n6219), .B2(n5871), .C1(n9809), .Y(n4963) );
	or4_1 U10264( .A(n7030), .B(n6314), .C(n7036), .D(n7347), .X(n9809) );
	nor2_1 U10265( .A(n7034), .B(n8885), .Y(n7036) );
	inv_1 U10266( .A(n10238), .Y(n7030) );
	inv_1 U10267( .A(n10249), .Y(n7040) );
	nand2_1 U10268( .A(n7347), .B(n6335), .Y(n7427) );
	inv_1 U10269( .A(n7522), .Y(n7347) );
	nand2_1 U10270( .A(n7525), .B(n7029), .Y(n7522) );
	o21ai_0 U10271( .A1(n9810), .A2(n7472), .B1(g17423), .Y(n7029) );
	inv_1 U10272( .A(n8726), .Y(n7472) );
	nor2_1 U10273( .A(n8723), .B(n6486), .Y(n8726) );
	and3_1 U10274( .A(n7527), .B(n9811), .C(n9812), .X(n7525) );
	nand3_1 U10275( .A(n10166), .B(n6803), .C(n10280), .Y(n9812) );
	nand2_1 U10276( .A(n10257), .B(n8070), .Y(n7527) );
	o221ai_1 U10277( .A1(n7168), .A2(n7172), .B1(n6219), .B2(n7004), .C1(n7173), .Y(n4962) );
	nand3_1 U10278( .A(n8242), .B(n6377), .C(n10322), .Y(n7173) );
	inv_1 U10279( .A(n10322), .Y(n7004) );
	inv_1 U10280( .A(n10635), .Y(n7172) );
	or2_0 U10281( .A(n6314), .B(n8242), .X(n7168) );
	nor3_1 U10282( .A(n6890), .B(n7578), .C(n5893), .Y(n8242) );
	o211ai_1 U10283( .A1(n9740), .A2(n9645), .B1(n9813), .C1(n8630), .Y(n7578) );
	inv_1 U10284( .A(n10335), .Y(n6890) );
	nor3_1 U10285( .A(n9814), .B(n10179), .C(n7469), .Y(n4961) );
	and3_1 U10286( .A(g12919), .B(n9815), .C(n10715), .X(n7469) );
	a222oi_1 U10287( .A1(n10715), .A2(n6341), .B1(n9816), .B2(g12919), .C1( n7083), .C2(n9817), .Y(n9814) );
	inv_1 U10288( .A(n9818), .Y(n9817) );
	inv_1 U10289( .A(n8300), .Y(n7083) );
	o32ai_1 U10290( .A1(n6311), .A2(g8277), .A3(n9819), .B1(n6199), .B2(n9820), .Y(n4960) );
	a21oi_1 U10291( .A1(g8215), .A2(n9820), .B1(n10620), .Y(n9819) );
	inv_1 U10292( .A(n10619), .Y(n9820) );
	o32ai_1 U10293( .A1(n9564), .A2(n6278), .A3(n7725), .B1(n6198), .B2(n9821), .Y(n4959) );
	inv_1 U10294( .A(n10655), .Y(n9821) );
	inv_1 U10295( .A(n10544), .Y(n7725) );
	nand2_1 U10296( .A(n10408), .B(n8758), .Y(n9564) );
	nor2_1 U10297( .A(n9822), .B(n8754), .Y(n8758) );
	o21ai_0 U10298( .A1(n6236), .A2(n9163), .B1(n9823), .Y(n4958) );
	mux2i_1 U10299( .A0(n9824), .A1(n6258), .S(n9825), .Y(n9823) );
	nor2_1 U10300( .A(n7386), .B(n8074), .Y(n9825) );
	nand2_1 U10301( .A(n9021), .B(n9600), .Y(n8074) );
	inv_1 U10302( .A(n10208), .Y(n9021) );
	nand2_1 U10303( .A(n11968), .B(n8558), .Y(n7386) );
	nor2_1 U10304( .A(n6293), .B(n5923), .Y(n9824) );
	inv_1 U10305( .A(n10813), .Y(n9163) );
	nor2_1 U10306( .A(n6352), .B(n9826), .Y(n4957) );
	o21ai_0 U10307( .A1(n6236), .A2(n8005), .B1(n9827), .Y(n4956) );
	a22oi_1 U10308( .A1(n6584), .A2(n6520), .B1(n7002), .B2(n11767), .Y(n9827) );
	inv_1 U10309( .A(n7605), .Y(n7002) );
	and2_0 U10310( .A(n6346), .B(n9828), .X(n6520) );
	o21ai_0 U10311( .A1(g23683), .A2(n9829), .B1(n6577), .Y(n9828) );
	o211ai_1 U10312( .A1(n10306), .A2(n9830), .B1(n9829), .C1(n9831), .Y(n6577) );
	a21oi_1 U10313( .A1(n9832), .A2(n9833), .B1(n6308), .Y(n4955) );
	o211ai_1 U10314( .A1(n9834), .A2(n9835), .B1(n6932), .C1(n8985), .Y(n9833) );
	inv_1 U10315( .A(n6936), .Y(n6932) );
	mux2_1 U10316( .A0(n6930), .A1(n7687), .S(n10416), .X(n9835) );
	nor2_1 U10317( .A(n6927), .B(n10194), .Y(n6930) );
	mux2i_1 U10318( .A0(n6933), .A1(n7694), .S(n5915), .Y(n9834) );
	inv_1 U10319( .A(n7682), .Y(n7694) );
	nor2_1 U10320( .A(n10368), .B(n10194), .Y(n7682) );
	nand2_1 U10321( .A(n10194), .B(n6927), .Y(n6933) );
	inv_1 U10322( .A(n10368), .Y(n6927) );
	o21ai_0 U10323( .A1(n8985), .A2(n6936), .B1(n10599), .Y(n9832) );
	nand2_1 U10324( .A(n10229), .B(n9836), .Y(n6936) );
	nand3_1 U10325( .A(n9837), .B(n9838), .C(n11967), .Y(n9836) );
	nor2_1 U10326( .A(n8400), .B(n9839), .Y(n8985) );
	o21ai_0 U10327( .A1(n6236), .A2(n9446), .B1(n9840), .Y(n4954) );
	a22oi_1 U10328( .A1(n10810), .A2(n6650), .B1(n7010), .B2(n6249), .Y(n9840) );
	inv_1 U10329( .A(n6546), .Y(n6650) );
	inv_1 U10330( .A(n10498), .Y(n9446) );
	nor3_1 U10331( .A(n9655), .B(n9841), .C(n6307), .Y(n4953) );
	a22oi_1 U10332( .A1(n10433), .A2(n8706), .B1(n10170), .B2(n10354), .Y(n9841) );
	nand2_1 U10333( .A(n7769), .B(n8705), .Y(n8706) );
	inv_1 U10334( .A(n10170), .Y(n8705) );
	inv_1 U10335( .A(n10354), .Y(n7769) );
	nand2_1 U10336( .A(n11955), .B(n9579), .Y(n9655) );
	o32ai_1 U10337( .A1(n6311), .A2(n10414), .A3(n7283), .B1(n6199), .B2(n9842), .Y(n4952) );
	nor2_1 U10338( .A(n9843), .B(n9842), .Y(n7283) );
	o22ai_1 U10339( .A1(n6210), .A2(n7142), .B1(n6302), .B2(n9844), .Y(n4951) );
	mux2i_1 U10340( .A0(n9845), .A1(n9846), .S(n7413), .Y(n9844) );
	xnor2_1 U10341( .A(n5883), .B(n10922), .Y(n9846) );
	nor2_1 U10342( .A(n10602), .B(n10460), .Y(n9845) );
	inv_1 U10343( .A(n10473), .Y(n7142) );
	o21ai_0 U10344( .A1(n6236), .A2(n9847), .B1(n9848), .Y(n4950) );
	a22oi_1 U10345( .A1(n11844), .A2(n8406), .B1(n8411), .B2(n9333), .Y(n9848) );
	nand2_1 U10346( .A(n9849), .B(n9850), .Y(n9333) );
	mux2i_1 U10347( .A0(n9851), .A1(n9852), .S(n9853), .Y(n9850) );
	xnor2_1 U10348( .A(n9165), .B(g12350), .Y(n9853) );
	nand3_1 U10349( .A(n9854), .B(n9855), .C(n9856), .Y(n9852) );
	nand3_1 U10350( .A(n8905), .B(g17607), .C(n10495), .Y(n9856) );
	nand3_1 U10351( .A(g17739), .B(n11806), .C(n8904), .Y(n9855) );
	nand3_1 U10352( .A(g14738), .B(n11815), .C(n8906), .Y(n9854) );
	nand3_1 U10353( .A(n9857), .B(n9858), .C(n9859), .Y(n9851) );
	nand3_1 U10354( .A(n8903), .B(n11817), .C(g17739), .Y(n9859) );
	nand3_1 U10355( .A(g17607), .B(n10777), .C(n8906), .Y(n9858) );
	nand3_1 U10356( .A(g14738), .B(n11883), .C(n8905), .Y(n9857) );
	mux2_1 U10357( .A0(n9860), .A1(n9861), .S(n9165), .X(n9849) );
	a221oi_1 U10358( .A1(n8905), .A2(n9862), .B1(n8903), .B2(n9863), .C1(n9864), .Y(n9861) );
	o32ai_1 U10359( .A1(n9865), .A2(n5924), .A3(n9866), .B1(n9867), .B2(n9421), .Y(n9864) );
	a22oi_1 U10360( .A1(n10769), .A2(g17646), .B1(g17715), .B2(n10770), .Y( n9867) );
	inv_1 U10361( .A(n8906), .Y(n9866) );
	o22ai_1 U10362( .A1(n7607), .A2(n9868), .B1(n8334), .B2(n9869), .Y(n9863) );
	inv_1 U10363( .A(n10768), .Y(n7607) );
	o22ai_1 U10364( .A1(n7230), .A2(n9870), .B1(n8154), .B2(n9871), .Y(n9862) );
	a221oi_1 U10365( .A1(n8906), .A2(n9872), .B1(n8903), .B2(n9873), .C1(n9874), .Y(n9860) );
	o32ai_1 U10366( .A1(n9865), .A2(n5926), .A3(n9420), .B1(n9875), .B2(n9421), .Y(n9874) );
	inv_1 U10367( .A(n8904), .Y(n9421) );
	nor2_1 U10368( .A(n8408), .B(n10193), .Y(n8904) );
	a22oi_1 U10369( .A1(g12350), .A2(n10773), .B1(n10774), .B2(g17819), .Y( n9875) );
	inv_1 U10370( .A(n8905), .Y(n9420) );
	nor2_1 U10371( .A(n9876), .B(n10367), .Y(n8905) );
	o22ai_1 U10372( .A1(n8267), .A2(n9877), .B1(n9878), .B2(n9847), .Y(n9873) );
	inv_1 U10373( .A(n10772), .Y(n8267) );
	o22ai_1 U10374( .A1(n6901), .A2(n9870), .B1(n9871), .B2(n9482), .Y(n9872) );
	inv_1 U10375( .A(n10775), .Y(n9482) );
	inv_1 U10376( .A(n10776), .Y(n6901) );
	nor2_1 U10377( .A(n10367), .B(n10193), .Y(n8906) );
	nor2_1 U10378( .A(n8902), .B(n6300), .Y(n8411) );
	nor2_1 U10379( .A(n6293), .B(n9879), .Y(n8406) );
	inv_1 U10380( .A(n10771), .Y(n9847) );
	o21ai_0 U10381( .A1(n6236), .A2(n9880), .B1(n9881), .Y(n4949) );
	mux2i_1 U10382( .A0(n9882), .A1(n8256), .S(n5941), .Y(n9881) );
	nor2_1 U10383( .A(n9880), .B(n6367), .Y(n8256) );
	nor2_1 U10384( .A(n10543), .B(n6301), .Y(n9882) );
	inv_1 U10385( .A(n10543), .Y(n9880) );
	o21ai_0 U10386( .A1(n6236), .A2(n6989), .B1(n9883), .Y(n4948) );
	a22oi_1 U10387( .A1(n11776), .A2(n9884), .B1(n7303), .B2(n6959), .Y(n9883) );
	inv_1 U10388( .A(n10733), .Y(n6989) );
	o32ai_1 U10389( .A1(n7321), .A2(n10158), .A3(n9885), .B1(n6198), .B2(n5904), .Y(n4947) );
	nor3_1 U10390( .A(n8025), .B(n10273), .C(n10156), .Y(n4946) );
	o21ai_0 U10391( .A1(n9512), .A2(n8830), .B1(n6343), .Y(n8025) );
	o21ai_0 U10392( .A1(n7465), .A2(n6039), .B1(n9886), .Y(n4945) );
	mux2i_1 U10393( .A0(n9887), .A1(n9888), .S(n9889), .Y(n9886) );
	nor3_1 U10394( .A(n9017), .B(n11884), .C(n6306), .Y(n9888) );
	nand2_1 U10395( .A(n6224), .B(n9890), .Y(n9887) );
	nand3_1 U10396( .A(n6663), .B(n6377), .C(n11884), .Y(n9890) );
	o22ai_1 U10397( .A1(n6211), .A2(n6065), .B1(n9891), .B2(n6295), .Y(n4944) );
	nor2_1 U10398( .A(n10211), .B(n10576), .Y(n9891) );
	o21ai_0 U10399( .A1(n6236), .A2(n9892), .B1(n9893), .Y(n4943) );
	mux2i_1 U10400( .A0(n9894), .A1(n6258), .S(n9895), .Y(n9893) );
	nor2_1 U10401( .A(n6906), .B(n7229), .Y(n9895) );
	inv_1 U10402( .A(n9212), .Y(n7229) );
	nor2_1 U10403( .A(n9805), .B(n10207), .Y(n9212) );
	nor2_1 U10404( .A(n6292), .B(n8154), .Y(n9894) );
	inv_1 U10405( .A(n10765), .Y(n8154) );
	mux2i_1 U10406( .A0(n9896), .A1(n6225), .S(n11799), .Y(n4942) );
	nand2_1 U10407( .A(g7540), .B(n6335), .Y(n9896) );
	o22ai_1 U10408( .A1(n6810), .A2(n9632), .B1(n7546), .B2(n8708), .Y(n4941) );
	inv_1 U10409( .A(n10428), .Y(n8708) );
	inv_1 U10410( .A(n10859), .Y(n9632) );
	o22ai_1 U10411( .A1(n7060), .A2(n6630), .B1(n6632), .B2(n7774), .Y(n4940) );
	inv_1 U10412( .A(n10449), .Y(n7774) );
	o22ai_1 U10413( .A1(n6815), .A2(n6810), .B1(n6817), .B2(n7775), .Y(n4939) );
	inv_1 U10414( .A(n10329), .Y(n7775) );
	inv_1 U10415( .A(n7746), .Y(n6817) );
	nor2_1 U10416( .A(n9195), .B(n6299), .Y(n7746) );
	inv_1 U10417( .A(n10168), .Y(n6815) );
	o22ai_1 U10418( .A1(n6304), .A2(n8986), .B1(n6193), .B2(n9897), .Y(n4938) );
	and2_0 U10419( .A(n6386), .B(g9617), .X(n4937) );
	o221ai_1 U10420( .A1(n8114), .A2(n9898), .B1(n6217), .B2(n9899), .C1(n9900), .Y(n4936) );
	nand3_1 U10421( .A(n6340), .B(n8118), .C(n10672), .Y(n9900) );
	nand2_1 U10422( .A(n9728), .B(n10244), .Y(n8118) );
	nor2_1 U10423( .A(n9424), .B(n6633), .Y(n9728) );
	o21ai_0 U10424( .A1(n6917), .A2(n9899), .B1(n9729), .Y(n9898) );
	inv_1 U10425( .A(n7531), .Y(n9729) );
	nand3_1 U10426( .A(g35), .B(n9901), .C(n9902), .Y(n7531) );
	nand2_1 U10427( .A(g111), .B(n9390), .Y(n9901) );
	inv_1 U10428( .A(n10735), .Y(n9899) );
	inv_1 U10429( .A(n9903), .Y(n8114) );
	o21ai_0 U10430( .A1(n6236), .A2(n5864), .B1(n9904), .Y(n4935) );
	mux2_1 U10431( .A0(n7814), .A1(n7809), .S(n10693), .X(n9904) );
	or2_0 U10432( .A(n6314), .B(n9107), .X(n7809) );
	o22ai_1 U10433( .A1(n6305), .A2(n9905), .B1(n6193), .B2(n8588), .Y(n4934) );
	o22ai_1 U10434( .A1(n8142), .A2(n8327), .B1(n8145), .B2(n9906), .Y(n4933) );
	o21ai_0 U10435( .A1(n9907), .A2(n10594), .B1(n6342), .Y(n9906) );
	a21oi_1 U10436( .A1(n9908), .A2(n9909), .B1(n9128), .Y(n9907) );
	mux2i_1 U10437( .A0(n9140), .A1(n9141), .S(n5916), .Y(n9909) );
	nor2_1 U10438( .A(n10369), .B(n10195), .Y(n9141) );
	nor2_1 U10439( .A(n9910), .B(n10369), .Y(n9140) );
	mux2i_1 U10440( .A0(n9145), .A1(n9139), .S(n9769), .Y(n9908) );
	inv_1 U10441( .A(n10418), .Y(n9769) );
	nor2_1 U10442( .A(n9213), .B(n10195), .Y(n9139) );
	inv_1 U10443( .A(n8148), .Y(n8145) );
	nor2_1 U10444( .A(n9068), .B(n9911), .Y(n8148) );
	inv_1 U10445( .A(n9771), .Y(n8327) );
	nor2_1 U10446( .A(n6294), .B(n8331), .Y(n9771) );
	inv_1 U10447( .A(n9128), .Y(n8331) );
	nand2_1 U10448( .A(n10197), .B(n9912), .Y(n9128) );
	nand3_1 U10449( .A(n11810), .B(n9913), .C(n9388), .Y(n9912) );
	inv_1 U10450( .A(n10594), .Y(n8142) );
	o21ai_0 U10451( .A1(n6236), .A2(n9914), .B1(n9915), .Y(n4932) );
	o32ai_1 U10452( .A1(n6684), .A2(n10937), .A3(n10380), .B1(n9916), .B2(n9917), .Y(n9915) );
	a21oi_1 U10453( .A1(n6684), .A2(n7799), .B1(n6308), .Y(n9917) );
	inv_1 U10454( .A(n10443), .Y(n7799) );
	nor4_1 U10455( .A(n9918), .B(n9914), .C(n6347), .D(n5951), .Y(n9916) );
	nand2_1 U10456( .A(n11885), .B(n11886), .Y(n9918) );
	inv_1 U10457( .A(g4564), .Y(n9914) );
	o21ai_0 U10458( .A1(n6236), .A2(n8749), .B1(n9919), .Y(n4931) );
	mux2i_1 U10459( .A0(n9920), .A1(n6259), .S(n9921), .Y(n9919) );
	nor2_1 U10460( .A(n7965), .B(n8941), .Y(n9921) );
	nor2_1 U10461( .A(n6294), .B(n8931), .Y(n9920) );
	inv_1 U10462( .A(n10826), .Y(n8931) );
	o21ai_0 U10463( .A1(n6236), .A2(n6006), .B1(n9922), .Y(n4930) );
	mux2i_1 U10464( .A0(n9923), .A1(n6259), .S(n9924), .Y(n9922) );
	nor2_1 U10465( .A(n6466), .B(n8483), .Y(n9924) );
	nand2_1 U10466( .A(n10201), .B(n6566), .Y(n6466) );
	nor2_1 U10467( .A(n6291), .B(n5987), .Y(n9923) );
	o32ai_1 U10468( .A1(n6311), .A2(n10420), .A3(n8380), .B1(n6200), .B2(n8769), .Y(n4929) );
	nor2_1 U10469( .A(n9925), .B(n8769), .Y(n8380) );
	o22ai_1 U10470( .A1(n6212), .A2(n8539), .B1(n9926), .B2(n6297), .Y(n4928) );
	nor4_1 U10471( .A(n10657), .B(n10577), .C(n10184), .D(n9927), .Y(n9926) );
	o21ai_0 U10472( .A1(n8673), .A2(n9928), .B1(n9929), .Y(n4927) );
	mux2i_1 U10473( .A0(n9930), .A1(n9931), .S(n9570), .Y(n9929) );
	inv_1 U10474( .A(n10654), .Y(n9570) );
	nor3_1 U10475( .A(n6720), .B(n11889), .C(n6306), .Y(n9931) );
	inv_1 U10476( .A(n8385), .Y(n6720) );
	nand2_1 U10477( .A(n6222), .B(n9932), .Y(n9930) );
	nand3_1 U10478( .A(n8385), .B(n6378), .C(n11889), .Y(n9932) );
	o21ai_0 U10479( .A1(n6236), .A2(n5925), .B1(n9933), .Y(n4926) );
	mux2i_1 U10480( .A0(n9934), .A1(n6259), .S(n9935), .Y(n9933) );
	nor2_1 U10481( .A(n6668), .B(n8251), .Y(n9935) );
	nor2_1 U10482( .A(n6293), .B(n7700), .Y(n9934) );
	o22ai_1 U10483( .A1(n6211), .A2(n9936), .B1(n9937), .B2(n7239), .Y(n4925) );
	inv_1 U10484( .A(n9938), .Y(n7239) );
	a211oi_1 U10485( .A1(n10289), .A2(n8357), .B1(n7824), .C1(n6298), .Y(n9938) );
	inv_1 U10486( .A(n8107), .Y(n7824) );
	nor2_1 U10487( .A(n8106), .B(n8353), .Y(n8357) );
	xnor2_1 U10488( .A(n7825), .B(n10277), .Y(n9937) );
	inv_1 U10489( .A(n10600), .Y(n9936) );
	o32ai_1 U10490( .A1(n9939), .A2(n6348), .A3(n8925), .B1(n8926), .B2(n9382), .Y(n4924) );
	inv_1 U10491( .A(n10625), .Y(n9382) );
	inv_1 U10492( .A(n10692), .Y(n9939) );
	o21ai_0 U10493( .A1(n6236), .A2(n9940), .B1(n9941), .Y(n4923) );
	mux2i_1 U10494( .A0(n9942), .A1(n9943), .S(n9944), .Y(n9941) );
	a21oi_1 U10495( .A1(n9945), .A2(n6408), .B1(n6307), .Y(n4922) );
	inv_1 U10496( .A(n8101), .Y(n6408) );
	nor4_1 U10497( .A(n7096), .B(n7098), .C(n9946), .D(n7097), .Y(n8101) );
	a21oi_1 U10498( .A1(n9780), .A2(n9781), .B1(n9947), .Y(n7097) );
	nor3_1 U10499( .A(n9540), .B(n8518), .C(n5907), .Y(n9781) );
	nor2_1 U10500( .A(n8103), .B(n6911), .Y(n9946) );
	nand3_1 U10501( .A(n10457), .B(n7091), .C(n10472), .Y(n7096) );
	inv_1 U10502( .A(n10875), .Y(n7091) );
	xnor2_1 U10503( .A(n10248), .B(g7916), .Y(n9945) );
	o21ai_0 U10504( .A1(n6237), .A2(n9557), .B1(n9948), .Y(n4921) );
	mux2_1 U10505( .A0(n8848), .A1(n8841), .S(n11919), .X(n9948) );
	nand2_1 U10506( .A(n6338), .B(n9949), .Y(n8841) );
	nand2_1 U10507( .A(n8847), .B(n6335), .Y(n8848) );
	inv_1 U10508( .A(n9949), .Y(n8847) );
	nand4_1 U10509( .A(g17646), .B(n10375), .C(n8903), .D(n9879), .Y(n9949) );
	inv_1 U10510( .A(n8902), .Y(n9879) );
	nand2_1 U10511( .A(n11872), .B(n9950), .Y(n8902) );
	nand3_1 U10512( .A(n8348), .B(n9838), .C(n11890), .Y(n9950) );
	inv_1 U10513( .A(n10212), .Y(n9557) );
	o32ai_1 U10514( .A1(n9951), .A2(n6348), .A3(n6988), .B1(n6952), .B2(n6956), .Y(n4920) );
	inv_1 U10515( .A(n10630), .Y(n6956) );
	inv_1 U10516( .A(n10697), .Y(n9951) );
	o32ai_1 U10517( .A1(n6033), .A2(n9952), .A3(n6312), .B1(n9953), .B2(n9954), .Y(n4919) );
	nor2_1 U10518( .A(n9955), .B(n6437), .Y(n9953) );
	nor4_1 U10519( .A(n11891), .B(n6367), .C(n6711), .D(n6715), .Y(n9955) );
	a21oi_1 U10520( .A1(n10517), .A2(n9954), .B1(n6715), .Y(n9952) );
	inv_1 U10521( .A(n10422), .Y(n9954) );
	o22ai_1 U10522( .A1(n9956), .A2(n9944), .B1(n9957), .B2(n6537), .Y(n4918) );
	a21oi_1 U10523( .A1(n6332), .A2(n9944), .B1(n9942), .Y(n9957) );
	o21ai_0 U10524( .A1(n10317), .A2(n6314), .B1(n9958), .Y(n9942) );
	inv_1 U10525( .A(n10925), .Y(n9944) );
	a21oi_1 U10526( .A1(n9943), .A2(n6537), .B1(n6437), .Y(n9956) );
	inv_1 U10527( .A(n10876), .Y(n6537) );
	nor3_1 U10528( .A(n9940), .B(n6350), .C(n9959), .Y(n9943) );
	o32ai_1 U10529( .A1(n9960), .A2(n10260), .A3(n7113), .B1(n7110), .B2(n7883), .Y(n4917) );
	nand2_1 U10530( .A(n7884), .B(n6335), .Y(n7110) );
	nor2_1 U10531( .A(n8092), .B(n8885), .Y(n7113) );
	o21ai_0 U10532( .A1(n10239), .A2(n9961), .B1(n6343), .Y(n9960) );
	o221ai_1 U10533( .A1(n9962), .A2(n9963), .B1(n6217), .B2(n9362), .C1(n9964), .Y(n4916) );
	nand3_1 U10534( .A(n6340), .B(n7098), .C(n10875), .Y(n9964) );
	o211ai_1 U10535( .A1(n9965), .A2(n8896), .B1(n9966), .C1(n6839), .Y(n4915) );
	nand3_1 U10536( .A(n9967), .B(n6330), .C(n11973), .Y(n6839) );
	nand3_1 U10537( .A(n6841), .B(n8897), .C(n11890), .Y(n9966) );
	inv_1 U10538( .A(n9968), .Y(n8897) );
	nor2_1 U10539( .A(n6294), .B(n9967), .Y(n6841) );
	inv_1 U10540( .A(n10598), .Y(n8896) );
	a21oi_1 U10541( .A1(n9968), .A2(n6843), .B1(n6437), .Y(n9965) );
	nor2_1 U10542( .A(n9967), .B(n6365), .Y(n6843) );
	nor3_1 U10543( .A(g8132), .B(n10601), .C(n9969), .Y(n9967) );
	nor2_1 U10544( .A(n8351), .B(n8400), .Y(n9968) );
	o21ai_0 U10545( .A1(n6237), .A2(n7462), .B1(n9970), .Y(n4914) );
	mux2i_1 U10546( .A0(n9971), .A1(n7118), .S(n9972), .Y(n9970) );
	nor2_1 U10547( .A(n10240), .B(n7760), .Y(n9972) );
	nand2_1 U10548( .A(n10251), .B(n9533), .Y(n7760) );
	inv_1 U10549( .A(n7433), .Y(n9533) );
	nor2_1 U10550( .A(n9535), .B(n8880), .Y(n7433) );
	inv_1 U10551( .A(n8877), .Y(n8880) );
	o21ai_0 U10552( .A1(n9810), .A2(n8722), .B1(g17320), .Y(n8877) );
	and2_0 U10553( .A(n6346), .B(n9973), .X(n7118) );
	o21ai_0 U10554( .A1(n9535), .A2(n9492), .B1(n9529), .Y(n9973) );
	o211ai_1 U10555( .A1(n10256), .A2(n9974), .B1(n9535), .C1(n9975), .Y(n9529) );
	inv_1 U10556( .A(n10469), .Y(n9492) );
	o211ai_1 U10557( .A1(n10508), .A2(n8565), .B1(n9976), .C1(n9811), .Y(n9535) );
	nand3_1 U10558( .A(n6804), .B(n6803), .C(n10166), .Y(n9976) );
	nor2_1 U10559( .A(n6292), .B(n6007), .Y(n9971) );
	inv_1 U10560( .A(n10722), .Y(n7462) );
	o221ai_1 U10561( .A1(n7387), .A2(n6485), .B1(n6217), .B2(n9481), .C1(n9977), .Y(n4913) );
	nand3_1 U10562( .A(n10468), .B(g35), .C(n61), .Y(n9977) );
	nor2_1 U10563( .A(n7281), .B(n6366), .Y(n61) );
	nand2_1 U10564( .A(n6337), .B(n7281), .Y(n6485) );
	inv_1 U10565( .A(g7946), .Y(n7281) );
	inv_1 U10566( .A(n10874), .Y(n7387) );
	o211ai_1 U10567( .A1(n6203), .A2(n9224), .B1(n8232), .C1(n9978), .Y(n4912) );
	mux2i_1 U10568( .A0(n9979), .A1(n9980), .S(n7122), .Y(n9978) );
	inv_1 U10569( .A(n10434), .Y(n7122) );
	and2_0 U10570( .A(n6387), .B(n9981), .X(n9980) );
	nor2_1 U10571( .A(n9981), .B(n6299), .Y(n9979) );
	nor2_1 U10572( .A(n9225), .B(n9224), .Y(n9981) );
	nand2_1 U10573( .A(n9581), .B(n10288), .Y(n9225) );
	nor2_1 U10574( .A(n9121), .B(n9322), .Y(n9581) );
	nand2_1 U10575( .A(n9120), .B(n10163), .Y(n9121) );
	nor2_1 U10576( .A(n9982), .B(n8818), .Y(n9120) );
	inv_1 U10577( .A(n10425), .Y(n9224) );
	o22ai_1 U10578( .A1(n6210), .A2(n6480), .B1(n9983), .B2(n9984), .Y(n4911) );
	a222oi_1 U10579( .A1(n4709), .A2(n6482), .B1(n9985), .B2(n6382), .C1(n9986), .C2(n6341), .Y(n9984) );
	o22ai_1 U10580( .A1(n6210), .A2(n9987), .B1(n9988), .B2(n6298), .Y(n4910) );
	nor2_1 U10581( .A(n10232), .B(n10575), .Y(n9988) );
	inv_1 U10582( .A(n10576), .Y(n9987) );
	and2_0 U10583( .A(n6346), .B(n10884), .X(n4909) );
	o22ai_1 U10584( .A1(n6210), .A2(n8070), .B1(n9989), .B2(n6297), .Y(n4908) );
	nor2_1 U10585( .A(n10590), .B(n9481), .Y(n9989) );
	o32ai_1 U10586( .A1(n9990), .A2(n7941), .A3(n6312), .B1(n9991), .B2(n7940), .Y(n4907) );
	inv_1 U10587( .A(n10877), .Y(n7940) );
	a21oi_1 U10588( .A1(n7941), .A2(n6383), .B1(n6437), .Y(n9991) );
	o32ai_1 U10589( .A1(n6310), .A2(n9992), .A3(n9993), .B1(n6199), .B2(n8565), .Y(n4906) );
	inv_1 U10590( .A(n10256), .Y(n8565) );
	a21oi_1 U10591( .A1(n9432), .A2(n8974), .B1(n10906), .Y(n9993) );
	nor3_1 U10592( .A(n9994), .B(n7922), .C(n7279), .Y(n9992) );
	xnor2_1 U10593( .A(n10258), .B(n8698), .Y(n9994) );
	o21ai_0 U10594( .A1(n6237), .A2(n9486), .B1(n9995), .Y(n4905) );
	mux2i_1 U10595( .A0(n9996), .A1(n6259), .S(n9997), .Y(n9995) );
	nor2_1 U10596( .A(n7611), .B(n8266), .Y(n9997) );
	nand2_1 U10597( .A(n9209), .B(n9805), .Y(n8266) );
	inv_1 U10598( .A(n10207), .Y(n9209) );
	nand2_1 U10599( .A(n11956), .B(n8688), .Y(n7611) );
	nor2_1 U10600( .A(n6293), .B(n5926), .Y(n9996) );
	inv_1 U10601( .A(n10774), .Y(n9486) );
	and2_0 U10602( .A(n6345), .B(n10885), .X(n4904) );
	o221ai_1 U10603( .A1(n9998), .A2(n5894), .B1(n9042), .B2(n8955), .C1(n9038), .Y(n4903) );
	inv_1 U10604( .A(n8958), .Y(n9038) );
	nor3_1 U10605( .A(n7633), .B(n7657), .C(n9043), .Y(n8958) );
	inv_1 U10606( .A(n7625), .Y(n8955) );
	a21oi_1 U10607( .A1(n9083), .A2(n6381), .B1(n6437), .Y(n9998) );
	o21ai_0 U10608( .A1(n6237), .A2(n5939), .B1(n9999), .Y(n4902) );
	mux2i_1 U10609( .A0(n10000), .A1(n6259), .S(n10001), .Y(n9999) );
	nor2_1 U10610( .A(n6492), .B(n7178), .Y(n10001) );
	nand2_1 U10611( .A(n11943), .B(n10274), .Y(n6492) );
	nor2_1 U10612( .A(n6282), .B(n8610), .Y(n10000) );
	inv_1 U10613( .A(n10796), .Y(n8610) );
	a21oi_1 U10614( .A1(n6198), .A2(n10002), .B1(n6879), .Y(n4901) );
	nand2_1 U10615( .A(n6882), .B(n8854), .Y(n10002) );
	and2_0 U10616( .A(n6387), .B(g26960), .X(n4900) );
	o21ai_0 U10617( .A1(n6240), .A2(n9617), .B1(n10003), .Y(n4899) );
	a22oi_1 U10618( .A1(n10771), .A2(n6861), .B1(n7248), .B2(n6249), .Y(n10003) );
	inv_1 U10619( .A(n6751), .Y(n6861) );
	inv_1 U10620( .A(n10495), .Y(n9617) );
	o32ai_1 U10621( .A1(n6801), .A2(n8699), .A3(n6312), .B1(n10004), .B2(n8424), .Y(n4898) );
	o21ai_0 U10622( .A1(n6237), .A2(n9258), .B1(n10005), .Y(n4897) );
	mux2i_1 U10623( .A0(n10006), .A1(n6259), .S(n10007), .Y(n10005) );
	nor2_1 U10624( .A(n6858), .B(n7880), .Y(n10007) );
	nand2_1 U10625( .A(n10271), .B(n5900), .Y(n7880) );
	nand2_1 U10626( .A(n10206), .B(n9046), .Y(n6858) );
	nor2_1 U10627( .A(n6280), .B(n6008), .Y(n10006) );
	o22ai_1 U10628( .A1(n6305), .A2(n10008), .B1(n6193), .B2(n10009), .Y(n4896) );
	o21ai_0 U10629( .A1(n6237), .A2(n6082), .B1(n10010), .Y(n4895) );
	mux2i_1 U10630( .A0(n10011), .A1(n10012), .S(n10013), .Y(n10010) );
	nor2_1 U10631( .A(n6353), .B(n10014), .Y(n10012) );
	nor2_1 U10632( .A(n10015), .B(n8048), .Y(n10011) );
	o221ai_1 U10633( .A1(n10016), .A2(n5895), .B1(n7722), .B2(n8551), .C1(n7718), .Y(n4894) );
	inv_1 U10634( .A(n8752), .Y(n7718) );
	a21oi_1 U10635( .A1(n7220), .A2(n6381), .B1(n6437), .Y(n10016) );
	o21ai_0 U10636( .A1(n6237), .A2(n7451), .B1(n10017), .Y(n4893) );
	mux2i_1 U10637( .A0(n10018), .A1(n7021), .S(n10019), .Y(n10017) );
	nor2_1 U10638( .A(n10243), .B(n10020), .Y(n10019) );
	nor2_1 U10639( .A(n6292), .B(n6009), .Y(n10018) );
	inv_1 U10640( .A(n10725), .Y(n7451) );
	o21ai_0 U10641( .A1(n6237), .A2(n7700), .B1(n10021), .Y(n4892) );
	mux2i_1 U10642( .A0(n10022), .A1(n6259), .S(n10023), .Y(n10021) );
	nor2_1 U10643( .A(n8185), .B(n6668), .Y(n10023) );
	nor2_1 U10644( .A(n6293), .B(n7899), .Y(n10022) );
	inv_1 U10645( .A(n10779), .Y(n7899) );
	inv_1 U10646( .A(n10783), .Y(n7700) );
	nor2_1 U10647( .A(n6352), .B(n10024), .Y(n4891) );
	o21ai_0 U10648( .A1(n6237), .A2(n7213), .B1(n10025), .Y(n4890) );
	a22oi_1 U10649( .A1(n10026), .A2(n9262), .B1(n9261), .B2(n10897), .Y(n10025) );
	xnor2_1 U10650( .A(n10027), .B(n9263), .Y(n10026) );
	nand2_1 U10651( .A(n10028), .B(n10029), .Y(n9263) );
	mux2i_1 U10652( .A0(n10030), .A1(n10031), .S(n10032), .Y(n10029) );
	xnor2_1 U10653( .A(n9842), .B(g12422), .Y(n10032) );
	nand3_1 U10654( .A(n10033), .B(n10034), .C(n10035), .Y(n10031) );
	nand3_1 U10655( .A(n8397), .B(g17760), .C(n11851), .Y(n10035) );
	nand3_1 U10656( .A(n8395), .B(g14779), .C(n11833), .Y(n10034) );
	nand3_1 U10657( .A(n8394), .B(g17649), .C(n10494), .Y(n10033) );
	nand3_1 U10658( .A(n10036), .B(n10037), .C(n10038), .Y(n10030) );
	nand3_1 U10659( .A(n8396), .B(n11893), .C(g17760), .Y(n10038) );
	nand3_1 U10660( .A(g17649), .B(n10764), .C(n8395), .Y(n10037) );
	nand3_1 U10661( .A(n11894), .B(g14779), .C(n8394), .Y(n10036) );
	mux2_1 U10662( .A0(n10039), .A1(n10040), .S(n9842), .X(n10028) );
	a221oi_1 U10663( .A1(n8397), .A2(n10041), .B1(n8396), .B2(n10042), .C1( n10043), .Y(n10040) );
	o32ai_1 U10664( .A1(n10044), .A2(n5928), .A3(n10045), .B1(n10046), .B2( n10047), .Y(n10043) );
	a22oi_1 U10665( .A1(g13085), .A2(n10752), .B1(n10753), .B2(n10222), .Y( n10046) );
	o22ai_1 U10666( .A1(n8930), .A2(n10048), .B1(n10049), .B2(n9283), .Y(n10042) );
	o22ai_1 U10667( .A1(n7497), .A2(n10050), .B1(n10051), .B2(n8078), .Y(n10041) );
	inv_1 U10668( .A(n10756), .Y(n8078) );
	a221oi_1 U10669( .A1(n8397), .A2(n10052), .B1(n8396), .B2(n10053), .C1( n10054), .Y(n10039) );
	o32ai_1 U10670( .A1(n10044), .A2(n5927), .A3(n10047), .B1(n10055), .B2( n10045), .Y(n10054) );
	inv_1 U10671( .A(n8395), .Y(n10045) );
	nor2_1 U10672( .A(n10366), .B(n10192), .Y(n8395) );
	a22oi_1 U10673( .A1(g13085), .A2(n10762), .B1(n10222), .B2(n10763), .Y( n10055) );
	o22ai_1 U10674( .A1(n6629), .A2(n10050), .B1(n10051), .B2(n9259), .Y(n10053) );
	inv_1 U10675( .A(n10758), .Y(n9259) );
	inv_1 U10676( .A(n10759), .Y(n6629) );
	o22ai_1 U10677( .A1(n7881), .A2(n10048), .B1(n10049), .B2(n9258), .Y(n10052) );
	inv_1 U10678( .A(n10760), .Y(n9258) );
	inv_1 U10679( .A(n10761), .Y(n7881) );
	nand2_1 U10680( .A(n10897), .B(n10056), .Y(n10027) );
	nand3_1 U10681( .A(g17685), .B(n8396), .C(n10374), .Y(n10056) );
	inv_1 U10682( .A(n10310), .Y(n7213) );
	o32ai_1 U10683( .A1(n6310), .A2(n10057), .A3(n10058), .B1(n6200), .B2(n6801), .Y(n4889) );
	inv_1 U10684( .A(n10430), .Y(n6801) );
	a21oi_1 U10685( .A1(n9432), .A2(n8567), .B1(n10909), .Y(n10058) );
	nor3_1 U10686( .A(n10430), .B(n11816), .C(n7922), .Y(n9432) );
	nor3_1 U10687( .A(n10059), .B(n7922), .C(n8722), .Y(n10057) );
	inv_1 U10688( .A(n8567), .Y(n8722) );
	nor2_1 U10689( .A(n8723), .B(n10237), .Y(n8567) );
	xnor2_1 U10690( .A(n10256), .B(n8698), .Y(n10059) );
	nand2_1 U10691( .A(n10060), .B(n19677), .Y(n8698) );
	o32ai_1 U10692( .A1(n8424), .A2(n8699), .A3(n6312), .B1(n10004), .B2(n5933), .Y(n4888) );
	a21oi_1 U10693( .A1(n6378), .A2(n8699), .B1(n6437), .Y(n10004) );
	nor3_1 U10694( .A(n10237), .B(n10923), .C(n7922), .Y(n8699) );
	inv_1 U10695( .A(g13272), .Y(n7922) );
	inv_1 U10696( .A(n10440), .Y(n8424) );
	and2_0 U10697( .A(n6387), .B(g8215), .X(n4887) );
	o22ai_1 U10698( .A1(n6208), .A2(n7307), .B1(n10061), .B2(n10062), .Y(n4886) );
	a22oi_1 U10699( .A1(n7662), .A2(g25167), .B1(n10586), .B2(n6337), .Y(n10062) );
	nor2_1 U10700( .A(n9377), .B(n6301), .Y(n7662) );
	nor4_1 U10701( .A(n10268), .B(n9377), .C(n7487), .D(n10063), .Y(n10061) );
	inv_1 U10702( .A(n10286), .Y(n7487) );
	o211ai_1 U10703( .A1(n9740), .A2(n8303), .B1(n8223), .C1(n9741), .Y(n9377) );
	inv_1 U10704( .A(n10737), .Y(n7307) );
	o21ai_0 U10705( .A1(n6237), .A2(n7109), .B1(n10064), .Y(n4885) );
	mux2i_1 U10706( .A0(n10065), .A1(n10066), .S(n10067), .Y(n10064) );
	nor2_1 U10707( .A(n10396), .B(n6366), .Y(n10066) );
	nor2_1 U10708( .A(n7108), .B(n7588), .Y(n10065) );
	o22ai_1 U10709( .A1(n6304), .A2(n10009), .B1(n6193), .B2(n7263), .Y(n4884) );
	inv_1 U10710( .A(n10705), .Y(n7263) );
	nor2_1 U10711( .A(n10068), .B(n10069), .Y(n4883) );
	o21ai_0 U10712( .A1(n6237), .A2(n10070), .B1(n10071), .Y(n4882) );
	mux2i_1 U10713( .A0(n10072), .A1(n6259), .S(n10073), .Y(n10071) );
	nor2_1 U10714( .A(n8082), .B(n9287), .Y(n10073) );
	nand3_1 U10715( .A(n8888), .B(n5900), .C(n8169), .Y(n8082) );
	nor2_1 U10716( .A(n6292), .B(n9283), .Y(n10072) );
	inv_1 U10717( .A(n10754), .Y(n9283) );
	o21ai_0 U10718( .A1(n6237), .A2(n9631), .B1(n10074), .Y(n4881) );
	mux2i_1 U10719( .A0(n10075), .A1(n10076), .S(n10077), .Y(n10074) );
	nor2_1 U10720( .A(n6353), .B(n10078), .Y(n10076) );
	and2_0 U10721( .A(n10078), .B(n7237), .X(n10075) );
	inv_1 U10722( .A(n10399), .Y(n9631) );
	o21ai_0 U10723( .A1(n6237), .A2(n6809), .B1(n10079), .Y(n4880) );
	mux2i_1 U10724( .A0(n10080), .A1(n6259), .S(n9023), .Y(n10079) );
	nor2_1 U10725( .A(n6680), .B(n6994), .Y(n9023) );
	nand2_1 U10726( .A(n10208), .B(n9600), .Y(n6680) );
	nor2_1 U10727( .A(n6292), .B(n9158), .Y(n10080) );
	inv_1 U10728( .A(n10808), .Y(n9158) );
	inv_1 U10729( .A(n10816), .Y(n6809) );
	o22ai_1 U10730( .A1(n6210), .A2(n10081), .B1(n10082), .B2(n6297), .Y(n4879) );
	nor3_1 U10731( .A(n10588), .B(n11895), .C(n11974), .Y(n10082) );
	o211ai_1 U10732( .A1(n6203), .A2(n8831), .B1(n8232), .C1(n10083), .Y(n4878) );
	mux2i_1 U10733( .A0(n10084), .A1(n10085), .S(n8818), .Y(n10083) );
	inv_1 U10734( .A(n10162), .Y(n8818) );
	nor2_1 U10735( .A(n6352), .B(n9982), .Y(n10085) );
	and2_0 U10736( .A(n9982), .B(n6345), .X(n10084) );
	nand2_1 U10737( .A(n8318), .B(n10328), .Y(n9982) );
	nor2_1 U10738( .A(n6647), .B(n6645), .Y(n8318) );
	nand2_1 U10739( .A(n10182), .B(n10362), .Y(n6645) );
	inv_1 U10740( .A(n10356), .Y(n6647) );
	nand2_1 U10741( .A(n6338), .B(n7207), .Y(n8232) );
	inv_1 U10742( .A(n10291), .Y(n7207) );
	inv_1 U10743( .A(n10328), .Y(n8831) );
	o221ai_1 U10744( .A1(n10086), .A2(n5966), .B1(n10337), .B2(n7794), .C1( n10087), .Y(n4877) );
	mux2i_1 U10745( .A0(n10088), .A1(n10089), .S(n7793), .Y(n10087) );
	nor4_1 U10746( .A(n7954), .B(n10090), .C(n6588), .D(n6744), .Y(n10089) );
	or2_0 U10747( .A(n6973), .B(n11962), .X(n6744) );
	inv_1 U10748( .A(n10337), .Y(n6588) );
	nand2_1 U10749( .A(n6224), .B(n7794), .Y(n10088) );
	inv_1 U10750( .A(n6591), .Y(n7794) );
	nor3_1 U10751( .A(n7954), .B(n7657), .C(n10090), .Y(n6591) );
	a211oi_1 U10752( .A1(n6329), .A2(n10090), .B1(n6746), .C1(n7358), .Y(n10086) );
	nor2_1 U10753( .A(n6292), .B(n7795), .Y(n7358) );
	inv_1 U10754( .A(n7954), .Y(n7795) );
	o211ai_1 U10755( .A1(n9740), .A2(n10091), .B1(n10152), .C1(n9741), .Y(n7954) );
	nor2_1 U10756( .A(n6292), .B(n9390), .Y(n6746) );
	o21ai_0 U10757( .A1(n6237), .A2(n7702), .B1(n10092), .Y(n4876) );
	mux2i_1 U10758( .A0(n10093), .A1(n6259), .S(n10094), .Y(n10092) );
	nor2_1 U10759( .A(n6668), .B(n7903), .Y(n10094) );
	nand3_1 U10760( .A(n8020), .B(n5899), .C(n8185), .Y(n7903) );
	inv_1 U10761( .A(n9056), .Y(n6668) );
	nor2_1 U10762( .A(n9618), .B(n10203), .Y(n9056) );
	nor2_1 U10763( .A(n6292), .B(n9494), .Y(n10093) );
	inv_1 U10764( .A(n10778), .Y(n9494) );
	o21ai_0 U10765( .A1(n6237), .A2(n8323), .B1(n10095), .Y(n4875) );
	mux2i_1 U10766( .A0(n10096), .A1(n10097), .S(n10098), .Y(n10095) );
	nor2_1 U10767( .A(n10410), .B(n6365), .Y(n10097) );
	nor2_1 U10768( .A(n8300), .B(n8294), .Y(n10096) );
	inv_1 U10769( .A(n10410), .Y(n8294) );
	o221ai_1 U10770( .A1(n7834), .A2(n6753), .B1(n6213), .B2(n5862), .C1(n10099), .Y(n4874) );
	a21oi_1 U10771( .A1(n6757), .A2(n10171), .B1(n6758), .Y(n10099) );
	nor3_1 U10772( .A(n7657), .B(n7833), .C(n7835), .Y(n6758) );
	nor2_1 U10773( .A(n7833), .B(n6301), .Y(n6757) );
	inv_1 U10774( .A(n7836), .Y(n6753) );
	nor2_1 U10775( .A(n6281), .B(n8506), .Y(n7836) );
	inv_1 U10776( .A(n7833), .Y(n8506) );
	o221ai_1 U10777( .A1(n7182), .A2(n10100), .B1(n6213), .B2(n10101), .C1( n9347), .Y(n4873) );
	nand3_1 U10778( .A(n10685), .B(n6378), .C(n7502), .Y(n9347) );
	inv_1 U10779( .A(n10685), .Y(n10101) );
	inv_1 U10780( .A(n10643), .Y(n10100) );
	or2_0 U10781( .A(n6314), .B(n7502), .X(n7182) );
	nor2_1 U10782( .A(n6704), .B(n8622), .Y(n7502) );
	nand3_1 U10783( .A(g25114), .B(g25219), .C(g17577), .Y(n6704) );
	nor2_1 U10784( .A(n6290), .B(n10102), .Y(n4872) );
	o22ai_1 U10785( .A1(n10103), .A2(n8048), .B1(n10104), .B2(n10105), .Y(n4871) );
	nor2_1 U10786( .A(n10106), .B(n6437), .Y(n10104) );
	o21ai_0 U10787( .A1(n6237), .A2(n8398), .B1(n10107), .Y(n4870) );
	mux2i_1 U10788( .A0(n9261), .A1(n10108), .S(n10109), .Y(n10107) );
	nor2_1 U10789( .A(n10110), .B(n10111), .Y(n10108) );
	inv_1 U10790( .A(n9262), .Y(n10111) );
	nor2_1 U10791( .A(n8393), .B(n6301), .Y(n9262) );
	inv_1 U10792( .A(n8388), .Y(n9261) );
	nand2_1 U10793( .A(n6338), .B(n8393), .Y(n8388) );
	inv_1 U10794( .A(n10414), .Y(n8398) );
	o21ai_0 U10795( .A1(n6238), .A2(n10112), .B1(n10113), .Y(n4869) );
	mux2i_1 U10796( .A0(n10114), .A1(n10115), .S(n6910), .Y(n10113) );
	nor2_1 U10797( .A(n6353), .B(n10116), .Y(n10115) );
	and2_0 U10798( .A(n10116), .B(n6344), .X(n10114) );
	nand3_1 U10799( .A(n7767), .B(n6552), .C(n10913), .Y(n10116) );
	nor3_1 U10800( .A(n6554), .B(n10441), .C(n6550), .Y(n7767) );
	inv_1 U10801( .A(n10913), .Y(n10112) );
	nor3_1 U10802( .A(n10117), .B(n6350), .C(n10118), .Y(n4868) );
	a21oi_1 U10803( .A1(n10850), .A2(n9735), .B1(n7257), .Y(n10118) );
	nor2_1 U10804( .A(n6934), .B(n9282), .Y(n9735) );
	nor3_1 U10805( .A(n9734), .B(n7259), .C(n9282), .Y(n10117) );
	inv_1 U10806( .A(n10850), .Y(n9734) );
	o22ai_1 U10807( .A1(n9069), .A2(n6630), .B1(n8886), .B2(n6632), .Y(n4867) );
	o21ai_0 U10808( .A1(n7776), .A2(n6934), .B1(n6383), .Y(n6632) );
	inv_1 U10809( .A(n10119), .Y(n7776) );
	nand2_1 U10810( .A(n6338), .B(n10119), .Y(n6630) );
	nand2_1 U10811( .A(n10120), .B(n7772), .Y(n10119) );
	mux2i_1 U10812( .A0(n10121), .A1(n10122), .S(n7043), .Y(n10120) );
	nand3_1 U10813( .A(n6811), .B(n7545), .C(n10168), .Y(n10122) );
	inv_1 U10814( .A(n10442), .Y(n7545) );
	inv_1 U10815( .A(n10421), .Y(n6811) );
	o21ai_0 U10816( .A1(n6238), .A2(n6503), .B1(n10123), .Y(n4866) );
	mux2i_1 U10817( .A0(n10124), .A1(n6259), .S(n10125), .Y(n10123) );
	nor2_1 U10818( .A(n6502), .B(n8483), .Y(n10125) );
	inv_1 U10819( .A(n9802), .Y(n6502) );
	nor2_1 U10820( .A(n6566), .B(n10201), .Y(n9802) );
	nor2_1 U10821( .A(n6289), .B(n5937), .Y(n10124) );
	inv_1 U10822( .A(n10833), .Y(n6503) );
	o221ai_1 U10823( .A1(n10126), .A2(n9963), .B1(n6214), .B2(n5884), .C1( n10127), .Y(n4865) );
	nand3_1 U10824( .A(n6341), .B(n7098), .C(n10472), .Y(n10127) );
	inv_1 U10825( .A(n9816), .Y(n9963) );
	nor2_1 U10826( .A(n6405), .B(n6934), .Y(n9816) );
	inv_1 U10827( .A(n88), .Y(n6405) );
	nor2_1 U10828( .A(n7098), .B(n6366), .Y(n88) );
	o32ai_1 U10829( .A1(n5907), .A2(n10128), .A3(n6312), .B1(n10129), .B2(n9545), .Y(n4864) );
	nor2_1 U10830( .A(n10130), .B(n6437), .Y(n10129) );
	nor4_1 U10831( .A(n11914), .B(n6367), .C(n9438), .D(n9544), .Y(n10130) );
	a21oi_1 U10832( .A1(n10131), .A2(n9545), .B1(n9544), .Y(n10128) );
	o21ai_0 U10833( .A1(n10560), .A2(n9438), .B1(n10132), .Y(n9544) );
	inv_1 U10834( .A(n10304), .Y(n9545) );
	nor2_1 U10835( .A(n5875), .B(n10069), .Y(n4863) );
	o22ai_1 U10836( .A1(n6304), .A2(n10133), .B1(n6194), .B2(n5865), .Y(n4862) );
	and3_1 U10837( .A(n6346), .B(n10134), .C(n10135), .X(n4861) );
	o22ai_1 U10838( .A1(n6211), .A2(n10136), .B1(n10137), .B2(n6298), .Y(n4860) );
	nor2_1 U10839( .A(g933), .B(n10455), .Y(n10137) );
	o32ai_1 U10840( .A1(n8384), .A2(n6348), .A3(n8383), .B1(n6476), .B2(n8673), .Y(n4859) );
	nand2_1 U10841( .A(n8383), .B(n6376), .Y(n8673) );
	inv_1 U10842( .A(n10316), .Y(n6476) );
	nor2_1 U10843( .A(n6934), .B(n8385), .Y(n8383) );
	inv_1 U10844( .A(n10856), .Y(n8384) );
	o22ai_1 U10845( .A1(n6304), .A2(n9515), .B1(n6194), .B2(n6083), .Y(n4858) );
	inv_1 U10846( .A(g6748), .Y(n9515) );
	nor2_1 U10847( .A(n10276), .B(n6479), .Y(n4857) );
	or3_1 U10848( .A(n9983), .B(n10158), .C(n6306), .X(n6479) );
	o21ai_0 U10849( .A1(n6238), .A2(n8609), .B1(n10138), .Y(n4856) );
	mux2i_1 U10850( .A0(n10139), .A1(n10140), .S(n9610), .Y(n10138) );
	and2_0 U10851( .A(n10392), .B(n8608), .X(n9610) );
	and2_0 U10852( .A(n10398), .B(n8458), .X(n8608) );
	nor2_1 U10853( .A(n10141), .B(n8454), .Y(n8458) );
	nor2_1 U10854( .A(n10383), .B(n6366), .Y(n10140) );
	nor2_1 U10855( .A(n7108), .B(n8367), .Y(n10139) );
	inv_1 U10856( .A(n10392), .Y(n8609) );
	o32ai_1 U10857( .A1(n10142), .A2(n6348), .A3(n6934), .B1(n6201), .B2(n10109), .Y(n4855) );
	mux2i_1 U10858( .A0(n10143), .A1(n10192), .S(n8393), .Y(n10142) );
	a21oi_1 U10859( .A1(n10047), .A2(n10144), .B1(n10110), .Y(n10143) );
	and2_0 U10860( .A(n7049), .B(n9175), .X(n10110) );
	and3_1 U10861( .A(n10255), .B(n9390), .C(n11769), .X(n9175) );
	inv_1 U10862( .A(n8397), .Y(n10144) );
	nor2_1 U10863( .A(n10109), .B(n10192), .Y(n8397) );
	inv_1 U10864( .A(n8394), .Y(n10047) );
	nor2_1 U10865( .A(n10145), .B(n10366), .Y(n8394) );
	o22ai_1 U10866( .A1(n6211), .A2(n5952), .B1(n10146), .B2(n6298), .Y(n4854) );
	a22oi_1 U10867( .A1(n10147), .A2(n8587), .B1(n10148), .B2(n8586), .Y(n10146) );
	xor2_1 U10868( .A(g115), .B(n9784), .X(n10148) );
	mux2i_1 U10869( .A0(g114), .A1(g116), .S(n10698), .Y(n9784) );
	inv_1 U10870( .A(n10465), .Y(n8587) );
	xor2_1 U10871( .A(g126), .B(n7123), .X(n10147) );
	mux2i_1 U10872( .A0(g120), .A1(g124), .S(n10465), .Y(n7123) );
	o22ai_1 U10873( .A1(n9566), .A2(n6564), .B1(n10149), .B2(n7618), .Y(n4853) );
	a21oi_1 U10874( .A1(n10150), .A2(n7616), .B1(n6437), .Y(n10149) );
	and2_0 U10875( .A(n10361), .B(n6565), .X(n7616) );
	nor2_1 U10876( .A(n6353), .B(n7617), .Y(n10150) );
	or2_0 U10877( .A(n7617), .B(n6310), .X(n6564) );
	nand2_1 U10878( .A(n8342), .B(n9568), .Y(n7617) );
	a21oi_1 U10879( .A1(n6198), .A2(n10892), .B1(n8282), .Y(n4852) );
	inv_1 U10880( .A(n10180), .Y(n8282) );
	nand2_1 U10881( .A(n10940), .B(n6370), .Y(n10892) );
	xnor2_1 U10882( .A(n11940), .B(n8283), .Y(n10940) );
	inv_1 U10883( .A(n9199), .Y(n8283) );
	nor2_1 U10884( .A(n8285), .B(n9195), .Y(n9199) );
	o21ai_0 U10885( .A1(n6238), .A2(n10941), .B1(n10942), .Y(n4851) );
	mux2i_1 U10886( .A0(n10943), .A1(n10944), .S(n7860), .Y(n10942) );
	nor2_1 U10887( .A(n10941), .B(n10945), .Y(n7860) );
	nor3_1 U10888( .A(n7861), .B(n10439), .C(n7862), .Y(n10944) );
	inv_1 U10889( .A(n10946), .Y(n7862) );
	nand2_1 U10890( .A(n10340), .B(n6375), .Y(n7861) );
	nor2_1 U10891( .A(n7855), .B(n7863), .Y(n10943) );
	o211ai_1 U10892( .A1(n10946), .A2(n10945), .B1(n6332), .C1(n10340), .Y( n7863) );
	nand4_1 U10893( .A(n10947), .B(n10857), .C(n10948), .D(n10949), .Y(n10946) );
	nor3_1 U10894( .A(n7060), .B(n11789), .C(n10449), .Y(n10949) );
	inv_1 U10895( .A(n10205), .Y(n7060) );
	xnor2_1 U10896( .A(n10220), .B(n10426), .Y(n10948) );
	xnor2_1 U10897( .A(n11966), .B(n10358), .Y(n10947) );
	inv_1 U10898( .A(n10439), .Y(n7855) );
	inv_1 U10899( .A(n10357), .Y(n10941) );
	o32ai_1 U10900( .A1(n10950), .A2(n10263), .A3(n7893), .B1(n7887), .B2(n8591), .Y(n4850) );
	nand2_1 U10901( .A(n8593), .B(n6337), .Y(n8591) );
	nor2_1 U10902( .A(n7891), .B(n8885), .Y(n7893) );
	o21ai_0 U10903( .A1(n10242), .A2(n9235), .B1(n6341), .Y(n10950) );
	nor2_1 U10904( .A(n10253), .B(n8593), .Y(n9235) );
	o21ai_0 U10905( .A1(n6238), .A2(n10951), .B1(n10952), .Y(n4849) );
	mux2i_1 U10906( .A0(n10953), .A1(n6259), .S(n10954), .Y(n10952) );
	nor2_1 U10907( .A(n8941), .B(n8949), .Y(n10954) );
	nor2_1 U10908( .A(n6291), .B(n6010), .Y(n10953) );
	nor2_1 U10909( .A(n10955), .B(n8761), .Y(n4848) );
	o21ai_0 U10910( .A1(n6934), .A2(n8352), .B1(n6383), .Y(n8761) );
	o21ai_0 U10911( .A1(n6238), .A2(n6053), .B1(n10956), .Y(n4847) );
	mux2i_1 U10912( .A0(n10957), .A1(n10958), .S(n10959), .Y(n10956) );
	nor2_1 U10913( .A(n10562), .B(n6366), .Y(n10958) );
	nor2_1 U10914( .A(n8486), .B(n10960), .Y(n10957) );
	o21ai_0 U10915( .A1(n6238), .A2(n6010), .B1(n10961), .Y(n4846) );
	mux2i_1 U10916( .A0(n10962), .A1(n6259), .S(n10963), .Y(n10961) );
	nor2_1 U10917( .A(n7072), .B(n8949), .Y(n10963) );
	nor2_1 U10918( .A(n6291), .B(n6011), .Y(n10962) );
	o32ai_1 U10919( .A1(n8887), .A2(n10154), .A3(n6628), .B1(n6201), .B2(n5900), .Y(n4845) );
	nand2_1 U10920( .A(n11972), .B(n10271), .Y(n6628) );
	inv_1 U10921( .A(n10964), .Y(n8887) );
	o221ai_1 U10922( .A1(n7723), .A2(n8551), .B1(n6214), .B2(n5965), .C1(n10965), .Y(n4844) );
	a21oi_1 U10923( .A1(n7158), .A2(n10175), .B1(n8752), .Y(n10965) );
	nor3_1 U10924( .A(n7222), .B(n7657), .C(n7724), .Y(n8752) );
	nand2_1 U10925( .A(n11962), .B(n10966), .Y(n7657) );
	inv_1 U10926( .A(n6973), .Y(n10966) );
	nand2_1 U10927( .A(n6917), .B(n6372), .Y(n6973) );
	nor2_1 U10928( .A(n7222), .B(n6301), .Y(n7158) );
	inv_1 U10929( .A(n7161), .Y(n8551) );
	nor2_1 U10930( .A(n6291), .B(n7220), .Y(n7161) );
	inv_1 U10931( .A(n7222), .Y(n7220) );
	o21ai_0 U10932( .A1(n6238), .A2(n5929), .B1(n10967), .Y(n4843) );
	mux2i_1 U10933( .A0(n10968), .A1(n6260), .S(n10969), .Y(n10967) );
	nor2_1 U10934( .A(n7015), .B(n7321), .Y(n10969) );
	inv_1 U10935( .A(n9986), .Y(n7015) );
	nor2_1 U10936( .A(n8745), .B(n10209), .Y(n9986) );
	nor2_1 U10937( .A(n6291), .B(n8645), .Y(n10968) );
	inv_1 U10938( .A(n10822), .Y(n8645) );
	o21ai_0 U10939( .A1(n6238), .A2(n8875), .B1(n10970), .Y(n4842) );
	mux2i_1 U10940( .A0(n10971), .A1(n6260), .S(n10972), .Y(n10970) );
	nor2_1 U10941( .A(n8614), .B(n8139), .Y(n10972) );
	nand2_1 U10942( .A(n8993), .B(n8921), .Y(n8139) );
	nor2_1 U10943( .A(n6291), .B(n6785), .Y(n10971) );
	nor2_1 U10944( .A(n10973), .B(n10069), .Y(n4841) );
	o21ai_0 U10945( .A1(n6934), .A2(n8107), .B1(n6382), .Y(n10069) );
	nand3_1 U10946( .A(n11777), .B(n9390), .C(n10974), .Y(n8107) );
	o32ai_1 U10947( .A1(n6550), .A2(n7572), .A3(n6312), .B1(n7573), .B2(n7571), .Y(n4840) );
	inv_1 U10948( .A(n10441), .Y(n7571) );
	a21oi_1 U10949( .A1(n6378), .A2(n7572), .B1(n6437), .Y(n7573) );
	nor3_1 U10950( .A(n10248), .B(n11957), .C(n6554), .Y(n7572) );
	inv_1 U10951( .A(g13259), .Y(n6554) );
	inv_1 U10952( .A(n10431), .Y(n6550) );
	o22ai_1 U10953( .A1(n6211), .A2(n6523), .B1(n6347), .B2(n8655), .Y(n4839) );
	nand3_1 U10954( .A(n10921), .B(n10294), .C(g8719), .Y(n8655) );
	o22ai_1 U10955( .A1(n6210), .A2(n10975), .B1(n10976), .B2(n6298), .Y(n4838) );
	nor4_1 U10956( .A(n10977), .B(n10978), .C(n9927), .D(n10979), .Y(n10976) );
	or2_0 U10957( .A(n9550), .B(n10980), .X(n10979) );
	or3_1 U10958( .A(n7299), .B(n6472), .C(n7298), .X(n10978) );
	nand4_1 U10959( .A(n10981), .B(n6873), .C(n8540), .D(n10982), .Y(n10977) );
	nor3_1 U10960( .A(n10211), .B(n10657), .C(n10538), .Y(n10982) );
	o22ai_1 U10961( .A1(n8008), .A2(n10983), .B1(n10984), .B2(n8010), .Y(n4837) );
	inv_1 U10962( .A(n10450), .Y(n8010) );
	a21oi_1 U10963( .A1(n4753), .A2(n8008), .B1(n6437), .Y(n10984) );
	inv_1 U10964( .A(n85), .Y(n10983) );
	nor2_1 U10965( .A(n8300), .B(n10450), .Y(n85) );
	nand2_1 U10966( .A(g12919), .B(n6337), .Y(n8300) );
	inv_1 U10967( .A(n10389), .Y(n8008) );
	o21ai_0 U10968( .A1(n6238), .A2(n7027), .B1(n10985), .Y(n4836) );
	mux2i_1 U10969( .A0(n10986), .A1(n6260), .S(n9211), .Y(n10985) );
	nor2_1 U10970( .A(n6905), .B(n7228), .Y(n9211) );
	nand2_1 U10971( .A(n10207), .B(n9805), .Y(n6905) );
	nor2_1 U10972( .A(n6291), .B(n9892), .Y(n10986) );
	inv_1 U10973( .A(n10769), .Y(n9892) );
	inv_1 U10974( .A(n10777), .Y(n7027) );
	o21ai_0 U10975( .A1(n6238), .A2(n7497), .B1(n10987), .Y(n4835) );
	mux2i_1 U10976( .A0(n10988), .A1(n6260), .S(n10989), .Y(n10987) );
	nor2_1 U10977( .A(n7496), .B(n8169), .Y(n10989) );
	nor2_1 U10978( .A(n6291), .B(n10070), .Y(n10988) );
	inv_1 U10979( .A(n10753), .Y(n10070) );
	inv_1 U10980( .A(n10757), .Y(n7497) );
	o21ai_0 U10981( .A1(n6238), .A2(n6996), .B1(n10990), .Y(n4834) );
	mux2i_1 U10982( .A0(n10991), .A1(n6260), .S(n10992), .Y(n10990) );
	nor2_1 U10983( .A(n7875), .B(n6681), .Y(n10992) );
	nand3_1 U10984( .A(n8558), .B(n5901), .C(n6994), .Y(n6681) );
	inv_1 U10985( .A(n10275), .Y(n8558) );
	nor2_1 U10986( .A(n6291), .B(n8162), .Y(n10991) );
	inv_1 U10987( .A(n10806), .Y(n8162) );
	inv_1 U10988( .A(n10805), .Y(n6996) );
	mux2i_1 U10989( .A0(n10993), .A1(n10994), .S(n10718), .Y(n4833) );
	a21oi_1 U10990( .A1(n6378), .A2(n7732), .B1(n6437), .Y(n10994) );
	nand2_1 U10991( .A(n10215), .B(n6336), .Y(n10993) );
	o21ai_0 U10992( .A1(n6238), .A2(n7998), .B1(n10995), .Y(n4832) );
	mux2i_1 U10993( .A0(n10996), .A1(n10997), .S(n8454), .Y(n10995) );
	inv_1 U10994( .A(n10527), .Y(n8454) );
	nor2_1 U10995( .A(n6353), .B(n10141), .Y(n10997) );
	nor2_1 U10996( .A(n10998), .B(n7108), .Y(n10996) );
	inv_1 U10997( .A(n10141), .Y(n10998) );
	nand2_1 U10998( .A(n10528), .B(n7997), .Y(n10141) );
	and2_0 U10999( .A(n8278), .B(n10401), .X(n7997) );
	and2_0 U11000( .A(n10394), .B(n7592), .X(n8278) );
	and2_0 U11001( .A(n10067), .B(n10396), .X(n7592) );
	and2_0 U11002( .A(n10390), .B(n7107), .X(n10067) );
	and2_0 U11003( .A(n8313), .B(n10531), .X(n7107) );
	and2_0 U11004( .A(n10532), .B(n9104), .X(n8313) );
	and2_0 U11005( .A(n10533), .B(n9229), .X(n9104) );
	nor2_1 U11006( .A(n8677), .B(n8678), .Y(n9229) );
	nand3_1 U11007( .A(n10999), .B(n11000), .C(n11857), .Y(n8678) );
	inv_1 U11008( .A(n10534), .Y(n8677) );
	inv_1 U11009( .A(n10528), .Y(n7998) );
	o22ai_1 U11010( .A1(n6209), .A2(n11001), .B1(n7108), .B2(n11002), .Y(n4831) );
	o21ai_0 U11011( .A1(n8372), .A2(n9607), .B1(n11003), .Y(n11002) );
	xnor2_1 U11012( .A(n5888), .B(n10999), .Y(n11003) );
	a21oi_1 U11013( .A1(n11004), .A2(g12368), .B1(n11005), .Y(n10999) );
	nand2_1 U11014( .A(n6339), .B(n11000), .Y(n7108) );
	nand2_1 U11015( .A(g9048), .B(n11001), .Y(n11000) );
	inv_1 U11016( .A(n10662), .Y(n11001) );
	o32ai_1 U11017( .A1(n7258), .A2(n6348), .A3(n6545), .B1(n6546), .B2(n8641), .Y(n4830) );
	inv_1 U11018( .A(n10314), .Y(n8641) );
	nand2_1 U11019( .A(n6545), .B(n6379), .Y(n6546) );
	nor2_1 U11020( .A(n6934), .B(n7010), .Y(n6545) );
	inv_1 U11021( .A(n10854), .Y(n7258) );
	o21ai_0 U11022( .A1(n6238), .A2(n11006), .B1(n11007), .Y(n4829) );
	mux2i_1 U11023( .A0(n11008), .A1(n6260), .S(n9057), .Y(n11007) );
	nor2_1 U11024( .A(n8099), .B(n8185), .Y(n9057) );
	nor2_1 U11025( .A(n6291), .B(n7702), .Y(n11008) );
	inv_1 U11026( .A(n10782), .Y(n7702) );
	o21ai_0 U11027( .A1(n6238), .A2(n10960), .B1(n11009), .Y(n4828) );
	mux2i_1 U11028( .A0(n11010), .A1(n11011), .S(n8754), .Y(n11009) );
	inv_1 U11029( .A(n10540), .Y(n8754) );
	nor2_1 U11030( .A(n6353), .B(n9822), .Y(n11011) );
	nor2_1 U11031( .A(n11012), .B(n8486), .Y(n11010) );
	nand2_1 U11032( .A(n8634), .B(n6336), .Y(n8486) );
	inv_1 U11033( .A(n9822), .Y(n11012) );
	nand2_1 U11034( .A(n10562), .B(n10959), .Y(n9822) );
	and3_1 U11035( .A(n11819), .B(n8634), .C(n10924), .X(n10959) );
	and3_1 U11036( .A(n10135), .B(n9654), .C(n11013), .X(n8634) );
	a21oi_1 U11037( .A1(n10895), .A2(n10134), .B1(n7043), .Y(n11013) );
	inv_1 U11038( .A(n10267), .Y(n7043) );
	nand4_1 U11039( .A(n10458), .B(n10463), .C(n10218), .D(n11014), .Y(n10134) );
	nor4_1 U11040( .A(n10459), .B(n10302), .C(n10187), .D(n7367), .Y(n11014) );
	o21ai_0 U11041( .A1(n11015), .A2(n11016), .B1(n8485), .Y(n10135) );
	inv_1 U11042( .A(n10895), .Y(n8485) );
	nand3_1 U11043( .A(n10302), .B(n10459), .C(n10187), .Y(n11016) );
	nand4_1 U11044( .A(n7367), .B(n7938), .C(n7934), .D(n7935), .Y(n11015) );
	inv_1 U11045( .A(n10463), .Y(n7935) );
	inv_1 U11046( .A(n10178), .Y(n7367) );
	inv_1 U11047( .A(n10562), .Y(n10960) );
	o21ai_0 U11048( .A1(n6238), .A2(n6012), .B1(n11017), .Y(n4827) );
	mux2i_1 U11049( .A0(n11018), .A1(n6260), .S(n11019), .Y(n11017) );
	nor2_1 U11050( .A(n8191), .B(n9287), .Y(n11019) );
	nor2_1 U11051( .A(n6291), .B(n6013), .Y(n11018) );
	nor2_1 U11052( .A(n6291), .B(n11020), .Y(n4826) );
	o22ai_1 U11053( .A1(n6209), .A2(n11021), .B1(n11022), .B2(n6297), .Y(n4825) );
	and2_0 U11054( .A(g4531), .B(n10380), .X(n11022) );
	inv_1 U11055( .A(n10880), .Y(n11021) );
	o211ai_1 U11056( .A1(n11023), .A2(n11024), .B1(n11025), .C1(n8144), .Y( n4824) );
	nand3_1 U11057( .A(n11026), .B(n6330), .C(n11879), .Y(n8144) );
	nand3_1 U11058( .A(n11916), .B(n11027), .C(n8146), .Y(n11025) );
	nor2_1 U11059( .A(n6291), .B(n11026), .Y(n8146) );
	inv_1 U11060( .A(n7197), .Y(n11027) );
	inv_1 U11061( .A(n10596), .Y(n11024) );
	a21oi_1 U11062( .A1(n8147), .A2(n7197), .B1(n6437), .Y(n11023) );
	nor2_1 U11063( .A(n9068), .B(n11028), .Y(n7197) );
	nor2_1 U11064( .A(n11026), .B(n6366), .Y(n8147) );
	nor3_1 U11065( .A(g8178), .B(n10600), .C(n9969), .Y(n11026) );
	o32ai_1 U11066( .A1(n6583), .A2(n6349), .A3(n7604), .B1(n7605), .B2(n8005), .Y(n4823) );
	inv_1 U11067( .A(n10730), .Y(n8005) );
	nand2_1 U11068( .A(n7604), .B(n6379), .Y(n7605) );
	nor2_1 U11069( .A(n6934), .B(n6584), .Y(n7604) );
	nor3_1 U11070( .A(n10241), .B(n10262), .C(n6579), .Y(n6584) );
	inv_1 U11071( .A(n6582), .Y(n6579) );
	nand2_1 U11072( .A(n6585), .B(n9303), .Y(n6582) );
	o21ai_0 U11073( .A1(n11029), .A2(n11030), .B1(n10718), .Y(n9303) );
	nand2_1 U11074( .A(n6406), .B(n5884), .Y(n11030) );
	inv_1 U11075( .A(n9829), .Y(n6585) );
	o211ai_1 U11076( .A1(n10507), .A2(n7455), .B1(n11031), .C1(n11032), .Y( n9829) );
	nand3_1 U11077( .A(n10281), .B(n10167), .C(n10382), .Y(n11031) );
	inv_1 U11078( .A(n10481), .Y(n6583) );
	and2_0 U11079( .A(n6346), .B(n10889), .X(n4822) );
	o21ai_0 U11080( .A1(n6238), .A2(n10077), .B1(n11033), .Y(n4821) );
	mux2i_1 U11081( .A0(n11034), .A1(n11035), .S(n11036), .Y(n11033) );
	nor2_1 U11082( .A(n10391), .B(n6366), .Y(n11035) );
	nor2_1 U11083( .A(n11037), .B(n8048), .Y(n11034) );
	o22ai_1 U11084( .A1(n9940), .A2(n9958), .B1(n11038), .B2(n9959), .Y(n4820) );
	inv_1 U11085( .A(n10436), .Y(n9959) );
	a21oi_1 U11086( .A1(n6383), .A2(n9940), .B1(n6437), .Y(n11038) );
	inv_1 U11087( .A(n22), .Y(n9958) );
	inv_1 U11088( .A(n10317), .Y(n9940) );
	o21ai_0 U11089( .A1(n6239), .A2(n5930), .B1(n11039), .Y(n4819) );
	mux2i_1 U11090( .A0(n11040), .A1(n6260), .S(n11041), .Y(n11039) );
	nor2_1 U11091( .A(n7321), .B(n7965), .Y(n11041) );
	nand2_1 U11092( .A(n6480), .B(n8745), .Y(n7965) );
	inv_1 U11093( .A(n10209), .Y(n6480) );
	nand2_1 U11094( .A(n10276), .B(n11960), .Y(n7321) );
	nor2_1 U11095( .A(n6290), .B(n7961), .Y(n11040) );
	o21ai_0 U11096( .A1(n6239), .A2(n6014), .B1(n11042), .Y(n4818) );
	mux2i_1 U11097( .A0(n11043), .A1(n6260), .S(n11044), .Y(n11042) );
	nor2_1 U11098( .A(n6669), .B(n8099), .Y(n11044) );
	nor2_1 U11099( .A(n6290), .B(n6016), .Y(n11043) );
	o21ai_0 U11100( .A1(n6239), .A2(n5970), .B1(n11045), .Y(n4817) );
	mux2i_1 U11101( .A0(n11046), .A1(n11047), .S(n9540), .Y(n11045) );
	inv_1 U11102( .A(n10560), .Y(n9540) );
	nor2_1 U11103( .A(n8520), .B(n11048), .Y(n11047) );
	nand2_1 U11104( .A(n10131), .B(n6336), .Y(n8520) );
	nor2_1 U11105( .A(n10132), .B(n6301), .Y(n11046) );
	inv_1 U11106( .A(n11048), .Y(n10132) );
	o21ai_0 U11107( .A1(n11834), .A2(n9438), .B1(n9435), .Y(n11048) );
	a21oi_1 U11108( .A1(n8518), .A2(n10131), .B1(n8519), .Y(n9435) );
	inv_1 U11109( .A(n9438), .Y(n10131) );
	inv_1 U11110( .A(n10387), .Y(n8518) );
	nand3_1 U11111( .A(n9782), .B(n7971), .C(n11049), .Y(n9438) );
	mux2i_1 U11112( .A0(n11050), .A1(n11051), .S(n7424), .Y(n11049) );
	inv_1 U11113( .A(n10518), .Y(n7424) );
	nor2_1 U11114( .A(n11051), .B(n9783), .Y(n11050) );
	nand2_1 U11115( .A(n11834), .B(n10304), .Y(n9783) );
	inv_1 U11116( .A(n10557), .Y(n7971) );
	nand2_1 U11117( .A(n11939), .B(n11051), .Y(n9782) );
	o22ai_1 U11118( .A1(n6304), .A2(n9897), .B1(n6194), .B2(n6066), .Y(n4816) );
	mux2i_1 U11119( .A0(n11052), .A1(n11053), .S(n8614), .Y(n4815) );
	nand2_1 U11120( .A(n9462), .B(n10204), .Y(n11053) );
	a21oi_1 U11121( .A1(n8817), .A2(n9762), .B1(n6307), .Y(n9462) );
	a21oi_1 U11122( .A1(n7558), .A2(n8993), .B1(n6437), .Y(n11052) );
	inv_1 U11123( .A(n10204), .Y(n8993) );
	a21oi_1 U11124( .A1(n8817), .A2(n9762), .B1(n6368), .Y(n7558) );
	inv_1 U11125( .A(n9512), .Y(n9762) );
	o21ai_0 U11126( .A1(n6239), .A2(n5945), .B1(n7544), .Y(n4814) );
	inv_1 U11127( .A(n7513), .Y(n7544) );
	nor2_1 U11128( .A(n7512), .B(n6934), .Y(n7513) );
	nand2_1 U11129( .A(g12923), .B(n6374), .Y(n7512) );
	o22ai_1 U11130( .A1(n5908), .A2(n6202), .B1(n6300), .B2(n11054), .Y(n4813) );
	mux2i_1 U11131( .A0(n11055), .A1(n10422), .S(n6715), .Y(n11054) );
	nor2_1 U11132( .A(n10422), .B(n6711), .Y(n11055) );
	inv_1 U11133( .A(n10517), .Y(n6711) );
	o21ai_0 U11134( .A1(n6239), .A2(n6030), .B1(n11056), .Y(n4812) );
	mux2i_1 U11135( .A0(n11057), .A1(n7064), .S(n11058), .Y(n11056) );
	nor2_1 U11136( .A(n7883), .B(n9320), .Y(n11058) );
	inv_1 U11137( .A(n9961), .Y(n9320) );
	nor2_1 U11138( .A(n10250), .B(n7884), .Y(n9961) );
	inv_1 U11139( .A(n10239), .Y(n7883) );
	nor2_1 U11140( .A(n6285), .B(n6025), .Y(n11057) );
	and2_0 U11141( .A(n6345), .B(n10887), .X(n4811) );
	o22ai_1 U11142( .A1(n6209), .A2(n9569), .B1(n11059), .B2(n8467), .Y(n4810) );
	nand2_1 U11143( .A(n11060), .B(n8472), .Y(n8467) );
	nand2_1 U11144( .A(n10719), .B(n8871), .Y(n8472) );
	xnor2_1 U11145( .A(n10269), .B(n8871), .Y(n11059) );
	nor2_1 U11146( .A(n9568), .B(n9569), .Y(n8871) );
	nand3_1 U11147( .A(n10246), .B(n6565), .C(n10279), .Y(n9568) );
	nor2_1 U11148( .A(n6880), .B(n11061), .Y(n6565) );
	o22ai_1 U11149( .A1(n8220), .A2(n8218), .B1(n11062), .B2(n9454), .Y(n4809) );
	a21oi_1 U11150( .A1(n8221), .A2(n8220), .B1(n6437), .Y(n11062) );
	inv_1 U11151( .A(n8350), .Y(n8221) );
	nand3_1 U11152( .A(n8352), .B(n6377), .C(n9455), .Y(n8350) );
	o211ai_1 U11153( .A1(n8220), .A2(n11063), .B1(n8352), .C1(n6331), .Y(n8218) );
	nand3_1 U11154( .A(n11064), .B(n9390), .C(n11777), .Y(n8352) );
	inv_1 U11155( .A(n9455), .Y(n11063) );
	nor2_1 U11156( .A(n9365), .B(n9366), .Y(n9455) );
	o21ai_0 U11157( .A1(n6239), .A2(n6027), .B1(n11065), .Y(n4808) );
	mux2i_1 U11158( .A0(n11066), .A1(n6559), .S(n11067), .Y(n11065) );
	nor2_1 U11159( .A(n10287), .B(n8015), .Y(n11067) );
	inv_1 U11160( .A(n9474), .Y(n8015) );
	nor2_1 U11161( .A(n8734), .B(n8431), .Y(n9474) );
	nor2_1 U11162( .A(n8435), .B(n9007), .Y(n8431) );
	inv_1 U11163( .A(n11068), .Y(n9007) );
	o21ai_0 U11164( .A1(n9810), .A2(n11069), .B1(n10717), .Y(n11068) );
	nand2_1 U11165( .A(n6486), .B(n8723), .Y(n11069) );
	inv_1 U11166( .A(n10923), .Y(n8723) );
	inv_1 U11167( .A(n10247), .Y(n8734) );
	and2_0 U11168( .A(n6345), .B(n11070), .X(n6559) );
	o21ai_0 U11169( .A1(n10469), .A2(n8435), .B1(n8429), .Y(n11070) );
	o211ai_1 U11170( .A1(n10285), .A2(n9974), .B1(n8435), .C1(n9975), .Y(n8429) );
	o211ai_1 U11171( .A1(n10508), .A2(n6799), .B1(n11071), .C1(n9811), .Y(n8435) );
	nand3_1 U11172( .A(n10280), .B(n10166), .C(n10432), .Y(n11071) );
	nor2_1 U11173( .A(n6290), .B(n6026), .Y(n11066) );
	o21ai_0 U11174( .A1(n6239), .A2(n8930), .B1(n11072), .Y(n4807) );
	mux2i_1 U11175( .A0(n11073), .A1(n6260), .S(n11074), .Y(n11072) );
	nor2_1 U11176( .A(n7496), .B(n8191), .Y(n11074) );
	nand2_1 U11177( .A(n11972), .B(n8888), .Y(n8191) );
	inv_1 U11178( .A(n10271), .Y(n8888) );
	inv_1 U11179( .A(n8171), .Y(n7496) );
	nor2_1 U11180( .A(n9046), .B(n10206), .Y(n8171) );
	nor2_1 U11181( .A(n6290), .B(n5928), .Y(n11073) );
	inv_1 U11182( .A(n10755), .Y(n8930) );
	o21ai_0 U11183( .A1(n6239), .A2(n7466), .B1(n11075), .Y(n4806) );
	a22oi_1 U11184( .A1(n11076), .A2(n6835), .B1(n10902), .B2(n6831), .Y(n11075) );
	nor2_1 U11185( .A(n6290), .B(n9173), .Y(n6831) );
	inv_1 U11186( .A(n9063), .Y(n9173) );
	nor2_1 U11187( .A(n9063), .B(n6300), .Y(n6835) );
	nand2_1 U11188( .A(n10535), .B(n11077), .Y(n9063) );
	nand3_1 U11189( .A(n11905), .B(n8229), .C(n9388), .Y(n11077) );
	inv_1 U11190( .A(n9706), .Y(n9388) );
	nand4_1 U11191( .A(n10462), .B(n10289), .C(n11961), .D(n11078), .Y(n9706) );
	nor3_1 U11192( .A(n7822), .B(n10347), .C(n10277), .Y(n11078) );
	xnor2_1 U11193( .A(n11079), .B(n9178), .Y(n11076) );
	nand2_1 U11194( .A(n11080), .B(n11081), .Y(n9178) );
	mux2i_1 U11195( .A0(n11082), .A1(n11083), .S(n11084), .Y(n11081) );
	xnor2_1 U11196( .A(n7167), .B(g11388), .Y(n11084) );
	nand3_1 U11197( .A(n11085), .B(n11086), .C(n11087), .Y(n11083) );
	nand3_1 U11198( .A(g16627), .B(n10499), .C(n9066), .Y(n11087) );
	nand3_1 U11199( .A(g16744), .B(n11785), .C(n9065), .Y(n11086) );
	nand3_1 U11200( .A(g13926), .B(n11824), .C(n9067), .Y(n11085) );
	nand3_1 U11201( .A(n11088), .B(n11089), .C(n11090), .Y(n11082) );
	nand3_1 U11202( .A(n9064), .B(g16744), .C(n11850), .Y(n11090) );
	nand3_1 U11203( .A(n10829), .B(g16627), .C(n9067), .Y(n11089) );
	nand3_1 U11204( .A(n9066), .B(g13926), .C(n11875), .Y(n11088) );
	mux2_1 U11205( .A0(n11091), .A1(n11092), .S(n7167), .X(n11080) );
	a221oi_1 U11206( .A1(n9066), .A2(n11093), .B1(n9064), .B2(n11094), .C1( n11095), .Y(n11092) );
	o32ai_1 U11207( .A1(n11096), .A2(n5929), .A3(n11097), .B1(n11098), .B2( n11099), .Y(n11095) );
	a22oi_1 U11208( .A1(g16656), .A2(n10821), .B1(g16722), .B2(n10822), .Y( n11098) );
	inv_1 U11209( .A(n9067), .Y(n11097) );
	o22ai_1 U11210( .A1(n7747), .A2(n11100), .B1(n11101), .B2(n8937), .Y(n11094) );
	inv_1 U11211( .A(n10819), .Y(n8937) );
	inv_1 U11212( .A(n10820), .Y(n7747) );
	o22ai_1 U11213( .A1(n8649), .A2(n11102), .B1(n7017), .B2(n11103), .Y(n11093) );
	inv_1 U11214( .A(n10817), .Y(n7017) );
	inv_1 U11215( .A(n10818), .Y(n8649) );
	a221oi_1 U11216( .A1(n9067), .A2(n11104), .B1(n9064), .B2(n11105), .C1( n11106), .Y(n11091) );
	o32ai_1 U11217( .A1(n11096), .A2(n5930), .A3(n9174), .B1(n11107), .B2( n11099), .Y(n11106) );
	inv_1 U11218( .A(n9065), .Y(n11099) );
	nor2_1 U11219( .A(n6833), .B(n10196), .Y(n9065) );
	a22oi_1 U11220( .A1(n10825), .A2(g11388), .B1(g16924), .B2(n10826), .Y( n11107) );
	inv_1 U11221( .A(n9066), .Y(n9174) );
	nor2_1 U11222( .A(n11108), .B(n10370), .Y(n9066) );
	o22ai_1 U11223( .A1(n7961), .A2(n9761), .B1(n9176), .B2(n11109), .Y(n11105) );
	inv_1 U11224( .A(n10823), .Y(n9176) );
	inv_1 U11225( .A(g16722), .Y(n9761) );
	inv_1 U11226( .A(n10824), .Y(n7961) );
	o22ai_1 U11227( .A1(n7966), .A2(n11102), .B1(n8749), .B2(n11103), .Y(n11104) );
	inv_1 U11228( .A(n10827), .Y(n8749) );
	nor2_1 U11229( .A(n10370), .B(n10196), .Y(n9067) );
	nand2_1 U11230( .A(n10902), .B(n11110), .Y(n11079) );
	nand3_1 U11231( .A(n9064), .B(n10378), .C(g16656), .Y(n11110) );
	inv_1 U11232( .A(n10315), .Y(n7466) );
	o21ai_0 U11233( .A1(n6239), .A2(n6015), .B1(n11111), .Y(n4805) );
	mux2i_1 U11234( .A0(n11112), .A1(n6260), .S(n11113), .Y(n11111) );
	nor2_1 U11235( .A(n6888), .B(n8251), .Y(n11113) );
	nor2_1 U11236( .A(n6290), .B(n6423), .Y(n11112) );
	inv_1 U11237( .A(n10496), .Y(n6423) );
	o32ai_1 U11238( .A1(n8482), .A2(n10164), .A3(n6467), .B1(n6201), .B2(n7254), .Y(n4804) );
	inv_1 U11239( .A(n10574), .Y(n7254) );
	nand2_1 U11240( .A(n10574), .B(n10295), .Y(n6467) );
	inv_1 U11241( .A(n9203), .Y(n8482) );
	a21oi_1 U11242( .A1(n9027), .A2(n9119), .B1(n6368), .Y(n9203) );
	inv_1 U11243( .A(n9323), .Y(n9027) );
	nor2_1 U11244( .A(n6353), .B(n10050), .Y(n4803) );
	inv_1 U11245( .A(g17743), .Y(n10050) );
	o21ai_0 U11246( .A1(n7208), .A2(n7909), .B1(n11114), .Y(n4802) );
	mux2i_1 U11247( .A0(n11115), .A1(n11116), .S(n10640), .Y(n11114) );
	nand2_1 U11248( .A(n6221), .B(n8208), .Y(n11116) );
	nand3_1 U11249( .A(n7214), .B(n6378), .C(n10502), .Y(n8208) );
	nor2_1 U11250( .A(n10502), .B(n7215), .Y(n11115) );
	nand2_1 U11251( .A(n7214), .B(n6336), .Y(n7215) );
	inv_1 U11252( .A(n10866), .Y(n7909) );
	or2_0 U11253( .A(n6314), .B(n7214), .X(n7208) );
	nor4_1 U11254( .A(n9842), .B(n10051), .C(n11117), .D(n8393), .Y(n7214) );
	nand2_1 U11255( .A(n10198), .B(n11118), .Y(n8393) );
	nand3_1 U11256( .A(n11119), .B(n9838), .C(n11801), .Y(n11118) );
	inv_1 U11257( .A(n8396), .Y(n11117) );
	o21ai_0 U11258( .A1(n6239), .A2(n7708), .B1(n11120), .Y(n4801) );
	mux2i_1 U11259( .A0(n11121), .A1(n6260), .S(n11122), .Y(n11120) );
	nor2_1 U11260( .A(n6669), .B(n8250), .Y(n11122) );
	nand2_1 U11261( .A(n8186), .B(n9618), .Y(n8250) );
	inv_1 U11262( .A(n10203), .Y(n8186) );
	nand2_1 U11263( .A(n11907), .B(n8020), .Y(n6669) );
	inv_1 U11264( .A(n10273), .Y(n8020) );
	nor2_1 U11265( .A(n6290), .B(n5938), .Y(n11121) );
	inv_1 U11266( .A(n10787), .Y(n7708) );
	o21ai_0 U11267( .A1(n6239), .A2(n11037), .B1(n11123), .Y(n4800) );
	mux2i_1 U11268( .A0(n11124), .A1(n11125), .S(n11126), .Y(n11123) );
	nor2_1 U11269( .A(n10397), .B(n6365), .Y(n11125) );
	nor2_1 U11270( .A(n8510), .B(n8048), .Y(n11124) );
	inv_1 U11271( .A(n10391), .Y(n11037) );
	o21ai_0 U11272( .A1(n6239), .A2(n11127), .B1(n11128), .Y(n4799) );
	nand2_1 U11273( .A(g6744), .B(n6336), .Y(n11128) );
	o221ai_1 U11274( .A1(n11129), .A2(n6307), .B1(n6214), .B2(n7418), .C1( n11130), .Y(n4798) );
	or3_1 U11275( .A(n6369), .B(n10330), .C(n11131), .X(n11130) );
	inv_1 U11276( .A(n10199), .Y(n7418) );
	a21oi_1 U11277( .A1(n10330), .A2(n11131), .B1(n7416), .Y(n11129) );
	nor2_1 U11278( .A(n8194), .B(n11938), .Y(n7416) );
	inv_1 U11279( .A(n10501), .Y(n8194) );
	nand2_1 U11280( .A(n7419), .B(n10199), .Y(n11131) );
	a211oi_1 U11281( .A1(n7414), .A2(n9578), .B1(n9577), .C1(n9575), .Y(n7419) );
	inv_1 U11282( .A(n9579), .Y(n9575) );
	nor2_1 U11283( .A(n8525), .B(n10300), .Y(n9579) );
	inv_1 U11284( .A(n9375), .Y(n9577) );
	nor3_1 U11285( .A(n6523), .B(n10921), .C(n7379), .Y(n9375) );
	o221ai_1 U11286( .A1(n11132), .A2(n5869), .B1(n6214), .B2(n9077), .C1( n11133), .Y(n4797) );
	nand3_1 U11287( .A(n7628), .B(n11134), .C(n7626), .Y(n11133) );
	nor2_1 U11288( .A(n7633), .B(n6299), .Y(n7626) );
	xnor2_1 U11289( .A(n8680), .B(n10674), .Y(n11134) );
	inv_1 U11290( .A(n10726), .Y(n8680) );
	inv_1 U11291( .A(n10674), .Y(n9077) );
	a21oi_1 U11292( .A1(n6331), .A2(n9084), .B1(n7625), .Y(n11132) );
	nor2_1 U11293( .A(n6290), .B(n9083), .Y(n7625) );
	inv_1 U11294( .A(n7633), .Y(n9083) );
	o211ai_1 U11295( .A1(n9740), .A2(n9726), .B1(n9813), .C1(n8630), .Y(n7633) );
	inv_1 U11296( .A(n7628), .Y(n9084) );
	nor2_1 U11297( .A(n9042), .B(n11946), .Y(n7628) );
	o21ai_0 U11298( .A1(n6239), .A2(n6016), .B1(n11135), .Y(n4796) );
	mux2i_1 U11299( .A0(n11136), .A1(n6260), .S(n11137), .Y(n11135) );
	nor2_1 U11300( .A(n8099), .B(n8251), .Y(n11137) );
	nand2_1 U11301( .A(n10273), .B(n11907), .Y(n8251) );
	nand2_1 U11302( .A(n10203), .B(n9618), .Y(n8099) );
	nor2_1 U11303( .A(n6290), .B(n11006), .Y(n11136) );
	inv_1 U11304( .A(n10790), .Y(n11006) );
	o22ai_1 U11305( .A1(n6458), .A2(n8853), .B1(n11138), .B2(n11139), .Y(n4795) );
	inv_1 U11306( .A(n10920), .Y(n11139) );
	a21oi_1 U11307( .A1(n8854), .A2(n6458), .B1(n6437), .Y(n11138) );
	nor2_1 U11308( .A(n8473), .B(n11847), .Y(n8854) );
	inv_1 U11309( .A(n36), .Y(n8853) );
	o21ai_0 U11310( .A1(n6239), .A2(n5876), .B1(n11140), .Y(n4794) );
	mux2i_1 U11311( .A0(n6616), .A1(n11141), .S(n8180), .Y(n11140) );
	inv_1 U11312( .A(n10695), .Y(n8180) );
	inv_1 U11313( .A(n8572), .Y(n11141) );
	nand2_1 U11314( .A(n9208), .B(n6336), .Y(n8572) );
	nor2_1 U11315( .A(n6290), .B(n9208), .Y(n6616) );
	nor3_1 U11316( .A(n7723), .B(n7222), .C(n5895), .Y(n9208) );
	o211ai_1 U11317( .A1(n9740), .A2(n5885), .B1(n9813), .C1(n11142), .Y(n7222) );
	inv_1 U11318( .A(n10336), .Y(n7723) );
	o21ai_0 U11319( .A1(n6239), .A2(n6035), .B1(n11143), .Y(n4793) );
	mux2i_1 U11320( .A0(n11144), .A1(n7021), .S(n11145), .Y(n11143) );
	nor2_1 U11321( .A(n7450), .B(n9087), .Y(n11145) );
	inv_1 U11322( .A(n10243), .Y(n9087) );
	inv_1 U11323( .A(n9800), .Y(n7450) );
	nor2_1 U11324( .A(n10254), .B(n9243), .Y(n9800) );
	nor2_1 U11325( .A(n6287), .B(n6017), .Y(n11144) );
	a21oi_1 U11326( .A1(n6198), .A2(n11146), .B1(n5917), .Y(n4792) );
	or2_0 U11327( .A(n7166), .B(n6369), .X(n11146) );
	nor2_1 U11328( .A(n7167), .B(n11147), .Y(n7166) );
	and2_0 U11329( .A(g4571), .B(n6383), .X(n4791) );
	o221ai_1 U11330( .A1(n6036), .A2(n7814), .B1(n11148), .B2(n11149), .C1( n11150), .Y(n4790) );
	a22oi_1 U11331( .A1(n10546), .A2(n8240), .B1(n10334), .B2(n6437), .Y(n11150) );
	nor2_1 U11332( .A(n6288), .B(n6771), .Y(n8240) );
	inv_1 U11333( .A(n9075), .Y(n6771) );
	inv_1 U11334( .A(n7586), .Y(n11149) );
	nor2_1 U11335( .A(n9075), .B(n6299), .Y(n7586) );
	a221oi_1 U11336( .A1(n9074), .A2(n10722), .B1(n7921), .B2(n11786), .C1( n11151), .Y(n11148) );
	o32ai_1 U11337( .A1(n7840), .A2(n11904), .A3(n10334), .B1(n10173), .B2( n11152), .Y(n11151) );
	a22oi_1 U11338( .A1(n10334), .A2(n11796), .B1(n11846), .B2(n11904), .Y( n11152) );
	inv_1 U11339( .A(n10489), .Y(n7840) );
	nor2_1 U11340( .A(n8238), .B(n11904), .Y(n7921) );
	nand2_1 U11341( .A(n9107), .B(n6335), .Y(n7814) );
	nor3_1 U11342( .A(n7584), .B(n9075), .C(n5890), .Y(n9107) );
	o211ai_1 U11343( .A1(n9740), .A2(n9053), .B1(n8223), .C1(n9741), .Y(n9075) );
	and2_0 U11344( .A(n8225), .B(n9813), .X(n9741) );
	inv_1 U11345( .A(n10334), .Y(n7584) );
	nor3_1 U11346( .A(n8484), .B(n10295), .C(n10164), .Y(n4789) );
	o21ai_0 U11347( .A1(n9323), .A2(n8830), .B1(n6342), .Y(n8484) );
	inv_1 U11348( .A(n9119), .Y(n8830) );
	o21ai_0 U11349( .A1(n6239), .A2(n6052), .B1(n11153), .Y(n4788) );
	mux2i_1 U11350( .A0(n9884), .A1(n11154), .S(n7132), .Y(n11153) );
	inv_1 U11351( .A(n10325), .Y(n7132) );
	nor2_1 U11352( .A(n6291), .B(n6957), .Y(n11154) );
	inv_1 U11353( .A(n6959), .Y(n6957) );
	inv_1 U11354( .A(n6952), .Y(n9884) );
	nand2_1 U11355( .A(n6988), .B(n6379), .Y(n6952) );
	nor2_1 U11356( .A(n6934), .B(n6959), .Y(n6988) );
	nor3_1 U11357( .A(n10266), .B(n10268), .C(n7742), .Y(n6959) );
	o21ai_0 U11358( .A1(n6239), .A2(n6028), .B1(n11155), .Y(n4787) );
	mux2i_1 U11359( .A0(n11156), .A1(n7303), .S(n11157), .Y(n11155) );
	nor2_1 U11360( .A(n10286), .B(n7306), .Y(n11157) );
	inv_1 U11361( .A(n7490), .Y(n7306) );
	nor2_1 U11362( .A(n7596), .B(n7742), .Y(n7490) );
	nor2_1 U11363( .A(n9757), .B(g27831), .Y(n7742) );
	inv_1 U11364( .A(n10268), .Y(n7596) );
	and2_0 U11365( .A(n6345), .B(n11158), .X(n7303) );
	o21ai_0 U11366( .A1(n9593), .A2(n9757), .B1(n9752), .Y(n11158) );
	o211ai_1 U11367( .A1(n10282), .A2(n9830), .B1(n9757), .C1(n9831), .Y(n9752) );
	o211ai_1 U11368( .A1(n10507), .A2(n6910), .B1(n11159), .C1(n11032), .Y( n9757) );
	nand3_1 U11369( .A(n8093), .B(n9378), .C(n10167), .Y(n11159) );
	inv_1 U11370( .A(n10282), .Y(n6910) );
	nor2_1 U11371( .A(n6290), .B(n9095), .Y(n11156) );
	inv_1 U11372( .A(n10738), .Y(n9095) );
	nor2_1 U11373( .A(n6353), .B(n11160), .Y(n4786) );
	o32ai_1 U11374( .A1(n6061), .A2(n6348), .A3(n7464), .B1(n7465), .B2(n9889), .Y(n4785) );
	inv_1 U11375( .A(n10653), .Y(n9889) );
	nand2_1 U11376( .A(n7464), .B(n6380), .Y(n7465) );
	nor2_1 U11377( .A(n6934), .B(n6663), .Y(n7464) );
	o21ai_0 U11378( .A1(n6240), .A2(n10013), .B1(n11161), .Y(n4784) );
	mux2i_1 U11379( .A0(n11162), .A1(n11163), .S(n9626), .Y(n11161) );
	nor2_1 U11380( .A(n6354), .B(n11164), .Y(n11163) );
	and2_0 U11381( .A(n11164), .B(n7237), .X(n11162) );
	inv_1 U11382( .A(n10530), .Y(n10013) );
	o221ai_1 U11383( .A1(n9885), .A2(n8941), .B1(n6214), .B2(n11165), .C1( n11166), .Y(n4783) );
	or3_1 U11384( .A(n6314), .B(n9983), .C(n7072), .X(n11166) );
	nand2_1 U11385( .A(n11960), .B(n11165), .Y(n7072) );
	nand2_1 U11386( .A(n10276), .B(n5904), .Y(n8941) );
	inv_1 U11387( .A(n6483), .Y(n9885) );
	nor2_1 U11388( .A(n9983), .B(n6365), .Y(n6483) );
	nor3_1 U11389( .A(n9323), .B(n10163), .C(n9322), .Y(n9983) );
	nand4_1 U11390( .A(n11839), .B(n10288), .C(n11167), .D(n9390), .Y(n9323) );
	o22ai_1 U11391( .A1(n6211), .A2(n11168), .B1(n11169), .B2(n6298), .Y(n4782) );
	nor2_1 U11392( .A(n11170), .B(n11171), .Y(n11169) );
	mux2i_1 U11393( .A0(n11172), .A1(n11173), .S(n7334), .Y(n11171) );
	nand2_1 U11394( .A(n8453), .B(n11174), .Y(n11173) );
	inv_1 U11395( .A(n6881), .Y(n8453) );
	o21ai_0 U11396( .A1(n11175), .A2(n11176), .B1(n11177), .Y(n6881) );
	inv_1 U11397( .A(g135), .Y(n11177) );
	mux2i_1 U11398( .A0(n11178), .A1(n11179), .S(n9569), .Y(n11176) );
	nand2_1 U11399( .A(n10515), .B(n8714), .Y(n11179) );
	nand3_1 U11400( .A(n8718), .B(n8469), .C(n10269), .Y(n11178) );
	nor3_1 U11401( .A(n11180), .B(n10719), .C(n11181), .Y(n11175) );
	xnor2_1 U11402( .A(n8469), .B(n10341), .Y(n11181) );
	inv_1 U11403( .A(n10515), .Y(n8469) );
	xnor2_1 U11404( .A(n8718), .B(n10269), .Y(n11180) );
	inv_1 U11405( .A(n10353), .Y(n8718) );
	nand2_1 U11406( .A(n10255), .B(n10160), .Y(n11172) );
	a21oi_1 U11407( .A1(n11182), .A2(n7334), .B1(n11174), .Y(n11170) );
	mux2i_1 U11408( .A0(n11183), .A1(n11184), .S(n9566), .Y(n11182) );
	nand2_1 U11409( .A(n11185), .B(n6684), .Y(n11184) );
	mux2_1 U11410( .A0(n10213), .A1(n11186), .S(n7618), .X(n11185) );
	nand2_1 U11411( .A(g90), .B(n5872), .Y(n11186) );
	nor2_1 U11412( .A(n10246), .B(n7612), .Y(n11183) );
	a21oi_1 U11413( .A1(n5960), .A2(n7912), .B1(n6307), .Y(n4781) );
	inv_1 U11414( .A(n10872), .Y(n7912) );
	o21ai_0 U11415( .A1(n11187), .A2(n11188), .B1(n11189), .Y(n4780) );
	o21ai_0 U11416( .A1(n11190), .A2(n11191), .B1(n6342), .Y(n11189) );
	a21oi_1 U11417( .A1(g12919), .A2(n7468), .B1(n10346), .Y(n11190) );
	inv_1 U11418( .A(n10715), .Y(n7468) );
	inv_1 U11419( .A(n10346), .Y(n11188) );
	nor2_1 U11420( .A(n6437), .B(n4753), .Y(n11187) );
	o22ai_1 U11421( .A1(n6810), .A2(n8285), .B1(n7546), .B2(n11192), .Y(n4779) );
	inv_1 U11422( .A(n10870), .Y(n11192) );
	o21ai_0 U11423( .A1(n6819), .A2(n6934), .B1(n6382), .Y(n7546) );
	inv_1 U11424( .A(n10308), .Y(n8285) );
	inv_1 U11425( .A(n8289), .Y(n6810) );
	nor2_1 U11426( .A(n6312), .B(n6819), .Y(n8289) );
	nor2_1 U11427( .A(n6354), .B(n9877), .Y(n4778) );
	inv_1 U11428( .A(g17715), .Y(n9877) );
	o21ai_0 U11429( .A1(n6240), .A2(n8869), .B1(n11193), .Y(n4777) );
	mux2i_1 U11430( .A0(n11194), .A1(n10106), .S(n10105), .Y(n11193) );
	and2_0 U11431( .A(n11195), .B(n6383), .X(n10106) );
	nor2_1 U11432( .A(n11195), .B(n8048), .Y(n11194) );
	inv_1 U11433( .A(n7237), .Y(n8048) );
	a21oi_1 U11434( .A1(n8268), .A2(g11678), .B1(n6308), .Y(n7237) );
	inv_1 U11435( .A(n10664), .Y(n8268) );
	and2_0 U11436( .A(n10385), .B(n8868), .X(n11195) );
	nor2_1 U11437( .A(n7236), .B(n7235), .Y(n8868) );
	inv_1 U11438( .A(n10384), .Y(n7235) );
	nand2_1 U11439( .A(n8047), .B(n10402), .Y(n7236) );
	and2_0 U11440( .A(n10400), .B(n8213), .X(n8047) );
	nor2_1 U11441( .A(n8209), .B(n8514), .Y(n8213) );
	nand2_1 U11442( .A(n10397), .B(n11126), .Y(n8514) );
	and2_0 U11443( .A(n10391), .B(n11036), .X(n11126) );
	nor2_1 U11444( .A(n10077), .B(n10078), .Y(n11036) );
	nand2_1 U11445( .A(n10399), .B(n9630), .Y(n10078) );
	nor2_1 U11446( .A(n11164), .B(n9626), .Y(n9630) );
	inv_1 U11447( .A(n10529), .Y(n9626) );
	nand2_1 U11448( .A(n10530), .B(n10015), .Y(n11164) );
	inv_1 U11449( .A(n10014), .Y(n10015) );
	o211ai_1 U11450( .A1(n10664), .A2(n9826), .B1(n8270), .C1(n11858), .Y( n10014) );
	a21oi_1 U11451( .A1(n9826), .A2(g12184), .B1(n9654), .Y(n8270) );
	o211ai_1 U11452( .A1(n10105), .A2(n10103), .B1(n7941), .C1(n11196), .Y( n9654) );
	mux2i_1 U11453( .A0(n11197), .A1(n11198), .S(n9990), .Y(n11196) );
	nor2_1 U11454( .A(n10426), .B(n10220), .Y(n11198) );
	nor2_1 U11455( .A(n9069), .B(n8886), .Y(n11197) );
	inv_1 U11456( .A(n10220), .Y(n8886) );
	inv_1 U11457( .A(n10426), .Y(n9069) );
	nor3_1 U11458( .A(n10121), .B(n11199), .C(n11200), .Y(n7941) );
	or3_1 U11459( .A(n10199), .B(n10371), .C(n10330), .X(n11200) );
	nand2_1 U11460( .A(n8523), .B(n8525), .Y(n10121) );
	inv_1 U11461( .A(n10926), .Y(n10103) );
	inv_1 U11462( .A(n10551), .Y(n10105) );
	inv_1 U11463( .A(g11678), .Y(n9826) );
	inv_1 U11464( .A(n10393), .Y(n10077) );
	inv_1 U11465( .A(n10385), .Y(n8869) );
	o22ai_1 U11466( .A1(n8166), .A2(n8131), .B1(n11201), .B2(n8169), .Y(n4776) );
	a21oi_1 U11467( .A1(n10964), .A2(n8166), .B1(n6437), .Y(n11201) );
	nor2_1 U11468( .A(n8167), .B(n6365), .Y(n10964) );
	or3_1 U11469( .A(n8167), .B(n10154), .C(n6307), .X(n8131) );
	nor3_1 U11470( .A(n9512), .B(n9322), .C(n9116), .Y(n8167) );
	inv_1 U11471( .A(n10342), .Y(n9322) );
	nand4_1 U11472( .A(n11839), .B(n11167), .C(n9390), .D(n8829), .Y(n9512) );
	inv_1 U11473( .A(n10206), .Y(n8166) );
	o21ai_0 U11474( .A1(n6240), .A2(n8950), .B1(n11202), .Y(n4775) );
	mux2i_1 U11475( .A0(n11203), .A1(n6261), .S(n9985), .Y(n11202) );
	nor2_1 U11476( .A(n8949), .B(n6482), .Y(n9985) );
	nor2_1 U11477( .A(n6310), .B(n7011), .Y(n11203) );
	inv_1 U11478( .A(n10821), .Y(n7011) );
	inv_1 U11479( .A(n10829), .Y(n8950) );
	o221ai_1 U11480( .A1(n7449), .A2(n9241), .B1(n6213), .B2(n7956), .C1(n11204), .Y(n4774) );
	or3_1 U11481( .A(n9093), .B(n6369), .C(n10020), .X(n11204) );
	nor2_1 U11482( .A(n9091), .B(n8885), .Y(n9093) );
	nand2_1 U11483( .A(n10165), .B(n9390), .Y(n8885) );
	inv_1 U11484( .A(n10254), .Y(n7956) );
	nand2_1 U11485( .A(n9243), .B(n6336), .Y(n9241) );
	inv_1 U11486( .A(n9406), .Y(n9243) );
	o21ai_0 U11487( .A1(n6240), .A2(n7230), .B1(n11205), .Y(n4773) );
	mux2i_1 U11488( .A0(n11206), .A1(n6261), .S(n11207), .Y(n11205) );
	nor2_1 U11489( .A(n8069), .B(n6906), .Y(n11207) );
	nand3_1 U11490( .A(n8688), .B(n5902), .C(n7228), .Y(n6906) );
	inv_1 U11491( .A(n10272), .Y(n8688) );
	nor2_1 U11492( .A(n6311), .B(n8334), .Y(n11206) );
	inv_1 U11493( .A(n10767), .Y(n8334) );
	inv_1 U11494( .A(n10766), .Y(n7230) );
	o21ai_0 U11495( .A1(n6240), .A2(n6017), .B1(n11208), .Y(n4772) );
	mux2i_1 U11496( .A0(n11209), .A1(n7021), .S(n11210), .Y(n11208) );
	nor2_1 U11497( .A(n10264), .B(n10020), .Y(n11210) );
	nand2_1 U11498( .A(n10254), .B(n9406), .Y(n10020) );
	nand2_1 U11499( .A(n9407), .B(n9086), .Y(n9406) );
	o21ai_0 U11500( .A1(n11029), .A2(n6407), .B1(g17316), .Y(n9086) );
	inv_1 U11501( .A(n6911), .Y(n6407) );
	nor2_1 U11502( .A(n5884), .B(n10248), .Y(n6911) );
	inv_1 U11503( .A(n11211), .Y(n9407) );
	and2_0 U11504( .A(n6345), .B(n11212), .X(n7021) );
	o21ai_0 U11505( .A1(g23683), .A2(n11211), .B1(n9402), .Y(n11212) );
	o211ai_1 U11506( .A1(n10284), .A2(n9830), .B1(n11211), .C1(n9831), .Y(n9402) );
	o211ai_1 U11507( .A1(n10507), .A2(n8151), .B1(n11213), .C1(n11032), .Y( n11211) );
	nand3_1 U11508( .A(n10167), .B(n8093), .C(n10382), .Y(n11213) );
	inv_1 U11509( .A(n10281), .Y(n8093) );
	inv_1 U11510( .A(n10284), .Y(n8151) );
	nor2_1 U11511( .A(n6309), .B(n5988), .Y(n11209) );
	o22ai_1 U11512( .A1(n6305), .A2(n6749), .B1(n6195), .B2(n11214), .Y(n4771) );
	o32ai_1 U11513( .A1(n7445), .A2(n6348), .A3(n6750), .B1(n6751), .B2(n8846), .Y(n4770) );
	inv_1 U11514( .A(n10311), .Y(n8846) );
	nand2_1 U11515( .A(n6750), .B(n6380), .Y(n6751) );
	nor2_1 U11516( .A(n6934), .B(n7248), .Y(n6750) );
	inv_1 U11517( .A(n10851), .Y(n7445) );
	o21ai_0 U11518( .A1(n6240), .A2(n9501), .B1(n11215), .Y(n4769) );
	mux2i_1 U11519( .A0(n11216), .A1(n6261), .S(n11217), .Y(n11215) );
	nor2_1 U11520( .A(n6870), .B(n7178), .Y(n11217) );
	inv_1 U11521( .A(n8995), .Y(n7178) );
	nor2_1 U11522( .A(n8921), .B(n10204), .Y(n8995) );
	nand2_1 U11523( .A(n10274), .B(n5903), .Y(n6870) );
	nor2_1 U11524( .A(n6308), .B(n7174), .Y(n11216) );
	o21ai_0 U11525( .A1(n6240), .A2(n7966), .B1(n11218), .Y(n4768) );
	mux2i_1 U11526( .A0(n11219), .A1(n6261), .S(n11220), .Y(n11218) );
	nor2_1 U11527( .A(n7016), .B(n8949), .Y(n11220) );
	nand2_1 U11528( .A(n10209), .B(n8745), .Y(n8949) );
	nand3_1 U11529( .A(n11165), .B(n5904), .C(n6482), .Y(n7016) );
	inv_1 U11530( .A(n10276), .Y(n11165) );
	nor2_1 U11531( .A(n6277), .B(n10951), .Y(n11219) );
	inv_1 U11532( .A(n10825), .Y(n10951) );
	inv_1 U11533( .A(n10828), .Y(n7966) );
	o22ai_1 U11534( .A1(n7768), .A2(n5919), .B1(n8890), .B2(n9181), .Y(n4767) );
	o21ai_0 U11535( .A1(n7772), .A2(n6934), .B1(n6382), .Y(n9181) );
	inv_1 U11536( .A(n11199), .Y(n7772) );
	inv_1 U11537( .A(n10881), .Y(n8890) );
	nand2_1 U11538( .A(n6338), .B(n11199), .Y(n7768) );
	nand2_1 U11539( .A(n6524), .B(n7114), .Y(n11199) );
	inv_1 U11540( .A(n10537), .Y(n7114) );
	o21ai_0 U11541( .A1(n6240), .A2(n6018), .B1(n11221), .Y(n4766) );
	mux2i_1 U11542( .A0(n11222), .A1(n6249), .S(n11223), .Y(n11221) );
	nor2_1 U11543( .A(n7186), .B(n8483), .Y(n11223) );
	nand2_1 U11544( .A(n10574), .B(n7253), .Y(n8483) );
	inv_1 U11545( .A(n10295), .Y(n7253) );
	and2_0 U11546( .A(n7257), .B(n6383), .X(n6426) );
	nor2_1 U11547( .A(n6934), .B(n7259), .Y(n7257) );
	nor2_1 U11548( .A(n11224), .B(n10666), .Y(n7259) );
	nor2_1 U11549( .A(n6307), .B(n6019), .Y(n11222) );
	nor2_1 U11550( .A(n6354), .B(n11004), .Y(n4765) );
	inv_1 U11551( .A(g9048), .Y(n11004) );
	o221ai_1 U11552( .A1(n6517), .A2(n8418), .B1(n6213), .B2(n8585), .C1(n8420), .Y(n4764) );
	nand3_1 U11553( .A(n8419), .B(n6376), .C(n10319), .Y(n8420) );
	inv_1 U11554( .A(n10319), .Y(n8585) );
	inv_1 U11555( .A(n10632), .Y(n8418) );
	or2_0 U11556( .A(n6313), .B(n8419), .X(n6517) );
	nor3_1 U11557( .A(n7834), .B(n7833), .C(n5896), .Y(n8419) );
	o211ai_1 U11558( .A1(n9740), .A2(n5886), .B1(n9813), .C1(n11142), .Y(n7833) );
	nand2_1 U11559( .A(n7537), .B(n11225), .Y(n9813) );
	nand3_1 U11560( .A(n10296), .B(n6391), .C(n9315), .Y(n11225) );
	inv_1 U11561( .A(n10332), .Y(n7834) );
	o21ai_0 U11562( .A1(n6240), .A2(n8128), .B1(n11226), .Y(n4763) );
	a22oi_1 U11563( .A1(n8501), .A2(n7064), .B1(n11762), .B2(n7802), .Y(n11226) );
	inv_1 U11564( .A(n8926), .Y(n7802) );
	nand2_1 U11565( .A(n8925), .B(n6380), .Y(n8926) );
	nor2_1 U11566( .A(n6934), .B(n8501), .Y(n8925) );
	and2_0 U11567( .A(n6345), .B(n11227), .X(n7064) );
	o21ai_0 U11568( .A1(n10469), .A2(n8502), .B1(n8495), .Y(n11227) );
	o211ai_1 U11569( .A1(n10258), .A2(n9974), .B1(n8502), .C1(n9975), .Y(n8495) );
	nand2_1 U11570( .A(n10508), .B(n7526), .Y(n9975) );
	inv_1 U11571( .A(n9974), .Y(n7526) );
	nand2_1 U11572( .A(n10670), .B(n9811), .Y(n9974) );
	nor3_1 U11573( .A(n10239), .B(n10260), .C(n7884), .Y(n8501) );
	nor2_1 U11574( .A(n8502), .B(n8088), .Y(n7884) );
	inv_1 U11575( .A(n8085), .Y(n8088) );
	o21ai_0 U11576( .A1(n9810), .A2(n7279), .B1(g17404), .Y(n8085) );
	inv_1 U11577( .A(n8974), .Y(n7279) );
	nor2_1 U11578( .A(n6486), .B(n10923), .Y(n8974) );
	inv_1 U11579( .A(n10237), .Y(n6486) );
	nand4_1 U11580( .A(n10326), .B(n6610), .C(n11861), .D(n11228), .Y(n9810) );
	nor3_1 U11581( .A(n10404), .B(n10470), .C(n10445), .Y(n11228) );
	inv_1 U11582( .A(n10214), .Y(n6610) );
	o211ai_1 U11583( .A1(n10508), .A2(n9431), .B1(n11229), .C1(n9811), .Y(n8502) );
	nand2_1 U11584( .A(n11230), .B(n11231), .Y(n9811) );
	nand3_1 U11585( .A(n10267), .B(n9009), .C(n10060), .Y(n11231) );
	nand3_1 U11586( .A(n10166), .B(n6804), .C(n10432), .Y(n11229) );
	inv_1 U11587( .A(n10728), .Y(n8128) );
	o21ai_0 U11588( .A1(n6240), .A2(n6020), .B1(n11232), .Y(n4762) );
	mux2i_1 U11589( .A0(n11233), .A1(n6430), .S(n11234), .Y(n11232) );
	nor3_1 U11590( .A(n7887), .B(n8593), .C(n7895), .Y(n11234) );
	inv_1 U11591( .A(n8964), .Y(n8593) );
	nand2_1 U11592( .A(n9356), .B(n7886), .Y(n8964) );
	o21ai_0 U11593( .A1(n6409), .A2(n11029), .B1(g17400), .Y(n7886) );
	inv_1 U11594( .A(n11235), .Y(n9356) );
	inv_1 U11595( .A(n10242), .Y(n7887) );
	and2_0 U11596( .A(n6346), .B(n11236), .X(n6430) );
	o21ai_0 U11597( .A1(n11235), .A2(n9593), .B1(n9352), .Y(n11236) );
	o211ai_1 U11598( .A1(n10283), .A2(n9830), .B1(n11235), .C1(n9831), .Y(n9352) );
	or2_0 U11599( .A(n7076), .B(n9830), .X(n9831) );
	nand2_1 U11600( .A(n10670), .B(n11032), .Y(n9830) );
	inv_1 U11601( .A(g23683), .Y(n9593) );
	o211ai_1 U11602( .A1(n10507), .A2(n6966), .B1(n11237), .C1(n11032), .Y( n11235) );
	nand2_1 U11603( .A(n11230), .B(n11238), .Y(n11032) );
	nand3_1 U11604( .A(n8153), .B(n9009), .C(n10267), .Y(n11238) );
	nand3_1 U11605( .A(n10167), .B(n9378), .C(n10281), .Y(n11237) );
	inv_1 U11606( .A(n10382), .Y(n9378) );
	inv_1 U11607( .A(n10283), .Y(n6966) );
	nor2_1 U11608( .A(n6294), .B(n7218), .Y(n11233) );
	inv_1 U11609( .A(n10491), .Y(n7218) );
	o221ai_1 U11610( .A1(n9648), .A2(n11239), .B1(n6213), .B2(n10091), .C1( n11240), .Y(n4761) );
	nand3_1 U11611( .A(n6340), .B(n7535), .C(n10524), .Y(n11240) );
	nand2_1 U11612( .A(n9316), .B(n7537), .Y(n7535) );
	o21ai_0 U11613( .A1(n6917), .A2(n7134), .B1(n7537), .Y(n11239) );
	inv_1 U11614( .A(n10848), .Y(n7134) );
	and2_0 U11615( .A(n9390), .B(g35), .X(n6917) );
	nand3_1 U11616( .A(g35), .B(n11241), .C(n9902), .Y(n9648) );
	nor2_1 U11617( .A(n9424), .B(n6365), .Y(n9902) );
	inv_1 U11618( .A(n9316), .Y(n9424) );
	nor4_1 U11619( .A(n5882), .B(n6397), .C(n6637), .D(n6391), .Y(n9316) );
	inv_1 U11620( .A(n10296), .Y(n6637) );
	nand2_1 U11621( .A(g85), .B(n9390), .Y(n11241) );
	o22ai_1 U11622( .A1(n6303), .A2(n9548), .B1(g23002), .B2(n6197), .Y(n4760) );
	inv_1 U11623( .A(g20652), .Y(n9548) );
	o21ai_0 U11624( .A1(n6240), .A2(n11242), .B1(n11243), .Y(n4759) );
	o221ai_1 U11625( .A1(n11244), .A2(n10603), .B1(g20763), .B2(n10593), .C1( n6382), .Y(n11243) );
	a21oi_1 U11626( .A1(n10593), .A2(n11245), .B1(n6934), .Y(n11244) );
	inv_1 U11627( .A(n10603), .Y(n11242) );
	o22ai_1 U11628( .A1(n6208), .A2(n6080), .B1(n11246), .B2(n6296), .Y(n4758) );
	a221oi_1 U11629( .A1(n11247), .A2(n10463), .B1(n10178), .B2(n6684), .C1( n11248), .Y(n11246) );
	o32ai_1 U11630( .A1(n7934), .A2(n11249), .A3(n11250), .B1(n7938), .B2( n11251), .Y(n11248) );
	inv_1 U11631( .A(n10218), .Y(n7938) );
	inv_1 U11632( .A(n10458), .Y(n7934) );
	o21ai_0 U11633( .A1(n6240), .A2(n5931), .B1(n11252), .Y(n4757) );
	mux2i_1 U11634( .A0(n11253), .A1(n11254), .S(n11255), .Y(n11252) );
	nor2_1 U11635( .A(n7152), .B(n5931), .Y(n11255) );
	nand2_1 U11636( .A(n10543), .B(n11948), .Y(n7152) );
	nor2_1 U11637( .A(g20557), .B(n6365), .Y(n11254) );
	and2_0 U11638( .A(n6346), .B(g20557), .X(n11253) );
	o32ai_1 U11639( .A1(n11256), .A2(g341), .A3(n6313), .B1(n6202), .B2(n11005), .Y(n4756) );
	inv_1 U11640( .A(g20763), .Y(n11005) );
	nand2_1 U11641( .A(n8600), .B(n10879), .Y(n11256) );
	mux2i_1 U11642( .A0(n10185), .A1(n10526), .S(n6975), .Y(n8600) );
	inv_1 U11643( .A(n10485), .Y(n6975) );
	o22ai_1 U11644( .A1(g23612), .A2(n6302), .B1(n6195), .B2(n11257), .Y(n4755) );
	o21ai_0 U11645( .A1(n6240), .A2(n11258), .B1(n11259), .Y(n4754) );
	a22oi_1 U11646( .A1(g21245), .A2(n6701), .B1(n6700), .B2(n6703), .Y(n11259) );
	nand2_1 U11647( .A(n11260), .B(n11261), .Y(n6703) );
	mux2i_1 U11648( .A0(n11262), .A1(n11263), .S(n11264), .Y(n11261) );
	xnor2_1 U11649( .A(n6505), .B(g12238), .Y(n11264) );
	nand3_1 U11650( .A(n11265), .B(n11266), .C(n11267), .Y(n11263) );
	nand3_1 U11651( .A(n10497), .B(g17519), .C(n11268), .Y(n11267) );
	nand3_1 U11652( .A(n11269), .B(g17674), .C(n11793), .Y(n11266) );
	nand3_1 U11653( .A(n11270), .B(g14662), .C(n11803), .Y(n11265) );
	nand3_1 U11654( .A(n11271), .B(n11272), .C(n11273), .Y(n11262) );
	nand3_1 U11655( .A(g17674), .B(n11902), .C(g25114), .Y(n11273) );
	nand3_1 U11656( .A(g17519), .B(n10803), .C(n11270), .Y(n11272) );
	nand3_1 U11657( .A(n11268), .B(g14662), .C(n11903), .Y(n11271) );
	mux2_1 U11658( .A0(n11274), .A1(n11275), .S(n6505), .X(n11260) );
	a221oi_1 U11659( .A1(n11268), .A2(n11276), .B1(g25114), .B2(n11277), .C1( n11278), .Y(n11275) );
	o32ai_1 U11660( .A1(n5939), .A2(n8626), .A3(n11279), .B1(n11280), .B2(n8628), .Y(n11278) );
	a22oi_1 U11661( .A1(n10795), .A2(g17577), .B1(n10796), .B2(g17639), .Y( n11280) );
	inv_1 U11662( .A(n11270), .Y(n8626) );
	o22ai_1 U11663( .A1(n11281), .A2(n7174), .B1(n11282), .B2(n7957), .Y(n11277) );
	inv_1 U11664( .A(n10793), .Y(n7957) );
	inv_1 U11665( .A(n10794), .Y(n7174) );
	o22ai_1 U11666( .A1(n11283), .A2(n8615), .B1(n11284), .B2(n9501), .Y(n11276) );
	inv_1 U11667( .A(n10791), .Y(n9501) );
	inv_1 U11668( .A(n10792), .Y(n8615) );
	inv_1 U11669( .A(n8625), .Y(n11268) );
	a221oi_1 U11670( .A1(n11270), .A2(n11285), .B1(g25114), .B2(n11286), .C1( n11287), .Y(n11274) );
	o32ai_1 U11671( .A1(n5940), .A2(n8625), .A3(n11279), .B1(n11288), .B2(n8628), .Y(n11287) );
	inv_1 U11672( .A(n11269), .Y(n8628) );
	nor2_1 U11673( .A(n8361), .B(n10188), .Y(n11269) );
	a22oi_1 U11674( .A1(n10799), .A2(g12238), .B1(n10800), .B2(g17787), .Y( n11288) );
	nand2_1 U11675( .A(n10188), .B(n8361), .Y(n8625) );
	inv_1 U11676( .A(n10381), .Y(n8361) );
	o22ai_1 U11677( .A1(n9785), .A2(n8875), .B1(n11258), .B2(n11289), .Y(n11286) );
	inv_1 U11678( .A(n10798), .Y(n8875) );
	inv_1 U11679( .A(g17639), .Y(n9785) );
	o22ai_1 U11680( .A1(n11283), .A2(n6785), .B1(n11284), .B2(n8135), .Y(n11285) );
	inv_1 U11681( .A(n10801), .Y(n8135) );
	inv_1 U11682( .A(n10802), .Y(n6785) );
	nor2_1 U11683( .A(n10381), .B(n10188), .Y(n11270) );
	nor2_1 U11684( .A(n8622), .B(n6299), .Y(n6700) );
	nor2_1 U11685( .A(n6284), .B(g28753), .Y(n6701) );
	inv_1 U11686( .A(n10797), .Y(n11258) );
	and2_0 U11687( .A(g12919), .B(n6383), .X(n4753) );
	o22ai_1 U11688( .A1(n11290), .A2(n5954), .B1(n6303), .B2(n11291), .Y(n4752) );
	mux2i_1 U11689( .A0(n10358), .A1(g20899), .S(n10945), .Y(n11291) );
	a21oi_1 U11690( .A1(n8196), .A2(n6381), .B1(n6437), .Y(n11290) );
	inv_1 U11691( .A(n10945), .Y(n8196) );
	nand4_1 U11692( .A(n8960), .B(n7414), .C(n6819), .D(n11292), .Y(n10945) );
	nor2_1 U11693( .A(n9578), .B(n8523), .Y(n11292) );
	inv_1 U11694( .A(n10550), .Y(n8523) );
	nand2_1 U11695( .A(n10199), .B(n10330), .Y(n9578) );
	inv_1 U11696( .A(n9195), .Y(n6819) );
	nand2_1 U11697( .A(n10537), .B(n6524), .Y(n9195) );
	nor3_1 U11698( .A(n7379), .B(n6523), .C(n6526), .Y(n6524) );
	inv_1 U11699( .A(n10921), .Y(n6526) );
	inv_1 U11700( .A(n10294), .Y(n6523) );
	inv_1 U11701( .A(n10669), .Y(n7379) );
	nor2_1 U11702( .A(n6354), .B(n8784), .Y(n4751) );
	inv_1 U11703( .A(g13865), .Y(n8784) );
	nor2_1 U11704( .A(n6354), .B(n7701), .Y(n4750) );
	nor2_1 U11705( .A(n6354), .B(n11096), .Y(n4749) );
	inv_1 U11706( .A(g13881), .Y(n11096) );
	nor2_1 U11707( .A(n6354), .B(n9151), .Y(n4748) );
	inv_1 U11708( .A(g13906), .Y(n9151) );
	nor2_1 U11709( .A(n6354), .B(n8794), .Y(n4747) );
	nor2_1 U11710( .A(n6355), .B(n10051), .Y(n4746) );
	nor2_1 U11711( .A(n6355), .B(n9878), .Y(n4745) );
	nor2_1 U11712( .A(n6355), .B(n9700), .Y(n4744) );
	nor2_1 U11713( .A(n6355), .B(n11293), .Y(n4743) );
	nor2_1 U11714( .A(n6358), .B(n10044), .Y(n4742) );
	inv_1 U11715( .A(g14705), .Y(n10044) );
	nor2_1 U11716( .A(n6355), .B(n11103), .Y(n4741) );
	nor2_1 U11717( .A(n6355), .B(n8789), .Y(n4740) );
	nor2_1 U11718( .A(n6355), .B(n9871), .Y(n4739) );
	nor2_1 U11719( .A(n6355), .B(n7693), .Y(n4738) );
	inv_1 U11720( .A(g14635), .Y(n7693) );
	nor2_1 U11721( .A(n6355), .B(n9695), .Y(n4737) );
	inv_1 U11722( .A(g14749), .Y(n9695) );
	nor2_1 U11723( .A(n6355), .B(n11284), .Y(n4736) );
	nor2_1 U11724( .A(n6355), .B(n11294), .Y(n4735) );
	nor2_1 U11725( .A(n6355), .B(n9157), .Y(n4734) );
	nor2_1 U11726( .A(n6355), .B(n11289), .Y(n4733) );
	nor2_1 U11727( .A(n6356), .B(n11295), .Y(n4732) );
	nor2_1 U11728( .A(n6356), .B(n11279), .Y(n4731) );
	inv_1 U11729( .A(g14597), .Y(n11279) );
	nor2_1 U11730( .A(n6356), .B(n9865), .Y(n4730) );
	inv_1 U11731( .A(g14673), .Y(n9865) );
	nor2_1 U11732( .A(n6356), .B(n9408), .Y(n4729) );
	nor2_1 U11733( .A(n6356), .B(n11109), .Y(n4728) );
	nor2_1 U11734( .A(n6356), .B(n11296), .Y(n4727) );
	nor2_1 U11735( .A(n6356), .B(n11297), .Y(n4726) );
	and2_0 U11736( .A(n6345), .B(g113), .X(n4725) );
	nor2_1 U11737( .A(n6356), .B(n11298), .Y(n4724) );
	nor2_1 U11738( .A(n6356), .B(n11299), .Y(n4723) );
	nor2_1 U11739( .A(n6357), .B(n11300), .Y(n4722) );
	o22ai_1 U11740( .A1(n6209), .A2(n11224), .B1(n6277), .B2(n11301), .Y(n4721) );
	nor2_1 U11741( .A(n6357), .B(n11302), .Y(n4720) );
	nor2_1 U11742( .A(n6357), .B(n11303), .Y(n4719) );
	nor2_1 U11743( .A(n6357), .B(n11304), .Y(n4718) );
	o22ai_1 U11744( .A1(n6209), .A2(n11305), .B1(n6277), .B2(n11306), .Y(n4717) );
	mux2i_1 U11745( .A0(n11302), .A1(n11307), .S(n11224), .Y(n11306) );
	inv_1 U11746( .A(n10670), .Y(n11224) );
	o21ai_0 U11747( .A1(n11308), .A2(n11309), .B1(n11302), .Y(n11307) );
	nand3_1 U11748( .A(n11297), .B(n11298), .C(n11300), .Y(n11309) );
	inv_1 U11749( .A(g11447), .Y(n11300) );
	inv_1 U11750( .A(g8784), .Y(n11298) );
	inv_1 U11751( .A(g8783), .Y(n11297) );
	nand4_1 U11752( .A(n11310), .B(n11311), .C(n11312), .D(n6536), .Y(n11308) );
	inv_1 U11753( .A(g8789), .Y(n6536) );
	inv_1 U11754( .A(g8786), .Y(n11302) );
	inv_1 U11755( .A(n10211), .Y(n11305) );
	nor2_1 U11756( .A(n6357), .B(n11312), .Y(n4716) );
	inv_1 U11757( .A(g8788), .Y(n11312) );
	and2_0 U11758( .A(n6384), .B(g8870), .X(n4715) );
	nor2_1 U11759( .A(n9046), .B(n6299), .Y(n4714) );
	inv_1 U11760( .A(n10510), .Y(n9046) );
	and2_0 U11761( .A(n6384), .B(g14201), .X(n4713) );
	and2_0 U11762( .A(n6384), .B(g8132), .X(n4712) );
	and2_0 U11763( .A(n6384), .B(g8178), .X(n4711) );
	nor2_1 U11764( .A(n6280), .B(n7327), .Y(n4710) );
	inv_1 U11765( .A(n10349), .Y(n7327) );
	nor2_1 U11766( .A(n8745), .B(n6299), .Y(n4709) );
	inv_1 U11767( .A(n10513), .Y(n8745) );
	and2_0 U11768( .A(n6386), .B(g14147), .X(n4708) );
	o22ai_1 U11769( .A1(n11799), .A2(n6302), .B1(n6195), .B2(n11245), .Y(n4707) );
	inv_1 U11770( .A(n10210), .Y(n11245) );
	nor2_1 U11771( .A(n6281), .B(n9618), .Y(n4706) );
	inv_1 U11772( .A(n10350), .Y(n9618) );
	inv_1 U11773( .A(n11313), .Y(n4705) );
	nor2_1 U11774( .A(n6283), .B(n11314), .Y(n4704) );
	and2_0 U11775( .A(n6384), .B(g14189), .X(n4703) );
	and2_0 U11776( .A(g125), .B(n6344), .X(n4702) );
	and2_0 U11777( .A(n6383), .B(g14096), .X(n4701) );
	and2_0 U11778( .A(n6384), .B(g14125), .X(n4700) );
	inv_1 U11779( .A(n11315), .Y(n47) );
	nor2_1 U11780( .A(n6282), .B(n6566), .Y(n4699) );
	inv_1 U11781( .A(n10352), .Y(n6566) );
	and2_0 U11782( .A(n6384), .B(g14217), .X(n4698) );
	nor2_1 U11783( .A(n9600), .B(n6300), .Y(n4697) );
	inv_1 U11784( .A(n10512), .Y(n9600) );
	nor2_1 U11785( .A(n9805), .B(n6299), .Y(n4696) );
	inv_1 U11786( .A(n10511), .Y(n9805) );
	and2_0 U11787( .A(n6385), .B(g8235), .X(n4695) );
	and2_0 U11788( .A(n6385), .B(g8283), .X(n4694) );
	o221ai_1 U11789( .A1(n6212), .A2(n5958), .B1(n6301), .B2(n6979), .C1(n6978), .Y(n4693) );
	inv_1 U11790( .A(n8598), .Y(n6978) );
	nor2_1 U11791( .A(n11127), .B(n6300), .Y(n8598) );
	inv_1 U11792( .A(n10185), .Y(n11127) );
	inv_1 U11793( .A(n10526), .Y(n6979) );
	mux2i_1 U11794( .A0(n11316), .A1(n11317), .S(n10914), .Y(n4692) );
	a21oi_1 U11795( .A1(n11318), .A2(n6382), .B1(n6437), .Y(n11317) );
	or2_0 U11796( .A(n11318), .B(n6286), .X(n11316) );
	o21ai_0 U11797( .A1(n6240), .A2(n6880), .B1(n11319), .Y(n4691) );
	nand4_1 U11798( .A(n8714), .B(n9569), .C(n11320), .D(n11321), .Y(n11319) );
	nor4_1 U11799( .A(n11322), .B(n7334), .C(n6879), .D(n11323), .Y(n11321) );
	inv_1 U11800( .A(n10407), .Y(n6879) );
	inv_1 U11801( .A(n6882), .Y(n11322) );
	nor3_1 U11802( .A(n10353), .B(n10719), .C(n10515), .Y(n11320) );
	inv_1 U11803( .A(n10341), .Y(n9569) );
	inv_1 U11804( .A(n10269), .Y(n8714) );
	nor2_1 U11805( .A(n6357), .B(n11324), .Y(n4690) );
	mux2i_1 U11806( .A0(n11325), .A1(n11326), .S(n10915), .Y(n4689) );
	a21oi_1 U11807( .A1(n11327), .A2(n6378), .B1(n6437), .Y(n11326) );
	or2_0 U11808( .A(n11327), .B(n6311), .X(n11325) );
	nor2_1 U11809( .A(n6357), .B(n11310), .Y(n4688) );
	inv_1 U11810( .A(g8785), .Y(n11310) );
	nor3_1 U11811( .A(n11328), .B(n6278), .C(n11329), .Y(n4687) );
	mux2i_1 U11812( .A0(n11330), .A1(g11388), .S(g13926), .Y(n11329) );
	nand3_1 U11813( .A(n11331), .B(n11109), .C(n11103), .Y(n11328) );
	inv_1 U11814( .A(g14451), .Y(n11103) );
	inv_1 U11815( .A(g16656), .Y(n11109) );
	nor3_1 U11816( .A(n11332), .B(n6278), .C(n11333), .Y(n4686) );
	mux2i_1 U11817( .A0(n11334), .A1(g12470), .S(g14828), .Y(n11333) );
	nand3_1 U11818( .A(n11335), .B(n9408), .C(n9700), .Y(n11332) );
	inv_1 U11819( .A(g13099), .Y(n9700) );
	inv_1 U11820( .A(g17722), .Y(n9408) );
	nor3_1 U11821( .A(n11336), .B(n6278), .C(n11337), .Y(n4685) );
	mux2i_1 U11822( .A0(n11338), .A1(g11418), .S(g13966), .Y(n11337) );
	nand3_1 U11823( .A(n11339), .B(n9157), .C(n11295), .Y(n11336) );
	inv_1 U11824( .A(g14518), .Y(n11295) );
	inv_1 U11825( .A(g16693), .Y(n9157) );
	nor3_1 U11826( .A(n11340), .B(n6278), .C(n11341), .Y(n4684) );
	mux2i_1 U11827( .A0(n11342), .A1(g11349), .S(g13895), .Y(n11341) );
	nand3_1 U11828( .A(n11343), .B(n8794), .C(n8789), .Y(n11340) );
	inv_1 U11829( .A(g14421), .Y(n8789) );
	inv_1 U11830( .A(g16624), .Y(n8794) );
	nor2_1 U11831( .A(n6289), .B(n8921), .Y(n4683) );
	inv_1 U11832( .A(n10351), .Y(n8921) );
	nor3_1 U11833( .A(n11344), .B(n6278), .C(n11345), .Y(n4682) );
	mux2i_1 U11834( .A0(n11346), .A1(g12422), .S(g14779), .Y(n11345) );
	nand3_1 U11835( .A(n11347), .B(n10051), .C(n11293), .Y(n11344) );
	inv_1 U11836( .A(g13085), .Y(n11293) );
	inv_1 U11837( .A(g17685), .Y(n10051) );
	o221ai_1 U11838( .A1(n6368), .A2(n11348), .B1(n6508), .B2(n11313), .C1( n6225), .Y(n4681) );
	nand2_1 U11839( .A(g4467), .B(n6379), .Y(n11313) );
	inv_1 U11840( .A(n10364), .Y(n6508) );
	nor2_1 U11841( .A(n7871), .B(n10297), .Y(n11348) );
	inv_1 U11842( .A(n7999), .Y(n7871) );
	nand3_1 U11843( .A(n11349), .B(n5957), .C(g26960), .Y(n7999) );
	o21ai_0 U11844( .A1(n11779), .A2(n9969), .B1(n6684), .Y(n11349) );
	o22ai_1 U11845( .A1(n6303), .A2(n6505), .B1(n6195), .B2(n9510), .Y(n4680) );
	inv_1 U11846( .A(n10151), .Y(n9510) );
	nor3_1 U11847( .A(n6307), .B(n10669), .C(g8719), .Y(n4679) );
	nor3_1 U11848( .A(n11350), .B(n6278), .C(n11351), .Y(n4678) );
	mux2i_1 U11849( .A0(n11352), .A1(g12238), .S(g14662), .Y(n11351) );
	nand3_1 U11850( .A(n11353), .B(n11289), .C(n11284), .Y(n11350) );
	inv_1 U11851( .A(g13039), .Y(n11284) );
	inv_1 U11852( .A(g17577), .Y(n11289) );
	nor3_1 U11853( .A(n11354), .B(n6278), .C(n11355), .Y(n4677) );
	mux2i_1 U11854( .A0(n11356), .A1(g12300), .S(g14694), .Y(n11355) );
	nand3_1 U11855( .A(n11357), .B(n7701), .C(n11294), .Y(n11354) );
	inv_1 U11856( .A(g13049), .Y(n11294) );
	inv_1 U11857( .A(g17604), .Y(n7701) );
	nor3_1 U11858( .A(n11358), .B(n6278), .C(n11359), .Y(n4676) );
	mux2i_1 U11859( .A0(n11360), .A1(g12350), .S(g14738), .Y(n11359) );
	nand3_1 U11860( .A(n11361), .B(n9878), .C(n9871), .Y(n11358) );
	inv_1 U11861( .A(g13068), .Y(n9871) );
	inv_1 U11862( .A(g17646), .Y(n9878) );
	nor4_1 U11863( .A(n11362), .B(g17291), .C(g17400), .D(g17316), .Y(n4675) );
	o21ai_0 U11864( .A1(n9553), .A2(n11363), .B1(n6342), .Y(n11362) );
	o21ai_0 U11865( .A1(n9947), .A2(n7425), .B1(n10405), .Y(n11363) );
	inv_1 U11866( .A(n7972), .Y(n7425) );
	inv_1 U11867( .A(n11364), .Y(n9947) );
	inv_1 U11868( .A(n7554), .Y(n9553) );
	nor2_1 U11869( .A(n7736), .B(n7737), .Y(n7554) );
	nand2_1 U11870( .A(n10215), .B(n10718), .Y(n7737) );
	inv_1 U11871( .A(n10471), .Y(n7736) );
	and2_0 U11872( .A(n6385), .B(g17320), .X(n4674) );
	and2_0 U11873( .A(n6385), .B(g17291), .X(n4673) );
	nor4_1 U11874( .A(n11365), .B(g17320), .C(g17423), .D(g17404), .Y(n4672) );
	o21ai_0 U11875( .A1(n7260), .A2(n11366), .B1(n6343), .Y(n11365) );
	o21ai_0 U11876( .A1(n8973), .A2(n6715), .B1(n6828), .Y(n11366) );
	nor2_1 U11877( .A(n6823), .B(n9524), .Y(n6828) );
	nand2_1 U11878( .A(n10214), .B(n10717), .Y(n9524) );
	inv_1 U11879( .A(n10470), .Y(n6823) );
	inv_1 U11880( .A(n6714), .Y(n6715) );
	inv_1 U11881( .A(n11367), .Y(n8973) );
	and2_0 U11882( .A(n6385), .B(g12184), .X(n4671) );
	and2_0 U11883( .A(n6386), .B(g12368), .X(n4670) );
	nor2_1 U11884( .A(n6357), .B(n7696), .Y(n4669) );
	inv_1 U11885( .A(g17813), .Y(n7696) );
	nor2_1 U11886( .A(n6357), .B(n9868), .Y(n4668) );
	inv_1 U11887( .A(g17819), .Y(n9868) );
	nor2_1 U11888( .A(n6357), .B(n10048), .Y(n4667) );
	inv_1 U11889( .A(g17845), .Y(n10048) );
	nor2_1 U11890( .A(n6358), .B(n9697), .Y(n4666) );
	inv_1 U11891( .A(g17871), .Y(n9697) );
	nor2_1 U11892( .A(n6358), .B(n9155), .Y(n4665) );
	inv_1 U11893( .A(g16955), .Y(n9155) );
	nor2_1 U11894( .A(n6358), .B(n11281), .Y(n4664) );
	inv_1 U11895( .A(g17787), .Y(n11281) );
	nor2_1 U11896( .A(n6358), .B(n11100), .Y(n4663) );
	inv_1 U11897( .A(g16924), .Y(n11100) );
	nor2_1 U11898( .A(n6358), .B(n8786), .Y(n4662) );
	inv_1 U11899( .A(g16874), .Y(n8786) );
	o22ai_1 U11900( .A1(n6211), .A2(n11368), .B1(n11369), .B2(n6296), .Y(n4661) );
	xnor2_1 U11901( .A(g8358), .B(n11370), .Y(n11369) );
	nor2_1 U11902( .A(n8031), .B(n8032), .Y(n11370) );
	nand2_1 U11903( .A(n10936), .B(g8291), .Y(n8032) );
	xnor2_1 U11904( .A(g8358), .B(n5920), .Y(n8031) );
	inv_1 U11905( .A(n10663), .Y(n11368) );
	nor2_1 U11906( .A(n6287), .B(n11371), .Y(n4660) );
	xnor2_1 U11907( .A(n9220), .B(n9584), .Y(n11371) );
	xor2_1 U11908( .A(g9251), .B(n11892), .X(n9584) );
	inv_1 U11909( .A(g9251), .Y(n9220) );
	and2_0 U11910( .A(n6371), .B(g17316), .X(n4659) );
	and2_0 U11911( .A(n6386), .B(g17404), .X(n4658) );
	o22ai_1 U11912( .A1(n6211), .A2(n11372), .B1(n6277), .B2(n11373), .Y(n4657) );
	xnor2_1 U11913( .A(n7773), .B(n8326), .Y(n11373) );
	xor2_1 U11914( .A(g9019), .B(n11964), .X(n8326) );
	inv_1 U11915( .A(g9019), .Y(n7773) );
	inv_1 U11916( .A(n10666), .Y(n11372) );
	o22ai_1 U11917( .A1(n6211), .A2(n7777), .B1(n6277), .B2(n11374), .Y(n4656) );
	xnor2_1 U11918( .A(g8839), .B(n6544), .Y(n11374) );
	xnor2_1 U11919( .A(g8839), .B(n11897), .Y(n6544) );
	nor2_1 U11920( .A(n6358), .B(n11343), .Y(n4655) );
	inv_1 U11921( .A(g16603), .Y(n11343) );
	nor2_1 U11922( .A(n6358), .B(n11342), .Y(n4654) );
	inv_1 U11923( .A(g16718), .Y(n11342) );
	nor2_1 U11924( .A(n6358), .B(n11334), .Y(n4653) );
	inv_1 U11925( .A(g17778), .Y(n11334) );
	nor2_1 U11926( .A(n6351), .B(n11335), .Y(n4652) );
	inv_1 U11927( .A(g17688), .Y(n11335) );
	nor2_1 U11928( .A(n6358), .B(n11352), .Y(n4651) );
	inv_1 U11929( .A(g17674), .Y(n11352) );
	nor2_1 U11930( .A(n6357), .B(n11339), .Y(n4650) );
	inv_1 U11931( .A(g16659), .Y(n11339) );
	nor2_1 U11932( .A(n6357), .B(n11361), .Y(n4649) );
	inv_1 U11933( .A(g17607), .Y(n11361) );
	nor2_1 U11934( .A(n6357), .B(n11353), .Y(n4648) );
	inv_1 U11935( .A(g17519), .Y(n11353) );
	nor2_1 U11936( .A(n6356), .B(n11346), .Y(n4647) );
	inv_1 U11937( .A(g17760), .Y(n11346) );
	nor2_1 U11938( .A(n6356), .B(n11356), .Y(n4646) );
	inv_1 U11939( .A(g17711), .Y(n11356) );
	nor2_1 U11940( .A(n6356), .B(n11330), .Y(n4645) );
	inv_1 U11941( .A(g16744), .Y(n11330) );
	nor2_1 U11942( .A(n6356), .B(n11338), .Y(n4644) );
	inv_1 U11943( .A(g16775), .Y(n11338) );
	nor2_1 U11944( .A(n6354), .B(n11347), .Y(n4643) );
	inv_1 U11945( .A(g17649), .Y(n11347) );
	nor2_1 U11946( .A(n6354), .B(n11360), .Y(n4642) );
	inv_1 U11947( .A(g17739), .Y(n11360) );
	nor2_1 U11948( .A(n6354), .B(n11357), .Y(n4641) );
	inv_1 U11949( .A(g17580), .Y(n11357) );
	nor2_1 U11950( .A(n6354), .B(n11331), .Y(n4640) );
	inv_1 U11951( .A(g16627), .Y(n11331) );
	o21ai_0 U11952( .A1(n6240), .A2(n7260), .B1(n11375), .Y(n4639) );
	nand2_1 U11953( .A(g496), .B(n6336), .Y(n11375) );
	inv_1 U11954( .A(n10404), .Y(n7260) );
	and2_0 U11955( .A(n6386), .B(g19357), .X(n4638) );
	o22ai_1 U11956( .A1(n6303), .A2(n11376), .B1(n6195), .B2(n7553), .Y(n4637) );
	inv_1 U11957( .A(n10405), .Y(n7553) );
	and2_0 U11958( .A(n6386), .B(g14828), .X(n4636) );
	and2_0 U11959( .A(n6386), .B(g13895), .X(n4635) );
	and2_0 U11960( .A(n6386), .B(g13926), .X(n4634) );
	and2_0 U11961( .A(n6387), .B(g14662), .X(n4633) );
	and2_0 U11962( .A(n6387), .B(g14738), .X(n4632) );
	and2_0 U11963( .A(n6387), .B(g14779), .X(n4631) );
	and2_0 U11964( .A(n6387), .B(g13966), .X(n4630) );
	and2_0 U11965( .A(n6387), .B(g14694), .X(n4629) );
	nor2_1 U11966( .A(n6353), .B(n11191), .Y(n4628) );
	inv_1 U11967( .A(g19334), .Y(n11191) );
	nor2_1 U11968( .A(n6353), .B(n7697), .Y(n4627) );
	inv_1 U11969( .A(g12300), .Y(n7697) );
	nor2_1 U11970( .A(n6353), .B(n9698), .Y(n4626) );
	inv_1 U11971( .A(g12470), .Y(n9698) );
	nor2_1 U11972( .A(n6353), .B(n11282), .Y(n4625) );
	inv_1 U11973( .A(g12238), .Y(n11282) );
	nor2_1 U11974( .A(n6352), .B(n8787), .Y(n4624) );
	inv_1 U11975( .A(g11349), .Y(n8787) );
	nor2_1 U11976( .A(n6352), .B(n11101), .Y(n4623) );
	inv_1 U11977( .A(g11388), .Y(n11101) );
	nor2_1 U11978( .A(n6352), .B(n9156), .Y(n4622) );
	inv_1 U11979( .A(g11418), .Y(n9156) );
	nor2_1 U11980( .A(n6352), .B(n9869), .Y(n4621) );
	inv_1 U11981( .A(g12350), .Y(n9869) );
	nor2_1 U11982( .A(n6351), .B(n10049), .Y(n4620) );
	inv_1 U11983( .A(g12422), .Y(n10049) );
	o22ai_1 U11984( .A1(n6212), .A2(n10126), .B1(n11377), .B2(n6295), .Y(n4619) );
	xor2_1 U11985( .A(n11327), .B(n11378), .X(n11377) );
	nor3_1 U11986( .A(n9815), .B(g8416), .C(g13259), .Y(n11378) );
	nand2_1 U11987( .A(n9818), .B(n7098), .Y(n9815) );
	nor2_1 U11988( .A(n10915), .B(g19334), .Y(n9818) );
	nand3_1 U11989( .A(n11364), .B(n11379), .C(n7972), .Y(n11327) );
	nor2_1 U11990( .A(n9780), .B(n8519), .Y(n7972) );
	nor2_1 U11991( .A(n10915), .B(n10179), .Y(n8519) );
	inv_1 U11992( .A(n11051), .Y(n9780) );
	xor2_1 U11993( .A(n10457), .B(n10179), .X(n11051) );
	xnor2_1 U11994( .A(n5944), .B(n10179), .Y(n11379) );
	inv_1 U11995( .A(n10457), .Y(n10126) );
	and2_0 U11996( .A(n6387), .B(g33079), .X(n4618) );
	and2_0 U11997( .A(n6387), .B(g33435), .X(n4617) );
	o22ai_1 U11998( .A1(n6212), .A2(g23759), .B1(n6347), .B2(n8304), .Y(n4616) );
	o221ai_1 U11999( .A1(n8224), .A2(n11380), .B1(n9425), .B2(n11381), .C1( n11382), .Y(n8304) );
	a21oi_1 U12000( .A1(n11383), .A2(n8225), .B1(n6934), .Y(n11382) );
	inv_1 U12001( .A(n11384), .Y(n11383) );
	mux4_2 U12002( .A0(n10547), .A1(n10548), .A2(n10091), .A3(n8303), .S0(n8223), .S1(n11385), .X(n11384) );
	inv_1 U12003( .A(n10524), .Y(n8303) );
	inv_1 U12004( .A(n10525), .Y(n10091) );
	mux2_1 U12005( .A0(n10554), .A1(n9645), .S(n11385), .X(n11381) );
	mux2_1 U12006( .A0(n10345), .A1(n5885), .S(n11385), .X(n11380) );
	o211ai_1 U12007( .A1(n6203), .A2(n5959), .B1(n6761), .C1(n11386), .Y(n4615) );
	nor2_1 U12008( .A(n6352), .B(n11387), .Y(n4614) );
	nand3_1 U12009( .A(n6760), .B(n6686), .C(n11388), .Y(n4613) );
	nand2_1 U12010( .A(g4567), .B(n6763), .Y(n11388) );
	nand3_1 U12011( .A(n6760), .B(n6889), .C(n11389), .Y(n4612) );
	nand2_1 U12012( .A(g4498), .B(n6763), .Y(n11389) );
	nand2_1 U12013( .A(n11390), .B(n11251), .Y(n6760) );
	inv_1 U12014( .A(n11391), .Y(n11251) );
	o211ai_1 U12015( .A1(n6203), .A2(n5957), .B1(n9513), .C1(n11386), .Y(n4611) );
	inv_1 U12016( .A(n11392), .Y(n11386) );
	o32ai_1 U12017( .A1(n19467), .A2(n10380), .A3(n6313), .B1(n11393), .B2( n6685), .Y(n11392) );
	nor2_1 U12018( .A(n11249), .B(n11250), .Y(n11393) );
	o32ai_1 U12019( .A1(n11323), .A2(n10245), .A3(n5949), .B1(n6202), .B2( n11394), .Y(n4610) );
	nand4_1 U12020( .A(n9566), .B(n7612), .C(n7618), .D(n11395), .Y(n11323) );
	nor2_1 U12021( .A(n6278), .B(n11174), .Y(n11395) );
	nand2_1 U12022( .A(n6880), .B(n7338), .Y(n11174) );
	inv_1 U12023( .A(n10246), .Y(n7618) );
	inv_1 U12024( .A(n10279), .Y(n9566) );
	and2_0 U12025( .A(g26959), .B(n6383), .X(n4609) );
	o22ai_1 U12026( .A1(n6303), .A2(n10133), .B1(n6196), .B2(n6086), .Y(n4608) );
	inv_1 U12027( .A(g6750), .Y(n10133) );
	nor2_1 U12028( .A(n6352), .B(n11396), .Y(n4607) );
	inv_1 U12029( .A(n11397), .Y(n4606) );
	a21oi_1 U12030( .A1(n6437), .A2(n11908), .B1(n39), .Y(n11397) );
	nand3_1 U12031( .A(n11398), .B(n9513), .C(n11399), .Y(n4605) );
	nand2_1 U12032( .A(g4495), .B(n6763), .Y(n11399) );
	nand2_1 U12033( .A(g20049), .B(n11390), .Y(n9513) );
	nand3_1 U12034( .A(n11398), .B(n6889), .C(n11400), .Y(n4604) );
	nand2_1 U12035( .A(g4480), .B(n6763), .Y(n11400) );
	nand2_1 U12036( .A(n11908), .B(n11390), .Y(n6889) );
	nand3_1 U12037( .A(n11398), .B(n6686), .C(n11401), .Y(n4603) );
	nand2_1 U12038( .A(g4540), .B(n6763), .Y(n11401) );
	nand2_1 U12039( .A(g4578), .B(n11390), .Y(n6686) );
	o22ai_1 U12040( .A1(n6211), .A2(n11376), .B1(n11402), .B2(n6295), .Y(n4602) );
	a222oi_1 U12041( .A1(n10187), .A2(n6684), .B1(n11391), .B2(n10302), .C1( n11247), .C2(n10459), .Y(n11402) );
	nor2_1 U12042( .A(n11250), .B(g73), .Y(n11391) );
	inv_1 U12043( .A(g72), .Y(n11250) );
	inv_1 U12044( .A(g20901), .Y(n11376) );
	nand3_1 U12045( .A(n11398), .B(n6761), .C(n11403), .Y(n4601) );
	nand2_1 U12046( .A(g4543), .B(n6763), .Y(n11403) );
	a21oi_1 U12047( .A1(g35), .A2(n10380), .B1(n6368), .Y(n6763) );
	nand2_1 U12048( .A(n11965), .B(n11390), .Y(n6761) );
	or2_0 U12049( .A(n6685), .B(n11247), .X(n11398) );
	nor2_1 U12050( .A(n11249), .B(g72), .Y(n11247) );
	inv_1 U12051( .A(g73), .Y(n11249) );
	nor2_1 U12052( .A(n6352), .B(n11394), .Y(n4600) );
	o22ai_1 U12053( .A1(n6212), .A2(n9962), .B1(n6277), .B2(n11404), .Y(n46) );
	mux2i_1 U12054( .A0(n10186), .A1(n10457), .S(n11405), .Y(n11404) );
	nor2_1 U12055( .A(n7098), .B(n6409), .Y(n11405) );
	inv_1 U12056( .A(n7766), .Y(n6409) );
	nor2_1 U12057( .A(n5884), .B(n6406), .Y(n7766) );
	inv_1 U12058( .A(g7916), .Y(n7098) );
	inv_1 U12059( .A(n10472), .Y(n9962) );
	nor2_1 U12060( .A(n6352), .B(n9450), .Y(n4599) );
	o22ai_1 U12061( .A1(n8975), .A2(n6202), .B1(n11406), .B2(n6295), .Y(n4598) );
	xor2_1 U12062( .A(n11318), .B(n11407), .X(n11406) );
	nor3_1 U12063( .A(n7898), .B(g8475), .C(g13272), .Y(n11407) );
	or3_1 U12064( .A(g7946), .B(n10914), .C(g19357), .X(n7898) );
	nand3_1 U12065( .A(n11367), .B(n11408), .C(n6714), .Y(n11318) );
	nor2_1 U12066( .A(n7787), .B(n7402), .Y(n6714) );
	nor2_1 U12067( .A(n10914), .B(n10326), .Y(n7402) );
	inv_1 U12068( .A(n9661), .Y(n7787) );
	xor2_1 U12069( .A(n10456), .B(n10326), .X(n9661) );
	xnor2_1 U12070( .A(n5945), .B(n10326), .Y(n11408) );
	inv_1 U12071( .A(n10456), .Y(n8975) );
	o22ai_1 U12072( .A1(n6304), .A2(n5958), .B1(n6196), .B2(n11314), .Y(n4597) );
	inv_1 U12073( .A(g21176), .Y(n11314) );
	o22ai_1 U12074( .A1(n6302), .A2(n7167), .B1(n6196), .B2(n11409), .Y(n4596) );
	inv_1 U12075( .A(n10618), .Y(n11409) );
	o22ai_1 U12076( .A1(n6300), .A2(n8769), .B1(n6196), .B2(n11410), .Y(n4595) );
	inv_1 U12077( .A(n10620), .Y(n11410) );
	o22ai_1 U12078( .A1(n6212), .A2(n11411), .B1(n6277), .B2(n11412), .Y(n4594) );
	mux2i_1 U12079( .A0(n11413), .A1(n11414), .S(g8870), .Y(n11412) );
	xnor2_1 U12080( .A(n11411), .B(n11301), .Y(n11414) );
	xnor2_1 U12081( .A(n11415), .B(n11301), .Y(n11413) );
	mux2_1 U12082( .A0(n11945), .A1(n11876), .S(n10466), .X(n11301) );
	o21ai_0 U12083( .A1(n11416), .A2(n11417), .B1(n11411), .Y(n11415) );
	nand3_1 U12084( .A(n11299), .B(n11296), .C(n11304), .Y(n11417) );
	inv_1 U12085( .A(g11770), .Y(n11304) );
	inv_1 U12086( .A(g8916), .Y(n11296) );
	inv_1 U12087( .A(g8915), .Y(n11299) );
	nand4_1 U12088( .A(n11324), .B(n11418), .C(n11303), .D(n11160), .Y(n11416) );
	inv_1 U12089( .A(g8920), .Y(n11160) );
	inv_1 U12090( .A(g8919), .Y(n11303) );
	inv_1 U12091( .A(g8917), .Y(n11324) );
	inv_1 U12092( .A(n10891), .Y(n11411) );
	a21oi_1 U12093( .A1(n6198), .A2(n11419), .B1(n8298), .Y(n4593) );
	inv_1 U12094( .A(n10905), .Y(n8298) );
	nand2_1 U12095( .A(n8297), .B(n6822), .Y(n11419) );
	and2_0 U12096( .A(n8299), .B(n6383), .X(n8297) );
	and2_0 U12097( .A(n10098), .B(n10410), .X(n8299) );
	nor2_1 U12098( .A(n8323), .B(n8324), .Y(n10098) );
	nand2_1 U12099( .A(n10566), .B(n9789), .Y(n8324) );
	and2_0 U12100( .A(n10568), .B(n9723), .X(n9789) );
	nor2_1 U12101( .A(n7082), .B(n7081), .Y(n9723) );
	inv_1 U12102( .A(n10570), .Y(n7081) );
	nand4_1 U12103( .A(n10450), .B(n10389), .C(n10572), .D(g12919), .Y(n7082) );
	inv_1 U12104( .A(n10542), .Y(n8323) );
	a21oi_1 U12105( .A1(n6198), .A2(n11420), .B1(n7542), .Y(n4592) );
	inv_1 U12106( .A(n10904), .Y(n7542) );
	nand2_1 U12107( .A(n7541), .B(n8113), .Y(n11420) );
	and2_0 U12108( .A(n7543), .B(n6383), .X(n7541) );
	and2_0 U12109( .A(n8179), .B(n10409), .X(n7543) );
	nor2_1 U12110( .A(n8175), .B(n9360), .Y(n8179) );
	nand2_1 U12111( .A(n10565), .B(n8041), .Y(n9360) );
	and2_0 U12112( .A(n10567), .B(n9417), .X(n8041) );
	nor2_1 U12113( .A(n8200), .B(n8201), .Y(n9417) );
	nand4_1 U12114( .A(n10571), .B(n10388), .C(n10621), .D(g12923), .Y(n8201) );
	inv_1 U12115( .A(n10569), .Y(n8200) );
	inv_1 U12116( .A(n10541), .Y(n8175) );
	o22ai_1 U12117( .A1(n6298), .A2(n7377), .B1(n6196), .B2(n11421), .Y(n4591) );
	inv_1 U12118( .A(n10612), .Y(n11421) );
	o22ai_1 U12119( .A1(n6295), .A2(n9135), .B1(n6196), .B2(n11422), .Y(n4590) );
	inv_1 U12120( .A(n10616), .Y(n11422) );
	o22ai_1 U12121( .A1(n6297), .A2(n9165), .B1(n6196), .B2(n11423), .Y(n4589) );
	inv_1 U12122( .A(n10609), .Y(n11423) );
	o22ai_1 U12123( .A1(n6302), .A2(n7474), .B1(n6197), .B2(n11424), .Y(n4588) );
	inv_1 U12124( .A(n10605), .Y(n11424) );
	o22ai_1 U12125( .A1(n6302), .A2(n9842), .B1(n6197), .B2(n11425), .Y(n4587) );
	inv_1 U12126( .A(n10607), .Y(n11425) );
	o22ai_1 U12127( .A1(n6212), .A2(n5870), .B1(n11426), .B2(n11427), .Y(n4586) );
	inv_1 U12128( .A(n11428), .Y(n11427) );
	o21ai_0 U12129( .A1(n11429), .A2(n6314), .B1(n11430), .Y(n11428) );
	nor3_1 U12130( .A(n11429), .B(n10443), .C(n8452), .Y(n11426) );
	nor4_1 U12131( .A(n5967), .B(n5880), .C(n5865), .D(n5870), .Y(n8452) );
	o221ai_1 U12132( .A1(n10024), .A2(n11431), .B1(n6219), .B2(n9534), .C1( n11432), .Y(n4585) );
	nand3_1 U12133( .A(g12923), .B(g35), .C(n75), .Y(n11432) );
	nor2_1 U12134( .A(n11433), .B(n6364), .Y(n75) );
	inv_1 U12135( .A(n10688), .Y(n9534) );
	nand2_1 U12136( .A(n6337), .B(n11433), .Y(n11431) );
	inv_1 U12137( .A(g17423), .Y(n11433) );
	inv_1 U12138( .A(g10527), .Y(n10024) );
	o21ai_0 U12139( .A1(n6240), .A2(n9990), .B1(n11315), .Y(n4584) );
	nand2_1 U12140( .A(g64), .B(n6336), .Y(n11315) );
	inv_1 U12141( .A(n10713), .Y(n9990) );
	o221ai_1 U12142( .A1(n8508), .A2(n11434), .B1(n6219), .B2(n6586), .C1( n11435), .Y(n4583) );
	nand3_1 U12143( .A(g12919), .B(g35), .C(n95), .Y(n11435) );
	nor2_1 U12144( .A(n11436), .B(n6363), .Y(n95) );
	inv_1 U12145( .A(n10689), .Y(n6586) );
	nand2_1 U12146( .A(n6339), .B(n11436), .Y(n11434) );
	inv_1 U12147( .A(g17400), .Y(n11436) );
	inv_1 U12148( .A(g10500), .Y(n8508) );
	o22ai_1 U12149( .A1(n10936), .A2(n6302), .B1(n6197), .B2(n9009), .Y(n4582) );
	inv_1 U12150( .A(n10447), .Y(n9009) );
	nor2_1 U12151( .A(n6351), .B(n11311), .Y(n4581) );
	inv_1 U12152( .A(g8787), .Y(n11311) );
	nor2_1 U12153( .A(n6354), .B(n11418), .Y(n4580) );
	inv_1 U12154( .A(g8918), .Y(n11418) );
	o32ai_1 U12155( .A1(n8804), .A2(n6278), .A3(n9268), .B1(n11437), .B2(n11438), .Y(n4579) );
	inv_1 U12156( .A(n10928), .Y(n11438) );
	o22ai_1 U12157( .A1(n11437), .A2(n11439), .B1(n6277), .B2(n11440), .Y(n4578) );
	inv_1 U12158( .A(n10922), .Y(n11439) );
	a21oi_1 U12159( .A1(n6382), .A2(n11882), .B1(n6437), .Y(n11437) );
	o221ai_1 U12160( .A1(n7412), .A2(n8804), .B1(n6220), .B2(n9264), .C1(n11441), .Y(n4577) );
	nand3_1 U12161( .A(n6339), .B(n5883), .C(n10928), .Y(n11441) );
	nand4_1 U12162( .A(n9536), .B(n8825), .C(n11442), .D(n9264), .Y(n8804) );
	inv_1 U12163( .A(n10873), .Y(n9264) );
	nor2_1 U12164( .A(n10928), .B(n10919), .Y(n11442) );
	inv_1 U12165( .A(g7260), .Y(n8825) );
	inv_1 U12166( .A(g7245), .Y(n9536) );
	o221ai_1 U12167( .A1(n7413), .A2(n7412), .B1(n6218), .B2(n9288), .C1(n11443), .Y(n4576) );
	nand3_1 U12168( .A(n6339), .B(n5883), .C(n10922), .Y(n11443) );
	nand2_1 U12169( .A(n6337), .B(n9268), .Y(n7412) );
	o32ai_1 U12170( .A1(n6294), .A2(n10665), .A3(g10122), .B1(n6200), .B2(n6079), .Y(n4575) );
	o21ai_0 U12171( .A1(n6368), .A2(n7968), .B1(n11444), .Y(n4574) );
	nand2_1 U12172( .A(g4455), .B(n6437), .Y(n11444) );
	nand3_1 U12173( .A(g35), .B(n11440), .C(n11445), .Y(n7968) );
	mux2i_1 U12174( .A0(n10602), .A1(n9268), .S(n7413), .Y(n11445) );
	inv_1 U12175( .A(n9291), .Y(n11440) );
	nor2_1 U12176( .A(n9268), .B(n7413), .Y(n9291) );
	nand4_1 U12177( .A(n7911), .B(n8976), .C(n11446), .D(n9288), .Y(n7413) );
	inv_1 U12178( .A(n10448), .Y(n9288) );
	nor2_1 U12179( .A(n11949), .B(n10922), .Y(n11446) );
	inv_1 U12180( .A(g7257), .Y(n8976) );
	inv_1 U12181( .A(g7243), .Y(n7911) );
	o22ai_1 U12182( .A1(n6210), .A2(g23652), .B1(n6347), .B2(n9054), .Y(n4573) );
	o221ai_1 U12183( .A1(n8224), .A2(n11447), .B1(n9425), .B2(n11448), .C1( n11449), .Y(n9054) );
	a21oi_1 U12184( .A1(n11450), .A2(n8225), .B1(n6934), .Y(n11449) );
	inv_1 U12185( .A(n11451), .Y(n11450) );
	mux4_2 U12186( .A0(n10545), .A1(n10546), .A2(n7533), .A3(n9053), .S0(n8223), .S1(n11385), .X(n11451) );
	inv_1 U12187( .A(n10522), .Y(n9053) );
	inv_1 U12188( .A(n10523), .Y(n7533) );
	mux2_1 U12189( .A0(n10553), .A1(n9726), .S(n11385), .X(n11448) );
	inv_1 U12190( .A(n8630), .Y(n9425) );
	nor2_1 U12191( .A(n8225), .B(n8223), .Y(n8630) );
	inv_1 U12192( .A(n10152), .Y(n8223) );
	mux2_1 U12193( .A0(n10344), .A1(n5886), .S(n11385), .X(n11447) );
	nor4_1 U12194( .A(n10296), .B(n10235), .C(n11452), .D(n9740), .Y(n11385) );
	inv_1 U12195( .A(n9315), .Y(n11452) );
	inv_1 U12196( .A(n11142), .Y(n8224) );
	nor2_1 U12197( .A(n8225), .B(n10152), .Y(n11142) );
	inv_1 U12198( .A(n10363), .Y(n8225) );
	o22ai_1 U12199( .A1(n6210), .A2(n11453), .B1(n11454), .B2(n11430), .Y(n4572) );
	a21oi_1 U12200( .A1(n6332), .A2(n10880), .B1(n11390), .Y(n11430) );
	nor3_1 U12201( .A(n11455), .B(g20049), .C(n11429), .Y(n11454) );
	inv_1 U12202( .A(n10213), .Y(n11453) );
	nor2_1 U12203( .A(n6197), .B(n9268), .Y(n4571) );
	inv_1 U12204( .A(n10460), .Y(n9268) );
	o22ai_1 U12205( .A1(n11456), .A2(n6685), .B1(n11457), .B2(n11458), .Y(n4570) );
	inv_1 U12206( .A(n10937), .Y(n11458) );
	inv_1 U12207( .A(n11459), .Y(n11457) );
	o21ai_0 U12208( .A1(n11456), .A2(n6369), .B1(n6248), .Y(n11459) );
	inv_1 U12209( .A(n11390), .Y(n6685) );
	nor2_1 U12210( .A(n11455), .B(n6301), .Y(n11390) );
	nor3_1 U12211( .A(n11429), .B(n11965), .C(n11455), .Y(n11456) );
	inv_1 U12212( .A(n10380), .Y(n11455) );
	and2_0 U12213( .A(g4519), .B(n6383), .X(n4569) );
	and2_0 U12214( .A(g4570), .B(n6383), .X(n4568) );
	o22ai_1 U12215( .A1(n6210), .A2(n8788), .B1(n11460), .B2(n6294), .Y(n4567) );
	xnor2_1 U12216( .A(n9925), .B(n8769), .Y(n11460) );
	inv_1 U12217( .A(n10379), .Y(n8769) );
	nand4_1 U12218( .A(g11349), .B(g16718), .C(g13895), .D(g16603), .Y(n9925) );
	inv_1 U12219( .A(n10228), .Y(n8788) );
	o22ai_1 U12220( .A1(n6210), .A2(n11102), .B1(n11461), .B2(n6294), .Y(n4566) );
	xnor2_1 U12221( .A(n11147), .B(n7167), .Y(n11461) );
	inv_1 U12222( .A(n10378), .Y(n7167) );
	nand4_1 U12223( .A(g16744), .B(g16627), .C(g13926), .D(g11388), .Y(n11147) );
	inv_1 U12224( .A(n10227), .Y(n11102) );
	o22ai_1 U12225( .A1(n6209), .A2(n11462), .B1(n11463), .B2(n6295), .Y(n4565) );
	xnor2_1 U12226( .A(n9586), .B(n9135), .Y(n11463) );
	inv_1 U12227( .A(n10377), .Y(n9135) );
	nand4_1 U12228( .A(g11418), .B(g16775), .C(g16659), .D(g13966), .Y(n9586) );
	inv_1 U12229( .A(n10226), .Y(n11462) );
	o22ai_1 U12230( .A1(n6209), .A2(n11283), .B1(n11464), .B2(n6294), .Y(n4564) );
	xnor2_1 U12231( .A(n6922), .B(n6505), .Y(n11464) );
	inv_1 U12232( .A(g25219), .Y(n6505) );
	nand4_1 U12233( .A(g17674), .B(g17519), .C(g14662), .D(g12238), .Y(n6922) );
	inv_1 U12234( .A(n10225), .Y(n11283) );
	o22ai_1 U12235( .A1(n6209), .A2(n11465), .B1(n11466), .B2(n6295), .Y(n4563) );
	xnor2_1 U12236( .A(n7378), .B(n7377), .Y(n11466) );
	inv_1 U12237( .A(n10376), .Y(n7377) );
	nand4_1 U12238( .A(g17711), .B(g17580), .C(g14694), .D(g12300), .Y(n7378) );
	inv_1 U12239( .A(n10224), .Y(n11465) );
	o22ai_1 U12240( .A1(n6209), .A2(n9870), .B1(n11467), .B2(n6294), .Y(n4562) );
	xnor2_1 U12241( .A(n9166), .B(n9165), .Y(n11467) );
	inv_1 U12242( .A(n10375), .Y(n9165) );
	nand4_1 U12243( .A(g17739), .B(g17607), .C(g14738), .D(g12350), .Y(n9166) );
	inv_1 U12244( .A(n10223), .Y(n9870) );
	o22ai_1 U12245( .A1(n6209), .A2(n11468), .B1(n11469), .B2(n6294), .Y(n4561) );
	xnor2_1 U12246( .A(n9843), .B(n9842), .Y(n11469) );
	inv_1 U12247( .A(n10374), .Y(n9842) );
	nand4_1 U12248( .A(g17760), .B(g17649), .C(g14779), .D(g12422), .Y(n9843) );
	inv_1 U12249( .A(n10222), .Y(n11468) );
	o22ai_1 U12250( .A1(n6208), .A2(n9699), .B1(n11470), .B2(n6295), .Y(n4560) );
	xnor2_1 U12251( .A(n8838), .B(n7474), .Y(n11470) );
	inv_1 U12252( .A(n10373), .Y(n7474) );
	nand4_1 U12253( .A(g17778), .B(g17688), .C(g14828), .D(g12470), .Y(n8838) );
	inv_1 U12254( .A(n10221), .Y(n9699) );
	o21ai_0 U12255( .A1(n6228), .A2(n7338), .B1(n11471), .Y(n4559) );
	mux2i_1 U12256( .A0(n11472), .A1(n11473), .S(n6880), .Y(n11471) );
	nor2_1 U12257( .A(n8473), .B(n11061), .Y(n11473) );
	nand2_1 U12258( .A(n8342), .B(n6379), .Y(n8473) );
	and2_0 U12259( .A(n11061), .B(n11060), .X(n11472) );
	inv_1 U12260( .A(n7341), .Y(n11060) );
	nand2_1 U12261( .A(n10160), .B(n7340), .Y(n11061) );
	nor2_1 U12262( .A(n7334), .B(n8341), .Y(n7340) );
	nand2_1 U12263( .A(n6882), .B(n10687), .Y(n8341) );
	nor2_1 U12264( .A(n6458), .B(n10920), .Y(n6882) );
	inv_1 U12265( .A(n10668), .Y(n6458) );
	inv_1 U12266( .A(n10245), .Y(n7334) );
	inv_1 U12267( .A(n11474), .Y(n39) );
	o21ai_0 U12268( .A1(n11475), .A2(n11476), .B1(n6343), .Y(n11474) );
	o21ai_0 U12269( .A1(n5875), .A2(n6090), .B1(n11477), .Y(n11476) );
	mux2i_1 U12270( .A0(n11478), .A1(n5968), .S(n10197), .Y(n11477) );
	a21oi_1 U12271( .A1(n11479), .A2(n9068), .B1(n8105), .Y(n11478) );
	nand3_1 U12272( .A(n10973), .B(n5875), .C(n10068), .Y(n8105) );
	mux2i_1 U12273( .A0(n11480), .A1(n11481), .S(n8353), .Y(n11479) );
	inv_1 U12274( .A(n10277), .Y(n8353) );
	nor2_1 U12275( .A(n10347), .B(n11482), .Y(n11481) );
	mux2i_1 U12276( .A0(n11483), .A1(n11484), .S(n7241), .Y(n11482) );
	inv_1 U12277( .A(n10289), .Y(n7241) );
	o211ai_1 U12278( .A1(n10658), .A2(n11485), .B1(n8231), .C1(n9911), .Y( n11484) );
	inv_1 U12279( .A(n8229), .Y(n9911) );
	inv_1 U12280( .A(n9387), .Y(n8231) );
	xor2_1 U12281( .A(n6422), .B(n11486), .X(n11483) );
	a221oi_1 U12282( .A1(n10706), .A2(n9387), .B1(n10711), .B2(n8229), .C1( n11487), .Y(n11486) );
	o22ai_1 U12283( .A1(n11485), .A2(n8693), .B1(n11028), .B2(n8588), .Y(n11487) );
	inv_1 U12284( .A(n9708), .Y(n11028) );
	nor2_1 U12285( .A(n10289), .B(n6422), .Y(n11480) );
	o22ai_1 U12286( .A1(n10973), .A2(n6081), .B1(n11821), .B2(n10068), .Y( n11475) );
	inv_1 U12287( .A(n10230), .Y(n10068) );
	inv_1 U12288( .A(n10535), .Y(n10973) );
	inv_1 U12289( .A(n11488), .Y(n37) );
	o21ai_0 U12290( .A1(n11489), .A2(n11490), .B1(n6344), .Y(n11488) );
	o21ai_0 U12291( .A1(n5874), .A2(n6091), .B1(n11491), .Y(n11490) );
	mux2i_1 U12292( .A0(n11492), .A1(n6087), .S(n10198), .Y(n11491) );
	a21oi_1 U12293( .A1(n11493), .A2(n8400), .B1(n8507), .Y(n11492) );
	nand3_1 U12294( .A(n10955), .B(n5874), .C(n8760), .Y(n8507) );
	mux2i_1 U12295( .A0(n11494), .A1(n11495), .S(n9366), .Y(n11493) );
	inv_1 U12296( .A(n10278), .Y(n9366) );
	nor2_1 U12297( .A(n10348), .B(n11496), .Y(n11495) );
	mux2i_1 U12298( .A0(n11497), .A1(n11498), .S(n8220), .Y(n11496) );
	inv_1 U12299( .A(n10290), .Y(n8220) );
	o211ai_1 U12300( .A1(n10659), .A2(n11499), .B1(n8399), .C1(n8351), .Y( n11498) );
	inv_1 U12301( .A(n9837), .Y(n8351) );
	inv_1 U12302( .A(n8348), .Y(n8399) );
	xor2_1 U12303( .A(n9442), .B(n11500), .X(n11497) );
	a221oi_1 U12304( .A1(n8348), .A2(n10710), .B1(n10705), .B2(n9837), .C1( n11501), .Y(n11500) );
	o22ai_1 U12305( .A1(n11499), .A2(n7394), .B1(n9839), .B2(n10009), .Y(n11501) );
	inv_1 U12306( .A(n10707), .Y(n10009) );
	inv_1 U12307( .A(n11502), .Y(n9839) );
	nor2_1 U12308( .A(n10290), .B(n9442), .Y(n11494) );
	o22ai_1 U12309( .A1(n11787), .A2(n8760), .B1(n10955), .B2(n11503), .Y( n11489) );
	inv_1 U12310( .A(g21245), .Y(n11503) );
	inv_1 U12311( .A(n10573), .Y(n10955) );
	inv_1 U12312( .A(n10229), .Y(n8760) );
	nor2_1 U12313( .A(n8852), .B(n10920), .Y(n36) );
	inv_1 U12314( .A(n8851), .Y(n8852) );
	nor2_1 U12315( .A(n7341), .B(n11847), .Y(n8851) );
	nand2_1 U12316( .A(n6337), .B(n8342), .Y(n7341) );
	o21ai_0 U12317( .A1(n9390), .A2(n11429), .B1(g65), .Y(n8342) );
	inv_1 U12318( .A(n6684), .Y(n11429) );
	nor2_1 U12319( .A(g73), .B(g72), .Y(n6684) );
	nor2_1 U12320( .A(n9969), .B(g113), .Y(n9390) );
	inv_1 U12321( .A(n11504), .Y(n9969) );
	nor2_1 U12322( .A(n6286), .B(n10436), .Y(n22) );
	o22ai_1 U12323( .A1(n8812), .A2(n6302), .B1(n6196), .B2(n6414), .Y(n21) );
	inv_1 U12324( .A(n10682), .Y(n6414) );
	inv_1 U12325( .A(n6437), .Y(n6390) );
	nor2_1 U12326( .A(n6934), .B(n6364), .Y(n6457) );
	and4_1 U12327( .A(n11505), .B(n10682), .C(n10183), .D(n6420), .X(n8812) );
	inv_1 U12328( .A(n10177), .Y(n6420) );
	mux2i_1 U12329( .A0(n10359), .A1(n10360), .S(g84), .Y(n11505) );
	nand2_1 U12330( .A(n10236), .B(n9450), .Y(g34972) );
	xnor2_1 U12331( .A(n11506), .B(n11507), .Y(n9450) );
	xor2_1 U12332( .A(n11508), .B(n11509), .X(n11507) );
	xor2_1 U12333( .A(n11510), .B(n11511), .X(n11509) );
	xor2_1 U12334( .A(n7124), .B(n8509), .X(n11511) );
	xor2_1 U12335( .A(n9125), .B(n9571), .X(n11510) );
	xor2_1 U12336( .A(n11512), .B(n11513), .X(n11508) );
	xnor2_1 U12337( .A(n11396), .B(n11387), .Y(n11513) );
	xnor2_1 U12338( .A(n9218), .B(n8965), .Y(n11512) );
	nand2_1 U12339( .A(g55), .B(n11514), .Y(n11506) );
	nand2_1 U12340( .A(n10236), .B(n8509), .Y(g34927) );
	and2_0 U12341( .A(n11515), .B(n11516), .X(n8509) );
	a221oi_1 U12342( .A1(n11517), .A2(n10281), .B1(n10864), .B2(n11518), .C1( n11519), .Y(n11516) );
	o21ai_0 U12343( .A1(n11520), .A2(n8111), .B1(n11521), .Y(n11519) );
	inv_1 U12344( .A(n10454), .Y(n8111) );
	a221oi_1 U12345( .A1(g51), .A2(n11522), .B1(n11523), .B2(n11524), .C1( n11525), .Y(n11515) );
	o22ai_1 U12346( .A1(n6804), .A2(n11526), .B1(n6820), .B2(n11527), .Y(n11525) );
	inv_1 U12347( .A(n10455), .Y(n6820) );
	inv_1 U12348( .A(n10280), .Y(n6804) );
	nand4_1 U12349( .A(n11528), .B(n11529), .C(n11530), .D(n11531), .Y(n11524) );
	a222oi_1 U12350( .A1(g127), .A2(n11532), .B1(n10575), .B2(n11533), .C1(g92), .C2(n11534), .Y(n11531) );
	inv_1 U12351( .A(n11535), .Y(n11533) );
	a222oi_1 U12352( .A1(n11536), .A2(g21292), .B1(n10402), .B2(n11537), .C1( n10530), .C2(n11538), .Y(n11530) );
	a222oi_1 U12353( .A1(n11539), .A2(n10216), .B1(n10576), .B2(n11540), .C1( n11541), .C2(n10465), .Y(n11529) );
	a222oi_1 U12354( .A1(n11542), .A2(n10534), .B1(n11543), .B2(n10699), .C1( n10528), .C2(n11544), .Y(n11528) );
	nand2_1 U12355( .A(n10236), .B(n7124), .Y(g34925) );
	and2_0 U12356( .A(n11545), .B(n11546), .X(n7124) );
	a221oi_1 U12357( .A1(n11517), .A2(n10167), .B1(g50), .B2(n11522), .C1( n11547), .Y(n11546) );
	o21ai_0 U12358( .A1(n6728), .A2(n11548), .B1(n11521), .Y(n11547) );
	inv_1 U12359( .A(n10466), .Y(n6728) );
	a221oi_1 U12360( .A1(n11523), .A2(n11549), .B1(n11550), .B2(n10136), .C1( n11551), .Y(n11545) );
	o22ai_1 U12361( .A1(n6974), .A2(n11526), .B1(n10590), .B2(n11520), .Y( n11551) );
	inv_1 U12362( .A(n10166), .Y(n6974) );
	inv_1 U12363( .A(n10591), .Y(n10136) );
	nand4_1 U12364( .A(n11552), .B(n11553), .C(n11554), .D(n11555), .Y(n11549) );
	a222oi_1 U12365( .A1(n10384), .A2(n11537), .B1(g20652), .B2(n11534), .C1( n10476), .C2(n11532), .Y(n11555) );
	a222oi_1 U12366( .A1(n11818), .A2(n11540), .B1(n10529), .B2(n11538), .C1( n11536), .C2(n11257), .Y(n11554) );
	inv_1 U12367( .A(n10516), .Y(n11257) );
	a222oi_1 U12368( .A1(n11543), .A2(n11838), .B1(n10878), .B2(n11541), .C1( n10716), .C2(n11539), .Y(n11553) );
	a22oi_1 U12369( .A1(n10527), .A2(n11544), .B1(n11542), .B2(n10533), .Y( n11552) );
	nand2_1 U12370( .A(n10236), .B(n9571), .Y(g34923) );
	and3_1 U12371( .A(n11556), .B(n11557), .C(n11558), .X(n9571) );
	a211oi_1 U12372( .A1(n11518), .A2(n10453), .B1(n11559), .C1(n11560), .Y( n11558) );
	inv_1 U12373( .A(n11521), .Y(n11560) );
	o22ai_1 U12374( .A1(n8070), .A2(n11520), .B1(n7076), .B2(n11527), .Y(n11559) );
	inv_1 U12375( .A(n10507), .Y(n7076) );
	inv_1 U12376( .A(n10508), .Y(n8070) );
	inv_1 U12377( .A(n11548), .Y(n11518) );
	a22oi_1 U12378( .A1(g49), .A2(n11522), .B1(n11561), .B2(n10008), .Y(n11557) );
	inv_1 U12379( .A(n10659), .Y(n10008) );
	a22oi_1 U12380( .A1(n11562), .A2(n9905), .B1(n11523), .B2(n11563), .Y( n11556) );
	nand4_1 U12381( .A(n11564), .B(n11565), .C(n11566), .D(n11567), .Y(n11563) );
	a221oi_1 U12382( .A1(n10702), .A2(n11532), .B1(n11534), .B2(n10704), .C1( n11568), .Y(n11567) );
	a222oi_1 U12383( .A1(n10233), .A2(n11536), .B1(n10385), .B2(n11537), .C1( n10399), .C2(n11538), .Y(n11566) );
	a222oi_1 U12384( .A1(n10538), .A2(n11539), .B1(n10622), .B2(n11540), .C1( n10872), .C2(n11541), .Y(n11565) );
	a222oi_1 U12385( .A1(n11542), .A2(n10532), .B1(n10712), .B2(n11543), .C1( n10398), .C2(n11544), .Y(n11564) );
	inv_1 U12386( .A(n10658), .Y(n9905) );
	inv_1 U12387( .A(n11569), .Y(n11562) );
	nand2_1 U12388( .A(n10236), .B(n9125), .Y(g34921) );
	and3_1 U12389( .A(n11570), .B(n11571), .C(n11572), .X(n9125) );
	a221oi_1 U12390( .A1(n11573), .A2(n10282), .B1(n11574), .B2(n10256), .C1( n11575), .Y(n11572) );
	o221ai_1 U12391( .A1(n8588), .A2(n11569), .B1(n11526), .B2(n9248), .C1( n11521), .Y(n11575) );
	inv_1 U12392( .A(n10886), .Y(n9248) );
	inv_1 U12393( .A(n10708), .Y(n8588) );
	a22oi_1 U12394( .A1(n10885), .A2(n11517), .B1(g48), .B2(n11522), .Y(n11571) );
	a22oi_1 U12395( .A1(n10707), .A2(n11561), .B1(n11523), .B2(n11576), .Y( n11570) );
	nand4_1 U12396( .A(n11577), .B(n11578), .C(n11579), .D(n11580), .Y(n11576) );
	a221oi_1 U12397( .A1(n11537), .A2(n10551), .B1(n10443), .B2(n11532), .C1( n11568), .Y(n11580) );
	inv_1 U12398( .A(n11581), .Y(n11568) );
	a222oi_1 U12399( .A1(n10577), .A2(n11540), .B1(n10393), .B2(n11538), .C1( n11536), .C2(n11826), .Y(n11579) );
	inv_1 U12400( .A(n11582), .Y(n11540) );
	a222oi_1 U12401( .A1(n11543), .A2(n10700), .B1(n11541), .B2(n10927), .C1( n10588), .C2(n11539), .Y(n11578) );
	inv_1 U12402( .A(n11583), .Y(n11541) );
	a22oi_1 U12403( .A1(n10392), .A2(n11544), .B1(n11542), .B2(n10531), .Y( n11577) );
	inv_1 U12404( .A(n11584), .Y(n11542) );
	inv_1 U12405( .A(n11585), .Y(n11544) );
	nand2_1 U12406( .A(n10236), .B(n11387), .Y(g34919) );
	and2_0 U12407( .A(n11586), .B(n11587), .X(n11387) );
	a221oi_1 U12408( .A1(n10884), .A2(n11588), .B1(n11573), .B2(n10284), .C1( n11589), .Y(n11587) );
	o221ai_1 U12409( .A1(n11590), .A2(n8619), .B1(n8332), .B2(n11569), .C1( n11521), .Y(n11589) );
	inv_1 U12410( .A(n10706), .Y(n8332) );
	nor2_1 U12411( .A(n11591), .B(n11592), .Y(n11590) );
	o221ai_1 U12412( .A1(n11582), .A2(n8539), .B1(n6659), .B2(n11583), .C1( n11593), .Y(n11592) );
	a222oi_1 U12413( .A1(n10587), .A2(n11536), .B1(n11532), .B2(n5872), .C1( n10391), .C2(n11538), .Y(n11593) );
	inv_1 U12414( .A(n11594), .Y(n11536) );
	inv_1 U12415( .A(n10860), .Y(n6659) );
	inv_1 U12416( .A(n10578), .Y(n8539) );
	o221ai_1 U12417( .A1(n11585), .A2(n8367), .B1(n7109), .B2(n11584), .C1( n11595), .Y(n11591) );
	a222oi_1 U12418( .A1(n11543), .A2(n11774), .B1(n11537), .B2(n10926), .C1( n10437), .C2(n11539), .Y(n11595) );
	inv_1 U12419( .A(n11596), .Y(n11539) );
	inv_1 U12420( .A(n11597), .Y(n11537) );
	inv_1 U12421( .A(n11598), .Y(n11543) );
	inv_1 U12422( .A(n10390), .Y(n7109) );
	inv_1 U12423( .A(n10383), .Y(n8367) );
	a221oi_1 U12424( .A1(g47), .A2(n11522), .B1(n11561), .B2(n10705), .C1( n11599), .Y(n11586) );
	o22ai_1 U12425( .A1(n11600), .A2(n11020), .B1(n9431), .B2(n11601), .Y( n11599) );
	inv_1 U12426( .A(n10258), .Y(n9431) );
	inv_1 U12427( .A(n10883), .Y(n11020) );
	inv_1 U12428( .A(n11602), .Y(n11561) );
	nand2_1 U12429( .A(n10236), .B(n11396), .Y(g34917) );
	and3_1 U12430( .A(n11603), .B(n11604), .C(n11605), .X(n11396) );
	a221oi_1 U12431( .A1(n10889), .A2(n11517), .B1(g46), .B2(n11522), .C1( n11606), .Y(n11605) );
	o22ai_1 U12432( .A1(n7264), .A2(n11602), .B1(n8333), .B2(n11569), .Y(n11606) );
	inv_1 U12433( .A(n10711), .Y(n8333) );
	inv_1 U12434( .A(n10710), .Y(n7264) );
	a221oi_1 U12435( .A1(n10890), .A2(n11588), .B1(n11574), .B2(n10257), .C1( n11607), .Y(n11604) );
	inv_1 U12436( .A(n11526), .Y(n11588) );
	a22oi_1 U12437( .A1(n11523), .A2(n11608), .B1(n11573), .B2(n10283), .Y( n11603) );
	or4_1 U12438( .A(n11609), .B(n11610), .C(n11611), .D(n11612), .X(n11608) );
	o22ai_1 U12439( .A1(n11583), .A2(n8986), .B1(n11582), .B2(n8537), .Y(n11612) );
	inv_1 U12440( .A(n10452), .Y(n8537) );
	inv_1 U12441( .A(n10862), .Y(n8986) );
	o22ai_1 U12442( .A1(n11613), .A2(n8510), .B1(n11614), .B2(n5955), .Y(n11611) );
	inv_1 U12443( .A(n10397), .Y(n8510) );
	o22ai_1 U12444( .A1(n11584), .A2(n7588), .B1(n11585), .B2(n8372), .Y(n11610) );
	inv_1 U12445( .A(n10307), .Y(n8372) );
	inv_1 U12446( .A(n10396), .Y(n7588) );
	o22ai_1 U12447( .A1(n6748), .A2(n11598), .B1(n11596), .B2(n8343), .Y(n11609) );
	nand2_1 U12448( .A(n10236), .B(n9218), .Y(g34915) );
	and2_0 U12449( .A(n11615), .B(n11616), .X(n9218) );
	a221oi_1 U12450( .A1(n10939), .A2(n11550), .B1(g52), .B2(n11522), .C1( n11617), .Y(n11616) );
	o21ai_0 U12451( .A1(n11548), .A2(n7777), .B1(n11521), .Y(n11617) );
	nand3_1 U12452( .A(n11618), .B(n6934), .C(n11523), .Y(n11521) );
	nand4_1 U12453( .A(n11613), .B(n11585), .C(n11584), .D(n11597), .Y(n11618) );
	inv_1 U12454( .A(n10863), .Y(n7777) );
	nand2_1 U12455( .A(n11619), .B(n11620), .Y(n11548) );
	inv_1 U12456( .A(n11527), .Y(n11550) );
	a221oi_1 U12457( .A1(n10938), .A2(n11621), .B1(n11517), .B2(n10382), .C1( n11622), .Y(n11615) );
	o22ai_1 U12458( .A1(n6803), .A2(n11526), .B1(n11623), .B2(n8619), .Y(n11622) );
	nor3_1 U12459( .A(n11624), .B(n11625), .C(n11626), .Y(n11623) );
	o22ai_1 U12460( .A1(n5888), .A2(n11584), .B1(n11585), .B2(n7993), .Y(n11626) );
	inv_1 U12461( .A(n10401), .Y(n7993) );
	o221ai_1 U12462( .A1(n11535), .A2(n11214), .B1(n11597), .B2(n8043), .C1( n11581), .Y(n11625) );
	nand3_1 U12463( .A(n11627), .B(n10200), .C(n11628), .Y(n11581) );
	inv_1 U12464( .A(n10400), .Y(n8043) );
	nand3_1 U12465( .A(n11629), .B(n11630), .C(n11620), .Y(n11597) );
	inv_1 U12466( .A(n10429), .Y(n11214) );
	nand4_1 U12467( .A(n11628), .B(n11835), .C(n11631), .D(n11632), .Y(n11535) );
	o221ai_1 U12468( .A1(n11594), .A2(n11633), .B1(n11583), .B2(n8586), .C1( n11634), .Y(n11624) );
	a222oi_1 U12469( .A1(n11858), .A2(n11538), .B1(g100), .B2(n11534), .C1( n11936), .C2(n11532), .Y(n11634) );
	inv_1 U12470( .A(n11614), .Y(n11532) );
	nand4_1 U12471( .A(n11835), .B(n11620), .C(n11630), .D(n11632), .Y(n11614) );
	and3_1 U12472( .A(n11635), .B(n11632), .C(n11835), .X(n11534) );
	inv_1 U12473( .A(n11613), .Y(n11538) );
	inv_1 U12474( .A(n10698), .Y(n8586) );
	inv_1 U12475( .A(n10234), .Y(n11633) );
	inv_1 U12476( .A(n10432), .Y(n6803) );
	inv_1 U12477( .A(n11520), .Y(n11621) );
	nand2_1 U12478( .A(n10236), .B(n8965), .Y(g34913) );
	nor4_1 U12479( .A(n11607), .B(n11636), .C(n11637), .D(n11638), .Y(n8965) );
	o221ai_1 U12480( .A1(n8693), .A2(n11569), .B1(n7394), .B2(n11602), .C1( n11639), .Y(n11638) );
	a22oi_1 U12481( .A1(n10887), .A2(n11517), .B1(g45), .B2(n11522), .Y(n11639) );
	nor2_1 U12482( .A(n11523), .B(g53), .Y(n11522) );
	inv_1 U12483( .A(n11600), .Y(n11517) );
	nand2_1 U12484( .A(n11619), .B(n11640), .Y(n11600) );
	nand3_1 U12485( .A(n11640), .B(n10555), .C(n11641), .Y(n11602) );
	inv_1 U12486( .A(n10474), .Y(n7394) );
	nand3_1 U12487( .A(n10555), .B(n11620), .C(n11641), .Y(n11569) );
	inv_1 U12488( .A(n10475), .Y(n8693) );
	o22ai_1 U12489( .A1(n7455), .A2(n11642), .B1(n11643), .B2(n8619), .Y(n11637) );
	inv_1 U12490( .A(n11523), .Y(n8619) );
	nor4_1 U12491( .A(n11644), .B(n11645), .C(n11646), .D(n11647), .Y(n11643) );
	o22ai_1 U12492( .A1(n11584), .A2(n7593), .B1(n11585), .B2(n9607), .Y(n11647) );
	inv_1 U12493( .A(n10589), .Y(n9607) );
	inv_1 U12494( .A(n10394), .Y(n7593) );
	o22ai_1 U12495( .A1(n6749), .A2(n11598), .B1(n11596), .B2(n8204), .Y(n11646) );
	nand3_1 U12496( .A(n11629), .B(n11631), .C(n11628), .Y(n11596) );
	nand3_1 U12497( .A(n11629), .B(n10200), .C(n11628), .Y(n11598) );
	and4_1 U12498( .A(n10509), .B(n11648), .C(n11971), .D(n11649), .X(n11628) );
	and2_0 U12499( .A(n11970), .B(n11969), .X(n11649) );
	o22ai_1 U12500( .A1(n11583), .A2(n9897), .B1(n11582), .B2(n7296), .Y(n11645) );
	inv_1 U12501( .A(n10451), .Y(n7296) );
	nand3_1 U12502( .A(n11620), .B(n11629), .C(n10509), .Y(n11582) );
	inv_1 U12503( .A(n10861), .Y(n9897) );
	nand3_1 U12504( .A(n11640), .B(n11629), .C(n10509), .Y(n11583) );
	o22ai_1 U12505( .A1(n7041), .A2(n11594), .B1(n11613), .B2(n8209), .Y(n11644) );
	inv_1 U12506( .A(n10395), .Y(n8209) );
	nand3_1 U12507( .A(n11629), .B(n11630), .C(n11640), .Y(n11594) );
	inv_1 U12508( .A(n10871), .Y(n7041) );
	inv_1 U12509( .A(n11573), .Y(n11642) );
	nor2_1 U12510( .A(n11527), .B(n10507), .Y(n11573) );
	nand3_1 U12511( .A(n11650), .B(n11620), .C(n11523), .Y(n11527) );
	and3_1 U12512( .A(n11651), .B(n11648), .C(n10200), .X(n11620) );
	inv_1 U12513( .A(n10306), .Y(n7455) );
	o22ai_1 U12514( .A1(n11526), .A2(n10102), .B1(n6799), .B2(n11601), .Y( n11636) );
	inv_1 U12515( .A(n11574), .Y(n11601) );
	nor2_1 U12516( .A(n11520), .B(n10508), .Y(n11574) );
	nand3_1 U12517( .A(n11640), .B(n11632), .C(n11641), .Y(n11520) );
	and3_1 U12518( .A(n11523), .B(n11630), .C(n11835), .X(n11641) );
	inv_1 U12519( .A(n10285), .Y(n6799) );
	inv_1 U12520( .A(n10888), .Y(n10102) );
	nand3_1 U12521( .A(n10343), .B(n11652), .C(n11619), .Y(n11526) );
	and3_1 U12522( .A(n11523), .B(n11627), .C(n10509), .X(n11619) );
	and3_1 U12523( .A(n11653), .B(n6934), .C(n11523), .X(n11607) );
	nor4_1 U12524( .A(g53), .B(n11514), .C(n10232), .D(g57), .Y(n11523) );
	nand2_1 U12525( .A(g54), .B(n11654), .Y(n11514) );
	inv_1 U12526( .A(g56), .Y(n11654) );
	nand3_1 U12527( .A(n11585), .B(n11584), .C(n11613), .Y(n11653) );
	nand2_1 U12528( .A(n11635), .B(n11629), .Y(n11613) );
	nor2_1 U12529( .A(n10555), .B(n11835), .Y(n11629) );
	and4_1 U12530( .A(n10343), .B(n10200), .C(n11651), .D(n11630), .X(n11635) );
	nand3_1 U12531( .A(n11652), .B(n11650), .C(n10343), .Y(n11584) );
	nand2_1 U12532( .A(n11640), .B(n11650), .Y(n11585) );
	and2_0 U12533( .A(n11627), .B(n11630), .X(n11650) );
	inv_1 U12534( .A(n10509), .Y(n11630) );
	nor2_1 U12535( .A(n11632), .B(n11835), .Y(n11627) );
	inv_1 U12536( .A(n10555), .Y(n11632) );
	and2_0 U12537( .A(n11652), .B(n11648), .X(n11640) );
	inv_1 U12538( .A(n10343), .Y(n11648) );
	and2_0 U12539( .A(n11651), .B(n11631), .X(n11652) );
	inv_1 U12540( .A(n10200), .Y(n11631) );
	nor3_1 U12541( .A(n11970), .B(n11969), .C(n11971), .Y(n11651) );
	a21oi_1 U12542( .A1(n11064), .A2(n11168), .B1(n5956), .Y(g34839) );
	inv_1 U12543( .A(n10667), .Y(n11168) );
	a21oi_1 U12544( .A1(n11843), .A2(n11655), .B1(n8489), .Y(g33894) );
	inv_1 U12545( .A(n10671), .Y(n8489) );
	nor4_1 U12546( .A(n10592), .B(n10362), .C(n10182), .D(n11656), .Y(g31521) );
	nor3_1 U12547( .A(n11657), .B(n10356), .C(n10328), .Y(n11656) );
	and4_1 U12548( .A(n8829), .B(n8817), .C(n10858), .D(n10162), .X(n11657) );
	inv_1 U12549( .A(n10288), .Y(n8829) );
	nand2_1 U12550( .A(n11658), .B(n8635), .Y(g34425) );
	mux2_1 U12551( .A0(n11659), .A1(n11660), .S(n6880), .X(n8635) );
	inv_1 U12552( .A(n10255), .Y(n6880) );
	a221oi_1 U12553( .A1(n9389), .A2(n6607), .B1(n7687), .B2(n7049), .C1(n11661), .Y(n11660) );
	o22ai_1 U12554( .A1(n8627), .A2(n11662), .B1(n11663), .B2(n8536), .Y(n11661) );
	nand2_1 U12555( .A(n10365), .B(n10191), .Y(n8536) );
	inv_1 U12556( .A(n9373), .Y(n11662) );
	and2_0 U12557( .A(n10194), .B(n10368), .X(n7687) );
	inv_1 U12558( .A(n7198), .Y(n6607) );
	nand2_1 U12559( .A(n11917), .B(n10327), .Y(n7198) );
	a221oi_1 U12560( .A1(n9064), .A2(n8262), .B1(n8903), .B2(n9373), .C1(n11664), .Y(n11659) );
	inv_1 U12561( .A(n11665), .Y(n11664) );
	a22oi_1 U12562( .A1(n7049), .A2(n8396), .B1(n9389), .B2(n9145), .Y(n11665) );
	nor2_1 U12563( .A(n9213), .B(n9910), .Y(n9145) );
	inv_1 U12564( .A(n10195), .Y(n9910) );
	inv_1 U12565( .A(n10369), .Y(n9213) );
	and2_0 U12566( .A(n10974), .B(n10160), .X(n9389) );
	nor2_1 U12567( .A(n10109), .B(n10145), .Y(n8396) );
	inv_1 U12568( .A(n10192), .Y(n10145) );
	inv_1 U12569( .A(n10366), .Y(n10109) );
	nor2_1 U12570( .A(n11666), .B(n7338), .Y(n7049) );
	nor2_1 U12571( .A(n11666), .B(n10160), .Y(n9373) );
	nor2_1 U12572( .A(n9876), .B(n8408), .Y(n8903) );
	inv_1 U12573( .A(n10367), .Y(n8408) );
	inv_1 U12574( .A(n10193), .Y(n9876) );
	inv_1 U12575( .A(n11663), .Y(n8262) );
	nand2_1 U12576( .A(n10974), .B(n7338), .Y(n11663) );
	inv_1 U12577( .A(n10160), .Y(n7338) );
	nor2_1 U12578( .A(n11108), .B(n6833), .Y(n9064) );
	inv_1 U12579( .A(n10370), .Y(n6833) );
	inv_1 U12580( .A(n10196), .Y(n11108) );
	o211ai_1 U12581( .A1(n11667), .A2(n11668), .B1(n11669), .C1(n7300), .Y( g34383) );
	and4_1 U12582( .A(n11670), .B(n11671), .C(n11672), .D(n11673), .X(n7300) );
	nor4_1 U12583( .A(n11674), .B(n11675), .C(n11676), .D(n11677), .Y(n11673) );
	nor3_1 U12584( .A(n7895), .B(n10253), .C(n7891), .Y(n11677) );
	inv_1 U12585( .A(n10263), .Y(n7895) );
	nor3_1 U12586( .A(n6573), .B(n10252), .C(n9307), .Y(n11676) );
	inv_1 U12587( .A(n10262), .Y(n6573) );
	nor3_1 U12588( .A(n7449), .B(n10254), .C(n9091), .Y(n11675) );
	inv_1 U12589( .A(n10264), .Y(n7449) );
	nor3_1 U12590( .A(n7038), .B(n10249), .C(n7034), .Y(n11674) );
	inv_1 U12591( .A(n10259), .Y(n7038) );
	a22oi_1 U12592( .A1(n9008), .A2(n6562), .B1(g25259), .B2(n7599), .Y(n11672) );
	inv_1 U12593( .A(n11678), .Y(n7599) );
	nor2_1 U12594( .A(n8014), .B(n10287), .Y(n6562) );
	inv_1 U12595( .A(n10265), .Y(n8014) );
	inv_1 U12596( .A(n11679), .Y(n9008) );
	nand3_1 U12597( .A(n8089), .B(n7089), .C(n10260), .Y(n11671) );
	inv_1 U12598( .A(n10250), .Y(n7089) );
	inv_1 U12599( .A(n8092), .Y(n8089) );
	nand3_1 U12600( .A(n8881), .B(n7430), .C(n10261), .Y(n11670) );
	inv_1 U12601( .A(n10251), .Y(n7430) );
	inv_1 U12602( .A(n8884), .Y(n8881) );
	nand4_1 U12603( .A(n9091), .B(n11679), .C(n7891), .D(n8884), .Y(n11668) );
	nand3_1 U12604( .A(n8525), .B(n8960), .C(n11680), .Y(n8884) );
	nand3_1 U12605( .A(n10161), .B(n11655), .C(n10293), .Y(n7891) );
	nand3_1 U12606( .A(n10161), .B(n8960), .C(n11680), .Y(n11679) );
	nand3_1 U12607( .A(n11655), .B(n8525), .C(n10293), .Y(n9091) );
	nand4_1 U12608( .A(n11678), .B(n8092), .C(n7034), .D(n9307), .Y(n11667) );
	nand3_1 U12609( .A(n11655), .B(n8960), .C(n10161), .Y(n9307) );
	nand3_1 U12610( .A(n11680), .B(n10161), .C(n10293), .Y(n7034) );
	nand3_1 U12611( .A(n11680), .B(n8525), .C(n10293), .Y(n8092) );
	and3_1 U12612( .A(n11681), .B(n11682), .C(n10371), .X(n11680) );
	nand3_1 U12613( .A(n8525), .B(n8960), .C(n11655), .Y(n11678) );
	and3_1 U12614( .A(n11682), .B(n7414), .C(n11681), .X(n11655) );
	xnor2_1 U12615( .A(n10330), .B(g73), .Y(n11681) );
	inv_1 U12616( .A(n10371), .Y(n7414) );
	xnor2_1 U12617( .A(n10199), .B(g72), .Y(n11682) );
	inv_1 U12618( .A(n10293), .Y(n8960) );
	inv_1 U12619( .A(n10161), .Y(n8525) );
	nand2_1 U12620( .A(n8490), .B(n11658), .Y(g34221) );
	inv_1 U12621( .A(n11683), .Y(n11658) );
	o21ai_0 U12622( .A1(n11064), .A2(n10974), .B1(n11669), .Y(n11683) );
	inv_1 U12623( .A(n11666), .Y(n11064) );
	inv_1 U12624( .A(n11684), .Y(n8490) );
	o32ai_1 U12625( .A1(n9365), .A2(n11666), .A3(n6840), .B1(n8528), .B2(n11685), .Y(n11684) );
	nand2_1 U12626( .A(n7825), .B(n10974), .Y(n11685) );
	and2_0 U12627( .A(n11686), .B(n10361), .X(n10974) );
	inv_1 U12628( .A(n8106), .Y(n7825) );
	nand2_1 U12629( .A(n7549), .B(n11961), .Y(n8106) );
	nor2_1 U12630( .A(n7826), .B(n7822), .Y(n7549) );
	inv_1 U12631( .A(n10190), .Y(n7822) );
	nand2_1 U12632( .A(n10197), .B(n10462), .Y(n7826) );
	inv_1 U12633( .A(n8532), .Y(n8528) );
	nor2_1 U12634( .A(n9068), .B(n11485), .Y(n8532) );
	inv_1 U12635( .A(n9913), .Y(n11485) );
	nand3_1 U12636( .A(n10289), .B(n8173), .C(n10277), .Y(n9068) );
	inv_1 U12637( .A(n10347), .Y(n8173) );
	inv_1 U12638( .A(n6842), .Y(n6840) );
	nor2_1 U12639( .A(n11499), .B(n8400), .Y(n6842) );
	nand3_1 U12640( .A(n10290), .B(n9454), .C(n10278), .Y(n8400) );
	inv_1 U12641( .A(n10348), .Y(n9454) );
	inv_1 U12642( .A(n11119), .Y(n11499) );
	nand2_1 U12643( .A(n11686), .B(n7612), .Y(n11666) );
	inv_1 U12644( .A(n10361), .Y(n7612) );
	and2_0 U12645( .A(n11687), .B(n11688), .X(n11686) );
	xnor2_1 U12646( .A(g72), .B(n10246), .Y(n11688) );
	xnor2_1 U12647( .A(n10279), .B(g73), .Y(n11687) );
	nand2_1 U12648( .A(n11898), .B(n8989), .Y(n9365) );
	and2_0 U12649( .A(n10189), .B(n6596), .X(n8989) );
	and2_0 U12650( .A(n10198), .B(n10461), .X(n6596) );
	o211ai_1 U12651( .A1(n11689), .A2(n11690), .B1(n11669), .C1(n9517), .Y( g34201) );
	nor4_1 U12652( .A(n11691), .B(n11692), .C(n11693), .D(n11694), .Y(n9517) );
	o22ai_1 U12653( .A1(n9339), .A2(n9076), .B1(n6743), .B2(n7090), .Y(n11694) );
	inv_1 U12654( .A(n7087), .Y(n7090) );
	nor2_1 U12655( .A(n6741), .B(n10333), .Y(n7087) );
	inv_1 U12656( .A(n10172), .Y(n6741) );
	inv_1 U12657( .A(n9074), .Y(n9076) );
	nor2_1 U12658( .A(n8238), .B(n10334), .Y(n9074) );
	inv_1 U12659( .A(n10173), .Y(n8238) );
	o22ai_1 U12660( .A1(n7835), .A2(n9428), .B1(n9276), .B2(n9043), .Y(n11693) );
	inv_1 U12661( .A(n7627), .Y(n9276) );
	nor2_1 U12662( .A(n9042), .B(n10331), .Y(n7627) );
	inv_1 U12663( .A(n10299), .Y(n9042) );
	inv_1 U12664( .A(n7926), .Y(n9428) );
	nor2_1 U12665( .A(n7832), .B(n10332), .Y(n7926) );
	inv_1 U12666( .A(n10171), .Y(n7832) );
	o22ai_1 U12667( .A1(n9598), .A2(n10063), .B1(n10090), .B2(n7955), .Y(n11692) );
	inv_1 U12668( .A(n7359), .Y(n7955) );
	nor2_1 U12669( .A(n7793), .B(n10337), .Y(n7359) );
	inv_1 U12670( .A(n10176), .Y(n7793) );
	inv_1 U12671( .A(g25167), .Y(n10063) );
	o22ai_1 U12672( .A1(n7223), .A2(n7724), .B1(n8316), .B2(n7579), .Y(n11691) );
	inv_1 U12673( .A(n6850), .Y(n8316) );
	nor2_1 U12674( .A(n7100), .B(n10335), .Y(n6850) );
	inv_1 U12675( .A(n10174), .Y(n7100) );
	inv_1 U12676( .A(n7219), .Y(n7223) );
	nor2_1 U12677( .A(n7722), .B(n10336), .Y(n7219) );
	inv_1 U12678( .A(n10175), .Y(n7722) );
	nand4_1 U12679( .A(n9043), .B(n7724), .C(n9339), .D(n7579), .Y(n11690) );
	nand3_1 U12680( .A(n10235), .B(n5882), .C(n11695), .Y(n7579) );
	nand2_1 U12681( .A(n11696), .B(n6391), .Y(n9339) );
	nand3_1 U12682( .A(n6391), .B(n5882), .C(n11695), .Y(n7724) );
	nand3_1 U12683( .A(n11963), .B(n10235), .C(n11695), .Y(n9043) );
	nand4_1 U12684( .A(n7835), .B(n6743), .C(n10090), .D(n9598), .Y(n11689) );
	nand3_1 U12685( .A(n9315), .B(n6391), .C(n11697), .Y(n9598) );
	nand3_1 U12686( .A(n9315), .B(n10235), .C(n11697), .Y(n10090) );
	nor2_1 U12687( .A(n11963), .B(n10552), .Y(n9315) );
	nand2_1 U12688( .A(n11696), .B(n10235), .Y(n6743) );
	and3_1 U12689( .A(n11697), .B(n6397), .C(n11963), .X(n11696) );
	inv_1 U12690( .A(n10552), .Y(n6397) );
	nand3_1 U12691( .A(n11963), .B(n6391), .C(n11695), .Y(n7835) );
	and2_0 U12692( .A(n11697), .B(n10552), .X(n11695) );
	and2_0 U12693( .A(n11698), .B(n11699), .X(n11697) );
	xnor2_1 U12694( .A(n10424), .B(g72), .Y(n11699) );
	xnor2_1 U12695( .A(n10435), .B(g73), .Y(n11698) );
	inv_1 U12696( .A(n10235), .Y(n6391) );
	nand4_1 U12697( .A(n6422), .B(g8283), .C(g8403), .D(n11504), .Y(g33935) );
	a221oi_1 U12698( .A1(n9387), .A2(n11916), .B1(n8229), .B2(n11905), .C1( n11700), .Y(n6422) );
	inv_1 U12699( .A(n11701), .Y(n11700) );
	a22oi_1 U12700( .A1(n11910), .A2(n9708), .B1(n11810), .B2(n9913), .Y(n11701) );
	nor2_1 U12701( .A(n7238), .B(n8226), .Y(n9913) );
	nor2_1 U12702( .A(n10181), .B(n10305), .Y(n9708) );
	nor2_1 U12703( .A(n8226), .B(n10305), .Y(n8229) );
	inv_1 U12704( .A(n10181), .Y(n8226) );
	nor2_1 U12705( .A(n7238), .B(n10181), .Y(n9387) );
	inv_1 U12706( .A(n10305), .Y(n7238) );
	nand3_1 U12707( .A(n11504), .B(n11394), .C(n11779), .Y(g33874) );
	inv_1 U12708( .A(g18881), .Y(n11394) );
	nand3_1 U12709( .A(n11167), .B(n9718), .C(n11669), .Y(g33659) );
	and2_0 U12710( .A(g113), .B(n11504), .X(n11669) );
	mux2_1 U12711( .A0(n11702), .A1(n11703), .S(n10288), .X(n9718) );
	a222oi_1 U12712( .A1(n11704), .A2(n10342), .B1(n9119), .B2(n8385), .C1( n8817), .C2(n6690), .Y(n11703) );
	nor2_1 U12713( .A(n7407), .B(n7353), .Y(n6690) );
	nand2_1 U12714( .A(n10349), .B(n10202), .Y(n7353) );
	inv_1 U12715( .A(n10153), .Y(n7407) );
	nor2_1 U12716( .A(n7186), .B(n6674), .Y(n8385) );
	inv_1 U12717( .A(n10164), .Y(n6674) );
	nand2_1 U12718( .A(n10352), .B(n10201), .Y(n7186) );
	mux2i_1 U12719( .A0(n6653), .A1(n9017), .S(n9116), .Y(n11704) );
	inv_1 U12720( .A(n6663), .Y(n9017) );
	nor2_1 U12721( .A(n7071), .B(n6482), .Y(n6663) );
	inv_1 U12722( .A(n10158), .Y(n6482) );
	nand2_1 U12723( .A(n10513), .B(n10209), .Y(n7071) );
	inv_1 U12724( .A(n7010), .Y(n6653) );
	nor2_1 U12725( .A(n6994), .B(n7875), .Y(n7010) );
	nand2_1 U12726( .A(n10512), .B(n10208), .Y(n7875) );
	inv_1 U12727( .A(n10157), .Y(n6994) );
	a222oi_1 U12728( .A1(n11705), .A2(n10342), .B1(n9119), .B2(n6427), .C1( n8817), .C2(g26801), .Y(n11702) );
	nor2_1 U12729( .A(n10342), .B(n10163), .Y(n8817) );
	nor2_1 U12730( .A(n8185), .B(n6888), .Y(n6427) );
	nand2_1 U12731( .A(n10350), .B(n10203), .Y(n6888) );
	inv_1 U12732( .A(n10156), .Y(n8185) );
	nor2_1 U12733( .A(n9116), .B(n10342), .Y(n9119) );
	mux2i_1 U12734( .A0(n9478), .A1(n6864), .S(n9116), .Y(n11705) );
	inv_1 U12735( .A(n10163), .Y(n9116) );
	inv_1 U12736( .A(n7248), .Y(n6864) );
	nor2_1 U12737( .A(n7228), .B(n8069), .Y(n7248) );
	nand2_1 U12738( .A(n10511), .B(n10207), .Y(n8069) );
	inv_1 U12739( .A(n10155), .Y(n7228) );
	inv_1 U12740( .A(n9282), .Y(n9478) );
	nor2_1 U12741( .A(n9287), .B(n8169), .Y(n9282) );
	inv_1 U12742( .A(n10154), .Y(n8169) );
	nand2_1 U12743( .A(n10510), .B(n10206), .Y(n9287) );
	inv_1 U12744( .A(n9719), .Y(n11167) );
	nand2_1 U12745( .A(n11706), .B(n11707), .Y(n9719) );
	xnor2_1 U12746( .A(n10425), .B(g72), .Y(n11707) );
	xnor2_1 U12747( .A(n10434), .B(g73), .Y(n11706) );
	nand4_1 U12748( .A(g8235), .B(n9442), .C(g8353), .D(n11504), .Y(g33636) );
	nand2_1 U12749( .A(n11230), .B(n11708), .Y(n11504) );
	nand2_1 U12750( .A(g99), .B(n10704), .Y(n11708) );
	inv_1 U12751( .A(g134), .Y(n11230) );
	a221oi_1 U12752( .A1(n8348), .A2(n11890), .B1(n9837), .B2(n11967), .C1( n11709), .Y(n9442) );
	inv_1 U12753( .A(n11710), .Y(n11709) );
	a22oi_1 U12754( .A1(n11941), .A2(n11502), .B1(n11801), .B2(n11119), .Y( n11710) );
	nor2_1 U12755( .A(n8345), .B(n8217), .Y(n11119) );
	nor2_1 U12756( .A(n8217), .B(n10403), .Y(n9837) );
	inv_1 U12757( .A(n10169), .Y(n8217) );
	nor2_1 U12758( .A(n8345), .B(n10169), .Y(n8348) );
	inv_1 U12759( .A(n10403), .Y(n8345) );
	o221ai_1 U12760( .A1(n10525), .A2(n6913), .B1(n10524), .B2(n9740), .C1( n11711), .Y(g33435) );
	a22oi_1 U12761( .A1(n9730), .A2(n5885), .B1(n9903), .B2(n9645), .Y(n11711) );
	inv_1 U12762( .A(n10673), .Y(n9645) );
	o221ai_1 U12763( .A1(n10523), .A2(n6913), .B1(n10522), .B2(n9740), .C1( n11712), .Y(g33079) );
	a22oi_1 U12764( .A1(n9730), .A2(n5886), .B1(n9903), .B2(n9726), .Y(n11712) );
	inv_1 U12765( .A(n10672), .Y(n9726) );
	nor2_1 U12766( .A(n6633), .B(n8365), .Y(n9903) );
	nor2_1 U12767( .A(n6633), .B(n10244), .Y(n9730) );
	inv_1 U12768( .A(n10338), .Y(n6633) );
	inv_1 U12769( .A(n7537), .Y(n9740) );
	nor2_1 U12770( .A(n10338), .B(n10244), .Y(n7537) );
	inv_1 U12771( .A(n9775), .Y(n6913) );
	nor2_1 U12772( .A(n8365), .B(n10338), .Y(n9775) );
	inv_1 U12773( .A(n10244), .Y(n8365) );
	nor2_1 U12774( .A(n8614), .B(n7570), .Y(g26801) );
	nand2_1 U12775( .A(n10351), .B(n10204), .Y(n7570) );
	inv_1 U12776( .A(n10159), .Y(n8614) );
	nor4_1 U12777( .A(n11713), .B(n11714), .C(n11715), .D(n11716), .Y(g32185) );
	o22ai_1 U12778( .A1(n5906), .A2(n9479), .B1(n6496), .B2(n6556), .Y(n11716) );
	inv_1 U12779( .A(n10216), .Y(n6556) );
	inv_1 U12780( .A(n10699), .Y(n6496) );
	inv_1 U12781( .A(n10716), .Y(n9479) );
	nor2_1 U12782( .A(n7404), .B(n8661), .Y(n11715) );
	inv_1 U12783( .A(n10538), .Y(n8661) );
	inv_1 U12784( .A(n10712), .Y(n7404) );
	o22ai_1 U12785( .A1(n6748), .A2(n8343), .B1(n5897), .B2(n10081), .Y(n11714) );
	inv_1 U12786( .A(n10437), .Y(n10081) );
	inv_1 U12787( .A(n10438), .Y(n8343) );
	inv_1 U12788( .A(n10709), .Y(n6748) );
	o22ai_1 U12789( .A1(n6937), .A2(n10975), .B1(n6749), .B2(n8204), .Y(n11713) );
	inv_1 U12790( .A(n10444), .Y(n8204) );
	inv_1 U12791( .A(n10701), .Y(n6749) );
	inv_1 U12792( .A(n10588), .Y(n10975) );
	inv_1 U12793( .A(n10700), .Y(n6937) );
	nor2_1 U12794( .A(n6707), .B(n10292), .Y(g25167) );
	inv_1 U12795( .A(n10301), .Y(n6707) );
	nor2_1 U12796( .A(n7305), .B(n10286), .Y(g25259) );
	inv_1 U12797( .A(n10266), .Y(n7305) );
	o21ai_0 U12798( .A1(n10980), .A2(n11717), .B1(n11718), .Y(g31793) );
	o211ai_1 U12799( .A1(n11719), .A2(n11720), .B1(n8541), .C1(n8540), .Y( n11718) );
	a21oi_1 U12800( .A1(n11802), .A2(g35), .B1(n11721), .Y(n11720) );
	a211oi_1 U12801( .A1(n11722), .A2(n11721), .B1(n10656), .C1(n10231), .Y( n11719) );
	o221ai_1 U12802( .A1(n11723), .A2(n11724), .B1(n5947), .B2(n5879), .C1( n11725), .Y(n11722) );
	a21oi_1 U12803( .A1(n11918), .A2(n11768), .B1(n11802), .Y(n11725) );
	o22ai_1 U12804( .A1(n8541), .A2(n8540), .B1(n5878), .B2(n5946), .Y(n11717) );
	o21ai_0 U12805( .A1(n11860), .A2(n11760), .B1(g35), .Y(n8540) );
	inv_1 U12806( .A(n6472), .Y(n8541) );
	nor2_1 U12807( .A(n6038), .B(n6934), .Y(n6472) );
	inv_1 U12808( .A(n8542), .Y(n10980) );
	nor4_1 U12809( .A(n11721), .B(n10231), .C(n10656), .D(n11802), .Y(n8542) );
	o21ai_0 U12810( .A1(n11723), .A2(n6934), .B1(n11724), .Y(n11721) );
	o21ai_0 U12811( .A1(n11918), .A2(n11768), .B1(g35), .Y(n11724) );
	nor2_1 U12812( .A(n11790), .B(n11798), .Y(n11723) );
	nand2_1 U12813( .A(g113), .B(n10702), .Y(g31665) );
	nand2_1 U12814( .A(g113), .B(n10476), .Y(g31656) );
	inv_1 U12815( .A(n10704), .Y(g23002) );
	inv_1 U12816( .A(n8622), .Y(g28753) );
	nand2_1 U12817( .A(n10573), .B(n11726), .Y(n8622) );
	nand3_1 U12818( .A(n11502), .B(n9838), .C(n11941), .Y(n11726) );
	and4_1 U12819( .A(n11898), .B(n10189), .C(n10290), .D(n11727), .X(n9838) );
	nor3_1 U12820( .A(n6592), .B(n10348), .C(n10278), .Y(n11727) );
	inv_1 U12821( .A(n10461), .Y(n6592) );
	nor2_1 U12822( .A(n10169), .B(n10403), .Y(n11502) );
	nand3_1 U12823( .A(n9362), .B(n9481), .C(g35), .Y(g28042) );
	inv_1 U12824( .A(n10467), .Y(n9481) );
	inv_1 U12825( .A(n10186), .Y(n9362) );
	nand3_1 U12826( .A(n8113), .B(n6822), .C(g35), .Y(g28041) );
	inv_1 U12827( .A(n8153), .Y(n6822) );
	nor2_1 U12828( .A(n8103), .B(n11364), .Y(n8153) );
	nor2_1 U12829( .A(n10557), .B(n10518), .Y(n11364) );
	inv_1 U12830( .A(n10412), .Y(n8103) );
	inv_1 U12831( .A(n10060), .Y(n8113) );
	nor2_1 U12832( .A(n7277), .B(n11367), .Y(n10060) );
	nor2_1 U12833( .A(n10556), .B(n10517), .Y(n11367) );
	inv_1 U12834( .A(n10411), .Y(n7277) );
	nand2_1 U12835( .A(n9927), .B(n11728), .Y(g28030) );
	nand3_1 U12836( .A(n6873), .B(n9928), .C(n11729), .Y(n11728) );
	o22ai_1 U12837( .A1(n11730), .A2(n11731), .B1(n11732), .B2(n11733), .Y( n11729) );
	a22oi_1 U12838( .A1(n11734), .A2(n11735), .B1(n11736), .B2(n11737), .Y( n11733) );
	o32ai_1 U12839( .A1(n11738), .A2(n10610), .A3(n10217), .B1(n11739), .B2( n11740), .Y(n11737) );
	o22ai_1 U12840( .A1(n11741), .A2(n11742), .B1(n11743), .B2(n11744), .Y( n11738) );
	o21ai_0 U12841( .A1(n11765), .A2(n10869), .B1(n11745), .Y(n11735) );
	inv_1 U12842( .A(n11730), .Y(n11734) );
	inv_1 U12843( .A(n10657), .Y(n9928) );
	inv_1 U12844( .A(n10184), .Y(n6873) );
	or3_1 U12845( .A(n11730), .B(n11732), .C(n11731), .X(n9927) );
	inv_1 U12846( .A(n11736), .Y(n11731) );
	nor2_1 U12847( .A(n11746), .B(n11745), .Y(n11736) );
	a21oi_1 U12848( .A1(n6040), .A2(n9392), .B1(n6934), .Y(n11745) );
	inv_1 U12849( .A(n10868), .Y(n9392) );
	a21oi_1 U12850( .A1(n6039), .A2(n8033), .B1(n6934), .Y(n11746) );
	inv_1 U12851( .A(n10869), .Y(n8033) );
	a21oi_1 U12852( .A1(n6041), .A2(n7179), .B1(n6934), .Y(n11732) );
	inv_1 U12853( .A(n10867), .Y(n7179) );
	o21ai_0 U12854( .A1(n11747), .A2(n6934), .B1(n11743), .Y(n11730) );
	inv_1 U12855( .A(n11740), .Y(n11743) );
	o21ai_0 U12856( .A1(n11741), .A2(n6934), .B1(n11742), .Y(n11740) );
	o21ai_0 U12857( .A1(n11887), .A2(n10866), .B1(g35), .Y(n11742) );
	nor2_1 U12858( .A(n11888), .B(n10865), .Y(n11741) );
	inv_1 U12859( .A(g35), .Y(n6934) );
	nor3_1 U12860( .A(n11739), .B(n10610), .C(n10217), .Y(n11747) );
	inv_1 U12861( .A(n11744), .Y(n11739) );
	nor2_1 U12862( .A(n10661), .B(n10212), .Y(n11744) );
	inv_1 U12863( .A(n11748), .Y(g27831) );
	o21ai_0 U12864( .A1(n6404), .A2(n11029), .B1(g17291), .Y(n11748) );
	nand4_1 U12865( .A(n10179), .B(n7732), .C(n10346), .D(n11749), .Y(n11029) );
	nor3_1 U12866( .A(n10405), .B(n10471), .C(n10446), .Y(n11749) );
	inv_1 U12867( .A(n10215), .Y(n7732) );
	inv_1 U12868( .A(n6552), .Y(n6404) );
	nor2_1 U12869( .A(n6406), .B(n11957), .Y(n6552) );
	inv_1 U12870( .A(n10248), .Y(n6406) );
	nand2_1 U12871( .A(n8664), .B(n8663), .Y(g26877) );
	nand2_1 U12872( .A(n11750), .B(n11751), .Y(n8663) );
	nor4_1 U12873( .A(n11794), .B(n11795), .C(n11836), .D(n11849), .Y(n11751) );
	nor4_1 U12874( .A(n11866), .B(n11867), .C(n11868), .D(n11869), .Y(n11750) );
	inv_1 U12875( .A(n11752), .Y(n8664) );
	o21ai_0 U12876( .A1(n11753), .A2(n11754), .B1(g35), .Y(n11752) );
	nand4_1 U12877( .A(n5918), .B(n5862), .C(n5867), .D(n5873), .Y(n11754) );
	nand4_1 U12878( .A(n5969), .B(n5866), .C(n5871), .D(n5881), .Y(n11753) );
	nand3_1 U12879( .A(n7299), .B(n7298), .C(g35), .Y(g26876) );
	nand2_1 U12880( .A(n11755), .B(n11756), .Y(n7298) );
	nor4_1 U12881( .A(n11920), .B(n11921), .C(n11922), .D(n11923), .Y(n11756) );
	nor4_1 U12882( .A(n11924), .B(n11925), .C(n11926), .D(n11927), .Y(n11755) );
	nand2_1 U12883( .A(n11757), .B(n11758), .Y(n7299) );
	nor4_1 U12884( .A(n11928), .B(n11929), .C(n11930), .D(n11931), .Y(n11758) );
	nor4_1 U12885( .A(n11932), .B(n11933), .C(n11934), .D(n11935), .Y(n11757) );
	nand2_1 U12886( .A(n9551), .B(n9550), .Y(g26875) );
	nand4_1 U12887( .A(n5942), .B(n5863), .C(n5868), .D(n5876), .Y(n9550) );
	inv_1 U12888( .A(n10981), .Y(n9551) );
	nand2_1 U12889( .A(g35), .B(n11759), .Y(n10981) );
	nand4_1 U12890( .A(n5943), .B(n5864), .C(n5869), .D(n5877), .Y(n11759) );
	inv_1 U12891( .A(n8627), .Y(g25114) );
	nand2_1 U12892( .A(n10381), .B(n10188), .Y(n8627) );
	inv_1 U12893( .A(g21292), .Y(g23612) );
	nor2_1 U12894( .A(n11944), .B(n10236), .Y(g23190) );
	nor2_1 U12895( .A(g35), .B(n20311), .Y(g21727) );
	inv_1 U12896( .A(g5), .Y(g12833) );
	dfrtp_1 troj0_0_counter_reg_0_( .D(troj0_0_n3), .CLK(CLK), .RESET_B(troj0_0_N5), .Q(troj0_0_counter_0_) );
	dfrtp_1 troj0_0_counter_reg_1_( .D(troj0_0_n2), .CLK(CLK), .RESET_B(troj0_0_N5), .Q(troj0_0_counter_1_) );
	dfrtp_1 troj0_0_counter_reg_2_( .D(troj0_0_n1), .CLK(CLK), .RESET_B(troj0_0_N5), .Q(troj0_0_counter_2_) );
	edfxtp_1 troj0_0_Trojan_out0_0_reg( .D(troj0_0_N7), .DE(troj0_0_N5), .CLK(CLK), .Q(Trojan_out_0_0) );
	mux2_1 troj0_0_U3( .A0(troj0_0_counter_2_), .A1(troj0_0_N4), .S(Trigger_en_0_0), .X(troj0_0_n1) );
	mux2_1 troj0_0_U4( .A0(troj0_0_counter_1_), .A1(troj0_0_N3), .S(Trigger_en_0_0), .X(troj0_0_n2) );
	xor2_1 troj0_0_U5( .A(troj0_0_counter_0_), .B(Trigger_en_0_0), .X(troj0_0_n3) );
	nor3_2 troj0_0_U6( .A(n4571), .B(n11169), .C(troj0_0_n5), .Y(Trigger_en_0_0) );
	xnor2_1 troj0_0_U7( .A(troj0_0_n4), .B(tempn5237), .Y(n5237) );
	nand2_1 troj0_0_U8( .A(Trojan_out_0_0), .B(Trigger_en_0_0), .Y(troj0_0_n4) );
	or3_1 troj0_0_U9( .A(n8387), .B(n6429), .C(n5354), .X(troj0_0_n5) );
	and3_1 troj0_0_U10( .A(troj0_0_counter_2_), .B(troj0_0_counter_0_), .C(troj0_0_counter_1_), .X(troj0_0_N7) );
	inv_1 troj0_0_U11( .A(RST), .Y(troj0_0_N5) );
	xnor2_1 troj0_0_U12( .A(troj0_0_counter_2_), .B(troj0_0_n6), .Y(troj0_0_N4) );
	nand2_1 troj0_0_U13( .A(troj0_0_counter_1_), .B(troj0_0_counter_0_), .Y(troj0_0_n6) );
	xnor2_1 troj0_0_U14( .A(troj0_0_counter_1_), .B(troj0_0_N2), .Y(troj0_0_N3) );
	inv_1 troj0_0_U15( .A(troj0_0_counter_0_), .Y(troj0_0_N2) );
endmodule
