module c3540 ( N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, 
    N116, N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, 
    N200, N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, 
    N274, N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, 
    N350, N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, 
    N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, 
    N5360, N5361 );
input  N1, N13, N20, N33, N41, N45, N50, N58, N68, N77, N87, N97, N107, N116, 
    N124, N125, N128, N132, N137, N143, N150, N159, N169, N179, N190, N200, 
    N213, N222, N223, N226, N232, N238, N244, N250, N257, N264, N270, N274, 
    N283, N294, N303, N311, N317, N322, N326, N329, N330, N343, N349, N350;
output N1713, N1947, N3195, N3833, N3987, N4028, N4145, N4589, N4667, N4815, 
    N4944, N5002, N5045, N5047, N5078, N5102, N5120, N5121, N5192, N5231, 
    N5360, N5361;
    wire n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
        n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
        n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
        n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
        n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
        n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
        n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
        n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
        n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
        n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
        n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
        n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
        n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
        n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
        n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, 
        n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, 
        n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, 
        n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
        n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, 
        n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
        n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
        n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
        n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, 
        n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, 
        n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, 
        n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, 
        n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
        n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
        n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
        n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, 
        n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, 
        n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
        n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, 
        n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, 
        n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, 
        n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
        n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
        n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
        n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
        n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
        n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
        n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
        n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
        n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
        n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
        n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
        n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
        n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
        n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
        n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
        n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
        n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
        n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
        n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
        n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
        n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
        n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
        n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
        n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
        n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
        n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
        n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
        n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
        n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
        n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
        n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
        n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
        n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
        n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
        n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
        n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
        n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
        n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
        n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
        n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
        n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
        n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
        n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
        n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
        n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
        n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
        n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
        n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
        n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
        n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
        n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
        n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
        n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
        n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
        n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
        n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
        n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
        n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
        n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
        n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
        n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
        n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
        n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669;

wire Trigger_en51_0,  troj51_0n1,  troj51_0n2,  troj51_0n3,  troj51_0n4,  tempn1000;

    nnd2s1 U1 ( .Q(N5121), .DIN1(n558), .DIN2(n559) );
    nnd2s1 U2 ( .Q(N5120), .DIN1(n560), .DIN2(n561) );
    nnd2s1 U3 ( .Q(N5102), .DIN1(n562), .DIN2(n563) );
    nnd2s1 U4 ( .Q(N5078), .DIN1(n564), .DIN2(n565) );
    nnd2s1 U5 ( .Q(N5047), .DIN1(n566), .DIN2(n567) );
    nnd2s1 U6 ( .Q(N4944), .DIN1(n568), .DIN2(n569) );
    nor2s1 U7 ( .Q(n570), .DIN1(n571), .DIN2(n572) );
    nor2s1 U8 ( .Q(n573), .DIN1(n571), .DIN2(n574) );
    nor2s1 U9 ( .Q(n575), .DIN1(n576), .DIN2(n577) );
    nor2s1 U10 ( .Q(n578), .DIN1(n579), .DIN2(n580) );
    nor2s1 U11 ( .Q(n581), .DIN1(n582), .DIN2(n583) );
    nnd2s1 U12 ( .Q(N5231), .DIN1(n584), .DIN2(N213) );
    nnd2s1 U13 ( .Q(N5192), .DIN1(n585), .DIN2(n586) );
    nnd2s1 U14 ( .Q(N5045), .DIN1(n587), .DIN2(n588) );
    nnd2s1 U15 ( .Q(N5002), .DIN1(n589), .DIN2(n590) );
    nnd2s1 U16 ( .Q(N4815), .DIN1(n591), .DIN2(n592) );
    nnd2s1 U17 ( .Q(N4667), .DIN1(n593), .DIN2(n594) );
    nnd2s1 U18 ( .Q(N4589), .DIN1(n595), .DIN2(n596) );
    nnd2s1 U19 ( .Q(N4145), .DIN1(n597), .DIN2(n598) );
    nor2s1 U20 ( .Q(N4028), .DIN1(n599), .DIN2(n600) );
    nor2s1 U21 ( .Q(N3195), .DIN1(n601), .DIN2(n602) );
    nnd2s1 U22 ( .Q(N1947), .DIN1(N87), .DIN2(n603) );
    nor2s1 U23 ( .Q(N1713), .DIN1(n604), .DIN2(n605) );
    nor2s1 U24 ( .Q(n606), .DIN1(N50), .DIN2(n607) );
    nor2s1 U25 ( .Q(n608), .DIN1(n606), .DIN2(n609) );
    nor2s1 U26 ( .Q(n610), .DIN1(N58), .DIN2(n608) );
    nor2s1 U27 ( .Q(n611), .DIN1(N349), .DIN2(N33) );
    nor2s1 U28 ( .Q(n612), .DIN1(n613), .DIN2(n614) );
    nor2s1 U29 ( .Q(n615), .DIN1(n616), .DIN2(n617) );
    nor2s1 U30 ( .Q(n618), .DIN1(n619), .DIN2(n620) );
    nor2s1 U31 ( .Q(n621), .DIN1(N50), .DIN2(n622) );
    nor2s1 U32 ( .Q(n623), .DIN1(n624), .DIN2(n625) );
    nor2s1 U33 ( .Q(n626), .DIN1(n627), .DIN2(n628) );
    nor2s1 U34 ( .Q(n629), .DIN1(n613), .DIN2(n619) );
    nor2s1 U35 ( .Q(n630), .DIN1(n616), .DIN2(n631) );
    nor2s1 U36 ( .Q(n632), .DIN1(n620), .DIN2(n633) );
    nor2s1 U37 ( .Q(n634), .DIN1(N159), .DIN2(n635) );
    nor2s1 U38 ( .Q(n636), .DIN1(n637), .DIN2(n638) );
    nor2s1 U39 ( .Q(n639), .DIN1(N77), .DIN2(n640) );
    nor2s1 U40 ( .Q(n641), .DIN1(N50), .DIN2(n635) );
    nor2s1 U41 ( .Q(n642), .DIN1(n643), .DIN2(n644) );
    nor2s1 U42 ( .Q(n645), .DIN1(n613), .DIN2(n633) );
    nor2s1 U43 ( .Q(n646), .DIN1(n616), .DIN2(n647) );
    nor2s1 U44 ( .Q(n648), .DIN1(n649), .DIN2(n620) );
    nor2s1 U45 ( .Q(n650), .DIN1(N87), .DIN2(n640) );
    nor2s1 U46 ( .Q(n651), .DIN1(N58), .DIN2(n635) );
    nor2s1 U47 ( .Q(n652), .DIN1(N77), .DIN2(n643) );
    nor2s1 U48 ( .Q(n653), .DIN1(n649), .DIN2(n613) );
    nor2s1 U49 ( .Q(n654), .DIN1(n616), .DIN2(n655) );
    nor2s1 U50 ( .Q(n656), .DIN1(n620), .DIN2(n657) );
    nor2s1 U51 ( .Q(n658), .DIN1(N87), .DIN2(n659) );
    nor2s1 U52 ( .Q(n660), .DIN1(n658), .DIN2(n609) );
    nor2s1 U53 ( .Q(n661), .DIN1(N97), .DIN2(n660) );
    nor2s1 U54 ( .Q(n662), .DIN1(n613), .DIN2(n657) );
    nor2s1 U55 ( .Q(n663), .DIN1(n616), .DIN2(n664) );
    nor2s1 U56 ( .Q(n665), .DIN1(n620), .DIN2(n666) );
    nor2s1 U57 ( .Q(n667), .DIN1(n613), .DIN2(n666) );
    nor2s1 U58 ( .Q(n668), .DIN1(n616), .DIN2(n669) );
    nor2s1 U59 ( .Q(n670), .DIN1(n620), .DIN2(n671) );
    nor2s1 U60 ( .Q(n672), .DIN1(N77), .DIN2(n635) );
    nor2s1 U61 ( .Q(n673), .DIN1(n674), .DIN2(n675) );
    nor2s1 U62 ( .Q(n676), .DIN1(N283), .DIN2(n640) );
    nor2s1 U63 ( .Q(n677), .DIN1(N97), .DIN2(n635) );
    nor2s1 U64 ( .Q(n678), .DIN1(N116), .DIN2(n643) );
    nor2s1 U65 ( .Q(n679), .DIN1(n613), .DIN2(n680) );
    nor2s1 U66 ( .Q(n681), .DIN1(n616), .DIN2(n682) );
    nor2s1 U67 ( .Q(n683), .DIN1(n620), .DIN2(n684) );
    nor2s1 U68 ( .Q(n685), .DIN1(N116), .DIN2(n640) );
    nor2s1 U69 ( .Q(n686), .DIN1(N87), .DIN2(n635) );
    nor2s1 U70 ( .Q(n687), .DIN1(n643), .DIN2(n655) );
    nor2s1 U71 ( .Q(n688), .DIN1(n613), .DIN2(n671) );
    nor2s1 U72 ( .Q(n689), .DIN1(n616), .DIN2(n690) );
    nor2s1 U73 ( .Q(n691), .DIN1(n620), .DIN2(n680) );
    nor2s1 U74 ( .Q(n692), .DIN1(n571), .DIN2(n693) );
    nnd2s1 U75 ( .Q(n694), .DIN1(n695), .DIN2(n696) );
    nor2s1 U76 ( .Q(n697), .DIN1(n698), .DIN2(n699) );
    nor2s1 U77 ( .Q(n700), .DIN1(n697), .DIN2(n701) );
    nor2s1 U78 ( .Q(n702), .DIN1(n700), .DIN2(n703) );
    nor2s1 U79 ( .Q(n704), .DIN1(n705), .DIN2(n706) );
    nor2s1 U80 ( .Q(n707), .DIN1(n708), .DIN2(n709) );
    nor2s1 U81 ( .Q(n710), .DIN1(n647), .DIN2(n711) );
    nor2s1 U82 ( .Q(n712), .DIN1(n655), .DIN2(n713) );
    nor2s1 U83 ( .Q(n714), .DIN1(n664), .DIN2(n715) );
    nor2s1 U84 ( .Q(n716), .DIN1(n669), .DIN2(n717) );
    nor2s1 U85 ( .Q(n718), .DIN1(n719), .DIN2(n720) );
    nor2s1 U86 ( .Q(n721), .DIN1(n722), .DIN2(n723) );
    nor2s1 U87 ( .Q(n724), .DIN1(n711), .DIN2(n725) );
    nnd2s1 U88 ( .Q(n726), .DIN1(n727), .DIN2(N137) );
    nor2s1 U89 ( .Q(n728), .DIN1(n715), .DIN2(n729) );
    nor2s1 U90 ( .Q(n730), .DIN1(n717), .DIN2(n731) );
    nor2s1 U91 ( .Q(n732), .DIN1(n733), .DIN2(n734) );
    nor2s1 U92 ( .Q(n735), .DIN1(n736), .DIN2(n737) );
    nor2s1 U93 ( .Q(n738), .DIN1(n739), .DIN2(n740) );
    nor2s1 U94 ( .Q(n741), .DIN1(n682), .DIN2(n742) );
    nor2s1 U95 ( .Q(n743), .DIN1(n647), .DIN2(n722) );
    nor2s1 U96 ( .Q(n744), .DIN1(n742), .DIN2(n731) );
    nor2s1 U97 ( .Q(n745), .DIN1(N68), .DIN2(n622) );
    nor2s1 U98 ( .Q(n746), .DIN1(n695), .DIN2(n628) );
    nor2s1 U99 ( .Q(n747), .DIN1(n748), .DIN2(n708) );
    nor2s1 U100 ( .Q(n749), .DIN1(n747), .DIN2(n750) );
    nor2s1 U101 ( .Q(n751), .DIN1(n742), .DIN2(n752) );
    nor2s1 U102 ( .Q(n753), .DIN1(n655), .DIN2(n722) );
    nor2s1 U103 ( .Q(n754), .DIN1(n742), .DIN2(n729) );
    nor2s1 U104 ( .Q(n755), .DIN1(N77), .DIN2(n622) );
    nor2s1 U105 ( .Q(n756), .DIN1(n628), .DIN2(n757) );
    nor2s1 U106 ( .Q(n758), .DIN1(n759), .DIN2(n596) );
    nor2s1 U107 ( .Q(n760), .DIN1(n761), .DIN2(n708) );
    nor2s1 U108 ( .Q(n762), .DIN1(n669), .DIN2(n722) );
    nor2s1 U109 ( .Q(n763), .DIN1(n690), .DIN2(n711) );
    nor2s1 U110 ( .Q(n764), .DIN1(n682), .DIN2(n713) );
    nor2s1 U111 ( .Q(n765), .DIN1(n715), .DIN2(n752) );
    nor2s1 U112 ( .Q(n766), .DIN1(n717), .DIN2(n767) );
    nor2s1 U113 ( .Q(n768), .DIN1(n742), .DIN2(n725) );
    nor2s1 U114 ( .Q(n769), .DIN1(n644), .DIN2(n722) );
    nor2s1 U115 ( .Q(n770), .DIN1(n771), .DIN2(n711) );
    nor2s1 U116 ( .Q(n772), .DIN1(n773), .DIN2(n713) );
    nor2s1 U117 ( .Q(n774), .DIN1(n715), .DIN2(n720) );
    nor2s1 U118 ( .Q(n775), .DIN1(n717), .DIN2(n723) );
    nor2s1 U119 ( .Q(n776), .DIN1(n777), .DIN2(n778) );
    nor2s1 U120 ( .Q(n779), .DIN1(n780), .DIN2(n781) );
    nor2s1 U121 ( .Q(n782), .DIN1(n783), .DIN2(n784) );
    nor2s1 U122 ( .Q(n785), .DIN1(n742), .DIN2(n767) );
    nor2s1 U123 ( .Q(n786), .DIN1(n655), .DIN2(n719) );
    nor2s1 U124 ( .Q(n787), .DIN1(n788), .DIN2(n789) );
    nor2s1 U125 ( .Q(n790), .DIN1(n787), .DIN2(n791) );
    nor2s1 U126 ( .Q(n792), .DIN1(n793), .DIN2(n794) );
    nor2s1 U127 ( .Q(n795), .DIN1(n759), .DIN2(n796) );
    nor2s1 U128 ( .Q(n797), .DIN1(n798), .DIN2(n675) );
    nor2s1 U129 ( .Q(n799), .DIN1(n800), .DIN2(n801) );
    nnd2s1 U130 ( .Q(n802), .DIN1(n803), .DIN2(N326) );
    nor2s1 U131 ( .Q(n804), .DIN1(n664), .DIN2(n805) );
    nor2s1 U132 ( .Q(n806), .DIN1(n799), .DIN2(n791) );
    nor2s1 U133 ( .Q(n807), .DIN1(n808), .DIN2(n793) );
    nor2s1 U134 ( .Q(n809), .DIN1(n810), .DIN2(n708) );
    nor2s1 U135 ( .Q(n811), .DIN1(n809), .DIN2(n750) );
    nor2s1 U136 ( .Q(n812), .DIN1(N77), .DIN2(N68) );
    nor2s1 U137 ( .Q(n813), .DIN1(n814), .DIN2(n815) );
    nnd2s1 U138 ( .Q(n816), .DIN1(n803), .DIN2(N329) );
    nor2s1 U139 ( .Q(n817), .DIN1(n669), .DIN2(n805) );
    nor2s1 U140 ( .Q(n818), .DIN1(n813), .DIN2(n791) );
    nor2s1 U141 ( .Q(n819), .DIN1(n793), .DIN2(n820) );
    nor2s1 U142 ( .Q(n821), .DIN1(N330), .DIN2(n820) );
    nor2s1 U143 ( .Q(n822), .DIN1(N343), .DIN2(n823) );
    nor2s1 U144 ( .Q(n824), .DIN1(n825), .DIN2(n826) );
    nor2s1 U145 ( .Q(n827), .DIN1(N264), .DIN2(N257) );
    nor2s1 U146 ( .Q(n828), .DIN1(n633), .DIN2(n773) );
    nor2s1 U147 ( .Q(n829), .DIN1(n771), .DIN2(n649) );
    nor2s1 U148 ( .Q(n830), .DIN1(n644), .DIN2(n657) );
    nor2s1 U149 ( .Q(n831), .DIN1(n617), .DIN2(n666) );
    nor2s1 U150 ( .Q(n832), .DIN1(n631), .DIN2(n671) );
    nor2s1 U151 ( .Q(n833), .DIN1(n647), .DIN2(n680) );
    nor2s1 U152 ( .Q(n834), .DIN1(n655), .DIN2(n684) );
    nor2s1 U153 ( .Q(n835), .DIN1(n664), .DIN2(n836) );
    nor2s1 U154 ( .Q(n837), .DIN1(n838), .DIN2(n839) );
    nor2s1 U155 ( .Q(n840), .DIN1(n841), .DIN2(n842) );
    nor2s1 U156 ( .Q(n843), .DIN1(n607), .DIN2(n771) );
    nor2s1 U157 ( .Q(n844), .DIN1(n647), .DIN2(n659) );
    nor2s1 U158 ( .Q(n800), .DIN1(n845), .DIN2(n846) );
    nor2s1 U159 ( .Q(n814), .DIN1(n847), .DIN2(n846) );
    nor2s1 U160 ( .Q(n825), .DIN1(N58), .DIN2(n848) );
    nor2s1 U161 ( .Q(n601), .DIN1(n849), .DIN2(n850) );
    hi1s1 U162 ( .Q(n851), .DIN(N45) );
    hi1s1 U163 ( .Q(n852), .DIN(N13) );
    hi1s1 U164 ( .Q(n853), .DIN(N1) );
    hi1s1 U165 ( .Q(n643), .DIN(N20) );
    nor2s1 U166 ( .Q(n854), .DIN1(n643), .DIN2(n853) );
    nnd2s1 U167 ( .Q(n855), .DIN1(n854), .DIN2(n852) );
    hi1s1 U168 ( .Q(n856), .DIN(N33) );
    nor2s1 U169 ( .Q(n857), .DIN1(n609), .DIN2(N20) );
    nor2s1 U170 ( .Q(n609), .DIN1(n856), .DIN2(N20) );
    hi1s1 U171 ( .Q(n644), .DIN(N68) );
    nnd2s1 U172 ( .Q(n607), .DIN1(N20), .DIN2(n644) );
    hi1s1 U173 ( .Q(n771), .DIN(N58) );
    nnd2s1 U174 ( .Q(n858), .DIN1(N20), .DIN2(n853) );
    nnd2s1 U175 ( .Q(n859), .DIN1(n860), .DIN2(n861) );
    nor2s1 U176 ( .Q(n862), .DIN1(n859), .DIN2(n863) );
    nor2s1 U177 ( .Q(n864), .DIN1(N1), .DIN2(n865) );
    hi1s1 U178 ( .Q(n866), .DIN(N41) );
    nnd2s1 U179 ( .Q(n860), .DIN1(N1), .DIN2(N13) );
    nor2s1 U180 ( .Q(n867), .DIN1(n864), .DIN2(n868) );
    hi1s1 U181 ( .Q(n649), .DIN(N232) );
    nor2s1 U182 ( .Q(n868), .DIN1(n860), .DIN2(n869) );
    nnd2s1 U183 ( .Q(n613), .DIN1(n868), .DIN2(n611) );
    hi1s1 U184 ( .Q(n619), .DIN(N223) );
    nnd2s1 U185 ( .Q(n616), .DIN1(n868), .DIN2(N33) );
    hi1s1 U186 ( .Q(n631), .DIN(N87) );
    nnd2s1 U187 ( .Q(n620), .DIN1(n870), .DIN2(n868) );
    hi1s1 U188 ( .Q(n633), .DIN(N226) );
    hi1s1 U189 ( .Q(n871), .DIN(N190) );
    hi1s1 U190 ( .Q(n872), .DIN(N200) );
    nnd2s1 U191 ( .Q(n873), .DIN1(n874), .DIN2(n875) );
    hi1s1 U192 ( .Q(n657), .DIN(N238) );
    hi1s1 U193 ( .Q(n647), .DIN(N97) );
    hi1s1 U194 ( .Q(n876), .DIN(N179) );
    nnd2s1 U195 ( .Q(n698), .DIN1(n638), .DIN2(n877) );
    hi1s1 U196 ( .Q(n773), .DIN(N50) );
    hi1s1 U197 ( .Q(n614), .DIN(N222) );
    hi1s1 U198 ( .Q(n617), .DIN(N77) );
    hi1s1 U199 ( .Q(n666), .DIN(N244) );
    hi1s1 U200 ( .Q(n655), .DIN(N107) );
    nnd2s1 U201 ( .Q(n705), .DIN1(n878), .DIN2(n879) );
    nnd2s1 U202 ( .Q(n706), .DIN1(n880), .DIN2(n881) );
    nnd2s1 U203 ( .Q(n881), .DIN1(n882), .DIN2(n883) );
    nnd2s1 U204 ( .Q(n884), .DIN1(n706), .DIN2(n885) );
    hi1s1 U205 ( .Q(n886), .DIN(N213) );
    nnd2s1 U206 ( .Q(n887), .DIN1(n888), .DIN2(n889) );
    hi1s1 U207 ( .Q(n664), .DIN(N116) );
    nor2s1 U208 ( .Q(n890), .DIN1(n851), .DIN2(N1) );
    nor2s1 U209 ( .Q(n891), .DIN1(n892), .DIN2(N41) );
    nor2s1 U210 ( .Q(n893), .DIN1(n868), .DIN2(n891) );
    hi1s1 U211 ( .Q(n836), .DIN(N270) );
    hi1s1 U212 ( .Q(n680), .DIN(N257) );
    hi1s1 U213 ( .Q(n682), .DIN(N303) );
    hi1s1 U214 ( .Q(n684), .DIN(N264) );
    nnd2s1 U215 ( .Q(n894), .DIN1(n895), .DIN2(n896) );
    nnd2s1 U216 ( .Q(n659), .DIN1(N20), .DIN2(n655) );
    hi1s1 U217 ( .Q(n671), .DIN(N250) );
    nnd2s1 U218 ( .Q(n897), .DIN1(n898), .DIN2(n899) );
    nnd2s1 U219 ( .Q(n900), .DIN1(n901), .DIN2(n902) );
    hi1s1 U220 ( .Q(n669), .DIN(N283) );
    nnd2s1 U221 ( .Q(n903), .DIN1(n904), .DIN2(n905) );
    nnd2s1 U222 ( .Q(n906), .DIN1(n907), .DIN2(n908) );
    hi1s1 U223 ( .Q(n690), .DIN(N294) );
    nnd2s1 U224 ( .Q(n909), .DIN1(n910), .DIN2(n911) );
    nnd2s1 U225 ( .Q(n912), .DIN1(n675), .DIN2(n913) );
    nnd2s1 U226 ( .Q(n674), .DIN1(n914), .DIN2(n915) );
    nnd2s1 U227 ( .Q(n579), .DIN1(n916), .DIN2(n917) );
    nnd2s1 U228 ( .Q(n580), .DIN1(n918), .DIN2(n919) );
    nnd2s1 U229 ( .Q(n675), .DIN1(n920), .DIN2(n906) );
    nnd2s1 U230 ( .Q(n921), .DIN1(n922), .DIN2(n923) );
    nor2s1 U231 ( .Q(n924), .DIN1(n884), .DIN2(n705) );
    nnd2s1 U232 ( .Q(n925), .DIN1(n926), .DIN2(n927) );
    nnd2s1 U233 ( .Q(n923), .DIN1(N343), .DIN2(n637) );
    nnd2s1 U234 ( .Q(n919), .DIN1(n928), .DIN2(n929) );
    nnd2s1 U235 ( .Q(n930), .DIN1(n580), .DIN2(n931) );
    nnd2s1 U236 ( .Q(n932), .DIN1(N330), .DIN2(n933) );
    nor2s1 U237 ( .Q(n934), .DIN1(n925), .DIN2(n935) );
    nor2s1 U238 ( .Q(n696), .DIN1(n932), .DIN2(n936) );
    nnd2s1 U239 ( .Q(n937), .DIN1(n934), .DIN2(n938) );
    nor2s1 U240 ( .Q(n939), .DIN1(n855), .DIN2(N41) );
    nnd2s1 U241 ( .Q(n750), .DIN1(N1), .DIN2(n940) );
    nnd2s1 U242 ( .Q(n572), .DIN1(n941), .DIN2(n695) );
    nnd2s1 U243 ( .Q(n574), .DIN1(n942), .DIN2(n695) );
    nnd2s1 U244 ( .Q(n638), .DIN1(n943), .DIN2(n873) );
    nnd2s1 U245 ( .Q(n693), .DIN1(n944), .DIN2(n945) );
    nor2s1 U246 ( .Q(n946), .DIN1(n947), .DIN2(n948) );
    nnd2s1 U247 ( .Q(n949), .DIN1(n950), .DIN2(n951) );
    nnd2s1 U248 ( .Q(n622), .DIN1(n628), .DIN2(n624) );
    nnd2s1 U249 ( .Q(n742), .DIN1(n952), .DIN2(n953) );
    nor2s1 U250 ( .Q(n954), .DIN1(n872), .DIN2(n643) );
    nnd2s1 U251 ( .Q(n805), .DIN1(n955), .DIN2(n954) );
    nor2s1 U252 ( .Q(n956), .DIN1(n957), .DIN2(n876) );
    nnd2s1 U253 ( .Q(n711), .DIN1(n956), .DIN2(n871) );
    nnd2s1 U254 ( .Q(n713), .DIN1(n958), .DIN2(n954) );
    nnd2s1 U255 ( .Q(n715), .DIN1(n956), .DIN2(N190) );
    nnd2s1 U256 ( .Q(n717), .DIN1(n959), .DIN2(n954) );
    nor2s1 U257 ( .Q(n960), .DIN1(n871), .DIN2(N179) );
    nnd2s1 U258 ( .Q(n722), .DIN1(n960), .DIN2(n954) );
    nor2s1 U259 ( .Q(n961), .DIN1(n954), .DIN2(n962) );
    hi1s1 U260 ( .Q(n720), .DIN(N159) );
    hi1s1 U261 ( .Q(n723), .DIN(N150) );
    hi1s1 U262 ( .Q(n725), .DIN(N143) );
    hi1s1 U263 ( .Q(n729), .DIN(N132) );
    hi1s1 U264 ( .Q(n731), .DIN(N128) );
    nor2s1 U265 ( .Q(n963), .DIN1(n860), .DIN2(n964) );
    nor2s1 U266 ( .Q(n788), .DIN1(N13), .DIN2(N33) );
    nor2s1 U267 ( .Q(n965), .DIN1(n750), .DIN2(n939) );
    nor2s1 U268 ( .Q(n966), .DIN1(n624), .DIN2(N33) );
    nor2s1 U269 ( .Q(n967), .DIN1(n624), .DIN2(n856) );
    nor2s1 U270 ( .Q(n968), .DIN1(n580), .DIN2(n798) );
    nnd2s1 U271 ( .Q(n969), .DIN1(N330), .DIN2(n820) );
    nnd2s1 U272 ( .Q(n970), .DIN1(n921), .DIN2(n932) );
    nnd2s1 U273 ( .Q(n596), .DIN1(n808), .DIN2(n971) );
    nnd2s1 U274 ( .Q(n972), .DIN1(n796), .DIN2(n973) );
    hi1s1 U275 ( .Q(n752), .DIN(N311) );
    hi1s1 U276 ( .Q(n767), .DIN(N317) );
    nor2s1 U277 ( .Q(n974), .DIN1(n856), .DIN2(n855) );
    nor2s1 U278 ( .Q(n975), .DIN1(n963), .DIN2(n976) );
    nor2s1 U279 ( .Q(n976), .DIN1(n628), .DIN2(N20) );
    nnd2s1 U280 ( .Q(n796), .DIN1(n977), .DIN2(n978) );
    nnd2s1 U281 ( .Q(n979), .DIN1(n980), .DIN2(n981) );
    nor2s1 U282 ( .Q(n982), .DIN1(n617), .DIN2(n644) );
    nnd2s1 U283 ( .Q(n849), .DIN1(n854), .DIN2(N13) );
    nnd2s1 U284 ( .Q(n850), .DIN1(N50), .DIN2(n604) );
    nnd2s1 U285 ( .Q(n983), .DIN1(n984), .DIN2(n985) );
    nnd2s1 U286 ( .Q(n986), .DIN1(n987), .DIN2(n988) );
    nnd2s1 U287 ( .Q(n604), .DIN1(n771), .DIN2(n644) );
    nor2s1 U288 ( .Q(n695), .DIN1(n989), .DIN2(n990) );
    nor2s1 U289 ( .Q(n936), .DIN1(n991), .DIN2(n992) );
    nor2s1 U290 ( .Q(n993), .DIN1(n994), .DIN2(n995) );
    nor2s1 U291 ( .Q(n571), .DIN1(n996), .DIN2(n997) );
    nor2s1 U292 ( .Q(n998), .DIN1(n999), .DIN2(n1000) );
    nor2s1 U293 ( .Q(n627), .DIN1(n1001), .DIN2(n1002) );
    nnd2s1 U294 ( .Q(n709), .DIN1(n1003), .DIN2(n1004) );
    nnd2s1 U295 ( .Q(n1005), .DIN1(n1006), .DIN2(n1007) );
    nnd2s1 U296 ( .Q(n820), .DIN1(n1008), .DIN2(n1009) );
    nnd2s1 U297 ( .Q(n576), .DIN1(n1010), .DIN2(n1011) );
    nor2s1 U298 ( .Q(n1012), .DIN1(n1013), .DIN2(n1014) );
    nnd2s1 U299 ( .Q(n794), .DIN1(n1015), .DIN2(n1016) );
    nor2s1 U300 ( .Q(n1017), .DIN1(n1018), .DIN2(n1019) );
    nor2s1 U301 ( .Q(n1020), .DIN1(n1021), .DIN2(n1022) );
    nnd2s1 U302 ( .Q(n1023), .DIN1(n1024), .DIN2(n1025) );
    nnd2s1 U303 ( .Q(N5360), .DIN1(n1026), .DIN2(n1027) );
    nnd2s1 U304 ( .Q(N3987), .DIN1(n1028), .DIN2(n1029) );
    nnd2s1 U305 ( .Q(N3833), .DIN1(n1030), .DIN2(n1031) );
    nnd2s1 U306 ( .Q(n1032), .DIN1(n1033), .DIN2(n582) );
    nor2s1 U307 ( .Q(n1034), .DIN1(N97), .DIN2(n643) );
    nnd2s1 U308 ( .Q(n1035), .DIN1(n1036), .DIN2(n1037) );
    nor2s1 U309 ( .Q(n1038), .DIN1(n868), .DIN2(n671) );
    nnd2s1 U310 ( .Q(n1039), .DIN1(n1040), .DIN2(n1041) );
    nor2s1 U311 ( .Q(n1042), .DIN1(n1043), .DIN2(n1044) );
    nor2s1 U312 ( .Q(n1045), .DIN1(n1046), .DIN2(n1047) );
    nnd2s1 U313 ( .Q(n1048), .DIN1(n1049), .DIN2(n699) );
    nor2s1 U314 ( .Q(n1050), .DIN1(N58), .DIN2(n643) );
    nnd2s1 U315 ( .Q(n1051), .DIN1(n1052), .DIN2(n1053) );
    nnd2s1 U316 ( .Q(n703), .DIN1(n1054), .DIN2(n927) );
    nnd2s1 U317 ( .Q(n625), .DIN1(n1055), .DIN2(n1056) );
    nnd2s1 U318 ( .Q(n1057), .DIN1(n1058), .DIN2(n1059) );
    nnd2s1 U319 ( .Q(n789), .DIN1(n1060), .DIN2(n1061) );
    nnd2s1 U320 ( .Q(n845), .DIN1(n1062), .DIN2(n1063) );
    nor2s1 U321 ( .Q(n1064), .DIN1(N107), .DIN2(n974) );
    nnd2s1 U322 ( .Q(n801), .DIN1(n1065), .DIN2(n1066) );
    nnd2s1 U323 ( .Q(n847), .DIN1(n1067), .DIN2(n1068) );
    nor2s1 U324 ( .Q(n1069), .DIN1(N116), .DIN2(n974) );
    nnd2s1 U325 ( .Q(n815), .DIN1(n1070), .DIN2(n1071) );
    nor2s1 U326 ( .Q(n1072), .DIN1(n617), .DIN2(n1073) );
    nnd2s1 U327 ( .Q(n826), .DIN1(n1074), .DIN2(n1075) );
    nor2s1 U328 ( .Q(n1076), .DIN1(n827), .DIN2(n671) );
    nor2s1 U329 ( .Q(n1077), .DIN1(n1078), .DIN2(n837) );
    nnd2s1 U330 ( .Q(n602), .DIN1(n1079), .DIN2(n1080) );
    nnd2s1 U331 ( .Q(n1081), .DIN1(n1082), .DIN2(n1083) );
    nor2s1 U332 ( .Q(n1084), .DIN1(n1085), .DIN2(n650) );
    nor2s1 U333 ( .Q(n1086), .DIN1(n651), .DIN2(n652) );
    nor2s1 U334 ( .Q(n870), .DIN1(N33), .DIN2(n611) );
    nnd2s1 U335 ( .Q(n1087), .DIN1(n1088), .DIN2(n1089) );
    nor2s1 U336 ( .Q(n1090), .DIN1(n653), .DIN2(n1087) );
    nor2s1 U337 ( .Q(n1091), .DIN1(n654), .DIN2(n656) );
    nor2s1 U338 ( .Q(n889), .DIN1(N1), .DIN2(N20) );
    nor2s1 U339 ( .Q(n888), .DIN1(n852), .DIN2(n886) );
    nnd2s1 U340 ( .Q(n1092), .DIN1(n1093), .DIN2(n1094) );
    nor2s1 U341 ( .Q(n911), .DIN1(n688), .DIN2(n1092) );
    nor2s1 U342 ( .Q(n910), .DIN1(n689), .DIN2(n691) );
    nor2s1 U343 ( .Q(n1095), .DIN1(n1085), .DIN2(n685) );
    nor2s1 U344 ( .Q(n1096), .DIN1(n686), .DIN2(n687) );
    nor2s1 U345 ( .Q(n1097), .DIN1(n1085), .DIN2(n672) );
    nor2s1 U346 ( .Q(n1098), .DIN1(n844), .DIN2(n1035) );
    nnd2s1 U347 ( .Q(n1099), .DIN1(n1100), .DIN2(n1094) );
    nor2s1 U348 ( .Q(n905), .DIN1(n667), .DIN2(n1099) );
    nor2s1 U349 ( .Q(n904), .DIN1(n668), .DIN2(n670) );
    nor2s1 U350 ( .Q(n1101), .DIN1(n1085), .DIN2(n661) );
    nor2s1 U351 ( .Q(n899), .DIN1(n662), .DIN2(n663) );
    nor2s1 U352 ( .Q(n898), .DIN1(n665), .DIN2(n1039) );
    nor2s1 U353 ( .Q(n916), .DIN1(n912), .DIN2(n1032) );
    nor2s1 U354 ( .Q(n1102), .DIN1(n1085), .DIN2(n676) );
    nor2s1 U355 ( .Q(n1103), .DIN1(n677), .DIN2(n678) );
    nnd2s1 U356 ( .Q(n1104), .DIN1(n1105), .DIN2(n1094) );
    nor2s1 U357 ( .Q(n896), .DIN1(n679), .DIN2(n1104) );
    nor2s1 U358 ( .Q(n895), .DIN1(n681), .DIN2(n683) );
    nnd2s1 U359 ( .Q(n582), .DIN1(n978), .DIN2(n1106) );
    nnd2s1 U360 ( .Q(n583), .DIN1(n917), .DIN2(n1107) );
    nor2s1 U361 ( .Q(n1108), .DIN1(n578), .DIN2(n581) );
    nor2s1 U362 ( .Q(n1109), .DIN1(n1110), .DIN2(n673) );
    nnd2s1 U363 ( .Q(n1046), .DIN1(n903), .DIN2(n897) );
    nnd2s1 U364 ( .Q(n1047), .DIN1(n909), .DIN2(n894) );
    nnd2s1 U365 ( .Q(n1043), .DIN1(n1111), .DIN2(n1112) );
    nnd2s1 U366 ( .Q(n1044), .DIN1(n1113), .DIN2(n1114) );
    nor2s1 U367 ( .Q(n1115), .DIN1(n941), .DIN2(n942) );
    nor2s1 U368 ( .Q(n1116), .DIN1(n1085), .DIN2(n639) );
    nor2s1 U369 ( .Q(n1117), .DIN1(n641), .DIN2(n642) );
    nnd2s1 U370 ( .Q(n1118), .DIN1(n1119), .DIN2(n1089) );
    nor2s1 U371 ( .Q(n1120), .DIN1(n645), .DIN2(n1118) );
    nor2s1 U372 ( .Q(n1121), .DIN1(n646), .DIN2(n648) );
    nor2s1 U373 ( .Q(n941), .DIN1(n936), .DIN2(n921) );
    nor2s1 U374 ( .Q(n942), .DIN1(n798), .DIN2(n706) );
    nor2s1 U375 ( .Q(n944), .DIN1(n798), .DIN2(n1122) );
    nnd2s1 U376 ( .Q(n1123), .DIN1(n572), .DIN2(n574) );
    nnd2s1 U377 ( .Q(n1124), .DIN1(n693), .DIN2(n694) );
    nor2s1 U378 ( .Q(n1125), .DIN1(n1085), .DIN2(n634) );
    nor2s1 U379 ( .Q(n1126), .DIN1(n843), .DIN2(n1051) );
    nnd2s1 U380 ( .Q(n1127), .DIN1(n1128), .DIN2(n1089) );
    nor2s1 U381 ( .Q(n1129), .DIN1(n629), .DIN2(n1127) );
    nor2s1 U382 ( .Q(n1130), .DIN1(n630), .DIN2(n632) );
    nnd2s1 U383 ( .Q(n1131), .DIN1(n1132), .DIN2(n1089) );
    nor2s1 U384 ( .Q(n1133), .DIN1(n612), .DIN2(n1131) );
    nor2s1 U385 ( .Q(n1134), .DIN1(n615), .DIN2(n618) );
    nor2s1 U386 ( .Q(n1135), .DIN1(n1085), .DIN2(n610) );
    nor2s1 U387 ( .Q(n878), .DIN1(n698), .DIN2(n703) );
    nnd2s1 U388 ( .Q(n699), .DIN1(n945), .DIN2(n1136) );
    nor2s1 U389 ( .Q(n926), .DIN1(n702), .DIN2(n704) );
    nor2s1 U390 ( .Q(n1137), .DIN1(N20), .DIN2(n851) );
    nnd2s1 U391 ( .Q(n948), .DIN1(n933), .DIN2(n1138) );
    nnd2s1 U392 ( .Q(n947), .DIN1(n757), .DIN2(n695) );
    nor2s1 U393 ( .Q(n951), .DIN1(n570), .DIN2(n573) );
    nor2s1 U394 ( .Q(n950), .DIN1(n636), .DIN2(n692) );
    nor2s1 U395 ( .Q(n953), .DIN1(N190), .DIN2(N200) );
    nor2s1 U396 ( .Q(n952), .DIN1(N179), .DIN2(n643) );
    nor2s1 U397 ( .Q(n955), .DIN1(N190), .DIN2(N179) );
    nnd2s1 U398 ( .Q(n957), .DIN1(n872), .DIN2(N20) );
    nor2s1 U399 ( .Q(n958), .DIN1(N190), .DIN2(n876) );
    nor2s1 U400 ( .Q(n959), .DIN1(n871), .DIN2(n876) );
    nnd2s1 U401 ( .Q(n1139), .DIN1(n1140), .DIN2(n1141) );
    nnd2s1 U402 ( .Q(n1142), .DIN1(n1143), .DIN2(n1144) );
    nor2s1 U403 ( .Q(n1145), .DIN1(n1139), .DIN2(n1142) );
    nnd2s1 U404 ( .Q(n1146), .DIN1(n1147), .DIN2(n1148) );
    nnd2s1 U405 ( .Q(n1149), .DIN1(n1150), .DIN2(n1151) );
    nor2s1 U406 ( .Q(n1152), .DIN1(n1146), .DIN2(n1149) );
    nnd2s1 U407 ( .Q(n1153), .DIN1(n1154), .DIN2(n1155) );
    nnd2s1 U408 ( .Q(n1156), .DIN1(n1157), .DIN2(n1158) );
    nor2s1 U409 ( .Q(n1159), .DIN1(n1153), .DIN2(n1156) );
    nnd2s1 U410 ( .Q(n1160), .DIN1(n1161), .DIN2(n1162) );
    nor2s1 U411 ( .Q(n1163), .DIN1(n1164), .DIN2(n1165) );
    nor2s1 U412 ( .Q(n1166), .DIN1(n1160), .DIN2(n1167) );
    nor2s1 U413 ( .Q(n1168), .DIN1(n621), .DIN2(n623) );
    nor2s1 U414 ( .Q(n1169), .DIN1(n626), .DIN2(n1170) );
    nnd2s1 U415 ( .Q(n1171), .DIN1(n1172), .DIN2(n1173) );
    nor2s1 U416 ( .Q(n1174), .DIN1(n718), .DIN2(n1171) );
    nor2s1 U417 ( .Q(n1175), .DIN1(n721), .DIN2(n724) );
    nnd2s1 U418 ( .Q(n733), .DIN1(n1175), .DIN2(n1174) );
    nor2s1 U419 ( .Q(n1176), .DIN1(n1177), .DIN2(n728) );
    nor2s1 U420 ( .Q(n1178), .DIN1(n730), .DIN2(n1179) );
    nnd2s1 U421 ( .Q(n734), .DIN1(n1178), .DIN2(n1176) );
    nnd2s1 U422 ( .Q(n1180), .DIN1(n1181), .DIN2(n1182) );
    nor2s1 U423 ( .Q(n1183), .DIN1(n710), .DIN2(n1180) );
    nor2s1 U424 ( .Q(n1184), .DIN1(n712), .DIN2(n714) );
    nnd2s1 U425 ( .Q(n736), .DIN1(n1184), .DIN2(n1183) );
    nor2s1 U426 ( .Q(n1185), .DIN1(n716), .DIN2(n1186) );
    nnd2s1 U427 ( .Q(n1187), .DIN1(n1188), .DIN2(n967) );
    nnd2s1 U428 ( .Q(n737), .DIN1(n1189), .DIN2(n1185) );
    nor2s1 U429 ( .Q(n1190), .DIN1(n732), .DIN2(n735) );
    nnd2s1 U430 ( .Q(n739), .DIN1(n1190), .DIN2(n1191) );
    nnd2s1 U431 ( .Q(n740), .DIN1(n965), .DIN2(n1192) );
    nor2s1 U432 ( .Q(n562), .DIN1(n707), .DIN2(n738) );
    nor2s1 U433 ( .Q(n977), .DIN1(n798), .DIN2(n1193) );
    nnd2s1 U434 ( .Q(n1194), .DIN1(n1195), .DIN2(n1188) );
    nor2s1 U435 ( .Q(n1196), .DIN1(n768), .DIN2(n1194) );
    nor2s1 U436 ( .Q(n1197), .DIN1(n769), .DIN2(n770) );
    nnd2s1 U437 ( .Q(n777), .DIN1(n1197), .DIN2(n1196) );
    nor2s1 U438 ( .Q(n1198), .DIN1(n772), .DIN2(n774) );
    nor2s1 U439 ( .Q(n1199), .DIN1(n775), .DIN2(n1179) );
    nnd2s1 U440 ( .Q(n778), .DIN1(n1199), .DIN2(n1198) );
    nnd2s1 U441 ( .Q(n1200), .DIN1(n1201), .DIN2(n1202) );
    nor2s1 U442 ( .Q(n1203), .DIN1(n762), .DIN2(n1200) );
    nor2s1 U443 ( .Q(n1204), .DIN1(n763), .DIN2(n764) );
    nnd2s1 U444 ( .Q(n780), .DIN1(n1204), .DIN2(n1203) );
    nor2s1 U445 ( .Q(n1205), .DIN1(n765), .DIN2(n766) );
    nnd2s1 U446 ( .Q(n1206), .DIN1(n1205), .DIN2(n967) );
    nnd2s1 U447 ( .Q(n781), .DIN1(n1207), .DIN2(n1208) );
    nor2s1 U448 ( .Q(n1209), .DIN1(n776), .DIN2(n779) );
    nnd2s1 U449 ( .Q(n783), .DIN1(n1209), .DIN2(n1210) );
    nnd2s1 U450 ( .Q(n784), .DIN1(n965), .DIN2(n1211) );
    nor2s1 U451 ( .Q(n564), .DIN1(n760), .DIN2(n782) );
    nnd2s1 U452 ( .Q(n577), .DIN1(n968), .DIN2(n1005) );
    nor2s1 U453 ( .Q(n1212), .DIN1(n575), .DIN2(n758) );
    nor2s1 U454 ( .Q(n1213), .DIN1(n795), .DIN2(n797) );
    nor2s1 U455 ( .Q(n1214), .DIN1(n1164), .DIN2(n1215) );
    nnd2s1 U456 ( .Q(n1216), .DIN1(n1214), .DIN2(n1217) );
    nnd2s1 U457 ( .Q(n1218), .DIN1(n1219), .DIN2(n1220) );
    nor2s1 U458 ( .Q(n1221), .DIN1(n1216), .DIN2(n1218) );
    nnd2s1 U459 ( .Q(n1222), .DIN1(n1223), .DIN2(n1224) );
    nnd2s1 U460 ( .Q(n1225), .DIN1(n966), .DIN2(n1226) );
    nor2s1 U461 ( .Q(n1227), .DIN1(n1222), .DIN2(n1225) );
    nor2s1 U462 ( .Q(n1228), .DIN1(n785), .DIN2(n786) );
    nnd2s1 U463 ( .Q(n1229), .DIN1(n1228), .DIN2(n1230) );
    nnd2s1 U464 ( .Q(n1231), .DIN1(n1232), .DIN2(n1233) );
    nor2s1 U465 ( .Q(n1234), .DIN1(n1229), .DIN2(n1231) );
    nnd2s1 U466 ( .Q(n1235), .DIN1(n1236), .DIN2(n1237) );
    nnd2s1 U467 ( .Q(n1238), .DIN1(n967), .DIN2(n1239) );
    nor2s1 U468 ( .Q(n1240), .DIN1(n1235), .DIN2(n1238) );
    nnd2s1 U469 ( .Q(n1241), .DIN1(n1242), .DIN2(n1243) );
    nor2s1 U470 ( .Q(n1244), .DIN1(n790), .DIN2(n1241) );
    nor2s1 U471 ( .Q(n1245), .DIN1(n792), .DIN2(n1170) );
    nor2s1 U472 ( .Q(n1246), .DIN1(n1165), .DIN2(n1247) );
    nnd2s1 U473 ( .Q(n1248), .DIN1(n1246), .DIN2(n1239) );
    nnd2s1 U474 ( .Q(n1249), .DIN1(n1250), .DIN2(n1251) );
    nor2s1 U475 ( .Q(n1252), .DIN1(n1248), .DIN2(n1249) );
    nnd2s1 U476 ( .Q(n1253), .DIN1(n1254), .DIN2(n1255) );
    nnd2s1 U477 ( .Q(n1256), .DIN1(n966), .DIN2(n1257) );
    nor2s1 U478 ( .Q(n1258), .DIN1(n1253), .DIN2(n1256) );
    nor2s1 U479 ( .Q(n1259), .DIN1(n1260), .DIN2(n804) );
    nnd2s1 U480 ( .Q(n1261), .DIN1(n1259), .DIN2(n1262) );
    nnd2s1 U481 ( .Q(n1263), .DIN1(n1264), .DIN2(n1265) );
    nor2s1 U482 ( .Q(n1266), .DIN1(n1261), .DIN2(n1263) );
    nnd2s1 U483 ( .Q(n1267), .DIN1(n1268), .DIN2(n1269) );
    nnd2s1 U484 ( .Q(n1270), .DIN1(n967), .DIN2(n1271) );
    nor2s1 U485 ( .Q(n1272), .DIN1(n1267), .DIN2(n1270) );
    nor2s1 U486 ( .Q(n981), .DIN1(N97), .DIN2(N116) );
    nor2s1 U487 ( .Q(n980), .DIN1(N107), .DIN2(N87) );
    nnd2s1 U488 ( .Q(n841), .DIN1(n848), .DIN2(n773) );
    nnd2s1 U489 ( .Q(n842), .DIN1(n1273), .DIN2(N58) );
    nnd2s1 U490 ( .Q(n1274), .DIN1(n1275), .DIN2(n1276) );
    nnd2s1 U491 ( .Q(n1277), .DIN1(n1278), .DIN2(n1279) );
    nnd2s1 U492 ( .Q(n1280), .DIN1(n1281), .DIN2(n1282) );
    nor2s1 U493 ( .Q(n1283), .DIN1(n806), .DIN2(n1280) );
    nor2s1 U494 ( .Q(n1284), .DIN1(n807), .DIN2(n1170) );
    nor2s1 U495 ( .Q(n1285), .DIN1(n971), .DIN2(n821) );
    nor2s1 U496 ( .Q(n1286), .DIN1(n1186), .DIN2(n1287) );
    nnd2s1 U497 ( .Q(n1288), .DIN1(n1286), .DIN2(n1208) );
    nnd2s1 U498 ( .Q(n1289), .DIN1(n1290), .DIN2(n1291) );
    nor2s1 U499 ( .Q(n1292), .DIN1(n1288), .DIN2(n1289) );
    nnd2s1 U500 ( .Q(n1293), .DIN1(n1294), .DIN2(n1295) );
    nnd2s1 U501 ( .Q(n1296), .DIN1(n966), .DIN2(n1297) );
    nor2s1 U502 ( .Q(n1298), .DIN1(n1293), .DIN2(n1296) );
    nor2s1 U503 ( .Q(n1299), .DIN1(n1300), .DIN2(n817) );
    nnd2s1 U504 ( .Q(n1301), .DIN1(n1299), .DIN2(n1302) );
    nnd2s1 U505 ( .Q(n1303), .DIN1(n1304), .DIN2(n1305) );
    nor2s1 U506 ( .Q(n1306), .DIN1(n1301), .DIN2(n1303) );
    nnd2s1 U507 ( .Q(n1307), .DIN1(n1308), .DIN2(n1309) );
    nnd2s1 U508 ( .Q(n1310), .DIN1(n967), .DIN2(n1311) );
    nor2s1 U509 ( .Q(n1312), .DIN1(n1307), .DIN2(n1310) );
    nor2s1 U510 ( .Q(n1313), .DIN1(n982), .DIN2(n812) );
    nnd2s1 U511 ( .Q(n1314), .DIN1(n1315), .DIN2(n1316) );
    nor2s1 U512 ( .Q(n1317), .DIN1(n818), .DIN2(n1314) );
    nor2s1 U513 ( .Q(n1318), .DIN1(n819), .DIN2(n1170) );
    nnd2s1 U514 ( .Q(n1319), .DIN1(n1320), .DIN2(n1321) );
    nnd2s1 U515 ( .Q(n1322), .DIN1(n1323), .DIN2(n1324) );
    nor2s1 U516 ( .Q(n1325), .DIN1(n1326), .DIN2(n744) );
    nnd2s1 U517 ( .Q(n1327), .DIN1(n1325), .DIN2(n1328) );
    nnd2s1 U518 ( .Q(n1329), .DIN1(n1330), .DIN2(n1331) );
    nor2s1 U519 ( .Q(n1332), .DIN1(n1327), .DIN2(n1329) );
    nnd2s1 U520 ( .Q(n1333), .DIN1(n1334), .DIN2(n1335) );
    nnd2s1 U521 ( .Q(n1336), .DIN1(n966), .DIN2(n1337) );
    nor2s1 U522 ( .Q(n1338), .DIN1(n1333), .DIN2(n1336) );
    nor2s1 U523 ( .Q(n1339), .DIN1(n741), .DIN2(n743) );
    nnd2s1 U524 ( .Q(n1340), .DIN1(n1339), .DIN2(n1341) );
    nnd2s1 U525 ( .Q(n1342), .DIN1(n1343), .DIN2(n1344) );
    nor2s1 U526 ( .Q(n1345), .DIN1(n1340), .DIN2(n1342) );
    nnd2s1 U527 ( .Q(n1346), .DIN1(n1347), .DIN2(n1348) );
    nnd2s1 U528 ( .Q(n1349), .DIN1(n967), .DIN2(n1350) );
    nor2s1 U529 ( .Q(n1351), .DIN1(n1346), .DIN2(n1349) );
    nnd2s1 U530 ( .Q(n1352), .DIN1(n1353), .DIN2(n1354) );
    nor2s1 U531 ( .Q(n1355), .DIN1(n745), .DIN2(n1352) );
    nor2s1 U532 ( .Q(n1356), .DIN1(n746), .DIN2(n1170) );
    nor2s1 U533 ( .Q(n1357), .DIN1(n1358), .DIN2(n754) );
    nnd2s1 U534 ( .Q(n1359), .DIN1(n1357), .DIN2(n1360) );
    nnd2s1 U535 ( .Q(n1361), .DIN1(n1362), .DIN2(n1363) );
    nor2s1 U536 ( .Q(n1364), .DIN1(n1359), .DIN2(n1361) );
    nnd2s1 U537 ( .Q(n1365), .DIN1(n1366), .DIN2(n1367) );
    nnd2s1 U538 ( .Q(n1368), .DIN1(n966), .DIN2(n1369) );
    nor2s1 U539 ( .Q(n1370), .DIN1(n1365), .DIN2(n1368) );
    nor2s1 U540 ( .Q(n1371), .DIN1(n751), .DIN2(n753) );
    nnd2s1 U541 ( .Q(n1372), .DIN1(n1371), .DIN2(n1373) );
    nnd2s1 U542 ( .Q(n1374), .DIN1(n1375), .DIN2(n1376) );
    nor2s1 U543 ( .Q(n1377), .DIN1(n1372), .DIN2(n1374) );
    nnd2s1 U544 ( .Q(n1378), .DIN1(n1379), .DIN2(n1380) );
    nnd2s1 U545 ( .Q(n1381), .DIN1(n967), .DIN2(n1195) );
    nor2s1 U546 ( .Q(n1382), .DIN1(n1378), .DIN2(n1381) );
    nnd2s1 U547 ( .Q(n1383), .DIN1(n1384), .DIN2(n1385) );
    nor2s1 U548 ( .Q(n1386), .DIN1(n755), .DIN2(n1383) );
    nor2s1 U549 ( .Q(n1387), .DIN1(n756), .DIN2(n1170) );
    nnd2s1 U550 ( .Q(n1388), .DIN1(n1389), .DIN2(n1390) );
    nor2s1 U551 ( .Q(n1391), .DIN1(n1392), .DIN2(n1393) );
    nnd2s1 U552 ( .Q(n1394), .DIN1(n1395), .DIN2(n1396) );
    nnd2s1 U553 ( .Q(n1397), .DIN1(n1398), .DIN2(n1399) );
    nnd2s1 U554 ( .Q(n1400), .DIN1(n1401), .DIN2(n1402) );
    nor2s1 U555 ( .Q(n586), .DIN1(n1397), .DIN2(n1400) );
    nnd2s1 U556 ( .Q(n1403), .DIN1(n1404), .DIN2(n1405) );
    nnd2s1 U557 ( .Q(n1406), .DIN1(n1407), .DIN2(n1408) );
    nor2s1 U558 ( .Q(n585), .DIN1(n1403), .DIN2(n1406) );
    nnd2s1 U559 ( .Q(n823), .DIN1(n1402), .DIN2(n1398) );
    nor2s1 U560 ( .Q(n584), .DIN1(n1409), .DIN2(n822) );
    nnd2s1 U561 ( .Q(n1073), .DIN1(N50), .DIN2(N58) );
    nor2s1 U562 ( .Q(n1410), .DIN1(N13), .DIN2(n824) );
    nnd2s1 U563 ( .Q(n1411), .DIN1(n1412), .DIN2(n1413) );
    nor2s1 U564 ( .Q(n1414), .DIN1(n930), .DIN2(n579) );
    nor2s1 U565 ( .Q(n1415), .DIN1(n828), .DIN2(n829) );
    nor2s1 U566 ( .Q(n1416), .DIN1(n830), .DIN2(n831) );
    nnd2s1 U567 ( .Q(n838), .DIN1(n1416), .DIN2(n1415) );
    nor2s1 U568 ( .Q(n1417), .DIN1(n832), .DIN2(n833) );
    nor2s1 U569 ( .Q(n1418), .DIN1(n834), .DIN2(n835) );
    nnd2s1 U570 ( .Q(n839), .DIN1(n1418), .DIN2(n1417) );
    nnd2s1 U571 ( .Q(n605), .DIN1(n773), .DIN2(n617) );
    nor2s1 U572 ( .Q(n863), .DIN1(n858), .DIN2(n852) );
    nnd2s1 U573 ( .Q(n1419), .DIN1(n862), .DIN2(n858) );
    nor2s1 U574 ( .Q(n1420), .DIN1(N77), .DIN2(n1421) );
    nor2s1 U575 ( .Q(n1422), .DIN1(n617), .DIN2(n1419) );
    nor2s1 U576 ( .Q(n882), .DIN1(n1420), .DIN2(n1422) );
    nnd2s1 U577 ( .Q(n1423), .DIN1(n1091), .DIN2(n1090) );
    nor2s1 U578 ( .Q(n1424), .DIN1(n1425), .DIN2(n872) );
    nor2s1 U579 ( .Q(n1426), .DIN1(n871), .DIN2(n1423) );
    nor2s1 U580 ( .Q(n1427), .DIN1(n1424), .DIN2(n1426) );
    nor2s1 U581 ( .Q(n1428), .DIN1(N179), .DIN2(n1423) );
    nor2s1 U582 ( .Q(n1429), .DIN1(N169), .DIN2(n1425) );
    nor2s1 U583 ( .Q(n880), .DIN1(n1428), .DIN2(n1429) );
    nor2s1 U584 ( .Q(n1430), .DIN1(n923), .DIN2(n1431) );
    nnd2s1 U585 ( .Q(n1432), .DIN1(n862), .DIN2(n1433) );
    nor2s1 U586 ( .Q(n1434), .DIN1(N87), .DIN2(n1421) );
    nor2s1 U587 ( .Q(n1435), .DIN1(n631), .DIN2(n1432) );
    nor2s1 U588 ( .Q(n901), .DIN1(n1434), .DIN2(n1435) );
    nor2s1 U589 ( .Q(n1436), .DIN1(n1111), .DIN2(n872) );
    nor2s1 U590 ( .Q(n1437), .DIN1(n871), .DIN2(n897) );
    nor2s1 U591 ( .Q(n1438), .DIN1(n1436), .DIN2(n1437) );
    nor2s1 U592 ( .Q(n1439), .DIN1(N179), .DIN2(n897) );
    nor2s1 U593 ( .Q(n1440), .DIN1(N169), .DIN2(n1111) );
    nor2s1 U594 ( .Q(n1441), .DIN1(n1439), .DIN2(n1440) );
    nor2s1 U595 ( .Q(n1442), .DIN1(N97), .DIN2(n1421) );
    nor2s1 U596 ( .Q(n1443), .DIN1(n647), .DIN2(n1432) );
    nor2s1 U597 ( .Q(n907), .DIN1(n1442), .DIN2(n1443) );
    nor2s1 U598 ( .Q(n1444), .DIN1(n1114), .DIN2(n872) );
    nor2s1 U599 ( .Q(n1445), .DIN1(n871), .DIN2(n903) );
    nor2s1 U600 ( .Q(n1446), .DIN1(n1444), .DIN2(n1445) );
    nor2s1 U601 ( .Q(n1447), .DIN1(N179), .DIN2(n903) );
    nor2s1 U602 ( .Q(n1448), .DIN1(N169), .DIN2(n1114) );
    nor2s1 U603 ( .Q(n920), .DIN1(n1447), .DIN2(n1448) );
    nor2s1 U604 ( .Q(n1449), .DIN1(N107), .DIN2(n1421) );
    nor2s1 U605 ( .Q(n1450), .DIN1(n655), .DIN2(n1432) );
    nor2s1 U606 ( .Q(n1451), .DIN1(n1449), .DIN2(n1450) );
    nnd2s1 U607 ( .Q(n1106), .DIN1(n1451), .DIN2(n1452) );
    nor2s1 U608 ( .Q(n1453), .DIN1(N116), .DIN2(n1421) );
    nor2s1 U609 ( .Q(n1454), .DIN1(n664), .DIN2(n1432) );
    nor2s1 U610 ( .Q(n928), .DIN1(n1453), .DIN2(n1454) );
    nor2s1 U611 ( .Q(n1455), .DIN1(n1112), .DIN2(n872) );
    nor2s1 U612 ( .Q(n1456), .DIN1(n871), .DIN2(n894) );
    nor2s1 U613 ( .Q(n1457), .DIN1(n1455), .DIN2(n1456) );
    nor2s1 U614 ( .Q(n1458), .DIN1(N179), .DIN2(n894) );
    nor2s1 U615 ( .Q(n1459), .DIN1(N169), .DIN2(n1112) );
    nor2s1 U616 ( .Q(n918), .DIN1(n1458), .DIN2(n1459) );
    nor2s1 U617 ( .Q(n1460), .DIN1(N68), .DIN2(n1421) );
    nor2s1 U618 ( .Q(n1461), .DIN1(n644), .DIN2(n1419) );
    nor2s1 U619 ( .Q(n1462), .DIN1(n1460), .DIN2(n1461) );
    nnd2s1 U620 ( .Q(n1463), .DIN1(n1121), .DIN2(n1120) );
    nnd2s1 U621 ( .Q(n1136), .DIN1(n1462), .DIN2(n1464) );
    nor2s1 U622 ( .Q(n1465), .DIN1(n923), .DIN2(n1122) );
    nor2s1 U623 ( .Q(n1466), .DIN1(n1467), .DIN2(n696) );
    nor2s1 U624 ( .Q(n1468), .DIN1(N58), .DIN2(n1421) );
    nor2s1 U625 ( .Q(n1469), .DIN1(n771), .DIN2(n1419) );
    nor2s1 U626 ( .Q(n874), .DIN1(n1468), .DIN2(n1469) );
    nnd2s1 U627 ( .Q(n1470), .DIN1(n1130), .DIN2(n1129) );
    nor2s1 U628 ( .Q(n1471), .DIN1(n1472), .DIN2(n872) );
    nor2s1 U629 ( .Q(n1473), .DIN1(n871), .DIN2(n1470) );
    nor2s1 U630 ( .Q(n1474), .DIN1(n1471), .DIN2(n1473) );
    nor2s1 U631 ( .Q(n1475), .DIN1(N179), .DIN2(n1470) );
    nor2s1 U632 ( .Q(n1476), .DIN1(N169), .DIN2(n1472) );
    nor2s1 U633 ( .Q(n943), .DIN1(n1475), .DIN2(n1476) );
    nor2s1 U634 ( .Q(n1477), .DIN1(n887), .DIN2(n1478) );
    nor2s1 U635 ( .Q(n1479), .DIN1(n1124), .DIN2(n1123) );
    nnd2s1 U636 ( .Q(n1480), .DIN1(n1134), .DIN2(n1133) );
    nor2s1 U637 ( .Q(n1481), .DIN1(N50), .DIN2(n1421) );
    nor2s1 U638 ( .Q(n1482), .DIN1(n773), .DIN2(n1419) );
    nor2s1 U639 ( .Q(n1483), .DIN1(n1481), .DIN2(n1482) );
    nnd2s1 U640 ( .Q(n1484), .DIN1(n1483), .DIN2(n1485) );
    nnd2s1 U641 ( .Q(n1486), .DIN1(n637), .DIN2(n1484) );
    nor2s1 U642 ( .Q(n1487), .DIN1(n949), .DIN2(n1488) );
    nor2s1 U643 ( .Q(n1489), .DIN1(n937), .DIN2(n993) );
    nnd2s1 U644 ( .Q(n1490), .DIN1(n798), .DIN2(n906) );
    nor2s1 U645 ( .Q(n1491), .DIN1(n923), .DIN2(n1492) );
    nnd2s1 U646 ( .Q(n1493), .DIN1(n798), .DIN2(n1106) );
    nor2s1 U647 ( .Q(n1494), .DIN1(n971), .DIN2(n968) );
    nnd2s1 U648 ( .Q(n1495), .DIN1(n810), .DIN2(n1496) );
    nor2s1 U649 ( .Q(n1497), .DIN1(n1057), .DIN2(n1495) );
    nnd2s1 U650 ( .Q(n1498), .DIN1(n1495), .DIN2(n1057) );
    nor2s1 U651 ( .Q(n761), .DIN1(n1497), .DIN2(n1499) );
    nor2s1 U652 ( .Q(n1500), .DIN1(N107), .DIN2(n664) );
    nor2s1 U653 ( .Q(n1501), .DIN1(N116), .DIN2(n655) );
    nor2s1 U654 ( .Q(n1502), .DIN1(n1500), .DIN2(n1501) );
    nor2s1 U655 ( .Q(n1503), .DIN1(N87), .DIN2(n647) );
    nor2s1 U656 ( .Q(n1504), .DIN1(N97), .DIN2(n631) );
    nor2s1 U657 ( .Q(n1505), .DIN1(n1503), .DIN2(n1504) );
    nor2s1 U658 ( .Q(n1506), .DIN1(N97), .DIN2(n974) );
    nor2s1 U659 ( .Q(n1507), .DIN1(n1508), .DIN2(n846) );
    nor2s1 U660 ( .Q(n1509), .DIN1(n1506), .DIN2(n1507) );
    nor2s1 U661 ( .Q(n1510), .DIN1(n923), .DIN2(n1511) );
    nnd2s1 U662 ( .Q(n1512), .DIN1(n1213), .DIN2(n1212) );
    nor2s1 U663 ( .Q(n1513), .DIN1(n794), .DIN2(n1512) );
    nnd2s1 U664 ( .Q(n1514), .DIN1(n1512), .DIN2(n794) );
    nor2s1 U665 ( .Q(n1515), .DIN1(n1513), .DIN2(n1516) );
    nor2s1 U666 ( .Q(n1517), .DIN1(N264), .DIN2(n836) );
    nor2s1 U667 ( .Q(n1518), .DIN1(N270), .DIN2(n684) );
    nor2s1 U668 ( .Q(n1519), .DIN1(n1517), .DIN2(n1518) );
    nor2s1 U669 ( .Q(n1520), .DIN1(N250), .DIN2(n680) );
    nor2s1 U670 ( .Q(n1521), .DIN1(N257), .DIN2(n671) );
    nor2s1 U671 ( .Q(n1522), .DIN1(n1520), .DIN2(n1521) );
    nnd2s1 U672 ( .Q(n1523), .DIN1(n810), .DIN2(n939) );
    nor2s1 U673 ( .Q(n1524), .DIN1(n1496), .DIN2(n1523) );
    nor2s1 U674 ( .Q(n1525), .DIN1(n811), .DIN2(n1012) );
    nor2s1 U675 ( .Q(n566), .DIN1(n1524), .DIN2(n1525) );
    nor2s1 U676 ( .Q(n1526), .DIN1(N50), .DIN2(n771) );
    nor2s1 U677 ( .Q(n1527), .DIN1(N58), .DIN2(n773) );
    nor2s1 U678 ( .Q(n1528), .DIN1(n1526), .DIN2(n1527) );
    nor2s1 U679 ( .Q(n1529), .DIN1(N68), .DIN2(n617) );
    nor2s1 U680 ( .Q(n1530), .DIN1(N77), .DIN2(n644) );
    nor2s1 U681 ( .Q(n1531), .DIN1(n1529), .DIN2(n1530) );
    nnd2s1 U682 ( .Q(n1532), .DIN1(n939), .DIN2(n748) );
    nor2s1 U683 ( .Q(n1533), .DIN1(n1534), .DIN2(n1532) );
    nor2s1 U684 ( .Q(n1535), .DIN1(n749), .DIN2(n993) );
    nor2s1 U685 ( .Q(n558), .DIN1(n1533), .DIN2(n1535) );
    nor2s1 U686 ( .Q(n1536), .DIN1(n757), .DIN2(n970) );
    nor2s1 U687 ( .Q(n1537), .DIN1(n810), .DIN2(n936) );
    nor2s1 U688 ( .Q(n1538), .DIN1(n1536), .DIN2(n1537) );
    nor2s1 U689 ( .Q(n1539), .DIN1(n1394), .DIN2(n1540) );
    nor2s1 U690 ( .Q(n1541), .DIN1(n1388), .DIN2(n1542) );
    nor2s1 U691 ( .Q(N5361), .DIN1(n1539), .DIN2(n1541) );
    nor2s1 U692 ( .Q(n1543), .DIN1(n1402), .DIN2(n1544) );
    nnd2s1 U693 ( .Q(n1545), .DIN1(n1546), .DIN2(n1547) );
    nnd2s1 U694 ( .Q(n1548), .DIN1(n924), .DIN2(n933) );
    nnd2s1 U695 ( .Q(n1549), .DIN1(N330), .DIN2(n1550) );
    nnd2s1 U696 ( .Q(n1551), .DIN1(n1552), .DIN2(n1553) );
    nnd2s1 U697 ( .Q(n1554), .DIN1(N116), .DIN2(n1555) );
    nor2s1 U698 ( .Q(n1556), .DIN1(n1078), .DIN2(n1551) );
    nor2s1 U699 ( .Q(n1557), .DIN1(n849), .DIN2(n1554) );
    nor2s1 U700 ( .Q(n589), .DIN1(n1556), .DIN2(n1557) );
    nnd2s1 U701 ( .Q(n1558), .DIN1(n1273), .DIN2(n708) );
    nor2s1 U702 ( .Q(n1559), .DIN1(n853), .DIN2(n1558) );
    nor2s1 U703 ( .Q(n1560), .DIN1(N1), .DIN2(n810) );
    nor2s1 U704 ( .Q(n593), .DIN1(n1559), .DIN2(n1560) );
    nnd2s1 U705 ( .Q(n922), .DIN1(n1109), .DIN2(n1108) );
    hi1s1 U706 ( .Q(n798), .DIN(n923) );
    hi1s1 U707 ( .Q(n624), .DIN(n963) );
    hi1s1 U708 ( .Q(n708), .DIN(n939) );
    hi1s1 U709 ( .Q(n1078), .DIN(n849) );
    nnd2s1 U710 ( .Q(n1089), .DIN1(n864), .DIN2(N274) );
    nnd2s1 U711 ( .Q(n1094), .DIN1(n891), .DIN2(N274) );
    hi1s1 U712 ( .Q(n635), .DIN(n857) );
    hi1s1 U713 ( .Q(n1179), .DIN(n966) );
    hi1s1 U714 ( .Q(n791), .DIN(n975) );
    hi1s1 U715 ( .Q(n848), .DIN(n982) );
    nor2s1 U716 ( .Q(n964), .DIN1(n643), .DIN2(N169) );
    hi1s1 U717 ( .Q(n628), .DIN(n788) );
    nnd2s1 U718 ( .Q(n940), .DIN1(n1137), .DIN2(N13) );
    hi1s1 U719 ( .Q(n1561), .DIN(n750) );
    hi1s1 U720 ( .Q(n1170), .DIN(n965) );
    nnd2s1 U721 ( .Q(n861), .DIN1(N33), .DIN2(n854) );
    hi1s1 U722 ( .Q(n640), .DIN(n609) );
    nnd2s1 U723 ( .Q(n1562), .DIN1(n857), .DIN2(n723) );
    nnd2s1 U724 ( .Q(n1485), .DIN1(n1135), .DIN2(n1562) );
    hi1s1 U725 ( .Q(n1563), .DIN(n1484) );
    nor2s1 U726 ( .Q(n869), .DIN1(n866), .DIN2(n856) );
    nor2s1 U727 ( .Q(n865), .DIN1(N41), .DIN2(N45) );
    nnd2s1 U728 ( .Q(n1132), .DIN1(N226), .DIN2(n867) );
    hi1s1 U729 ( .Q(n1564), .DIN(n1480) );
    hi1s1 U730 ( .Q(n803), .DIN(n742) );
    nnd2s1 U731 ( .Q(n1155), .DIN1(n803), .DIN2(N283) );
    hi1s1 U732 ( .Q(n1565), .DIN(n805) );
    nor2s1 U733 ( .Q(n1326), .DIN1(n805), .DIN2(n771) );
    hi1s1 U734 ( .Q(n1154), .DIN(n1326) );
    hi1s1 U735 ( .Q(n1566), .DIN(n711) );
    nnd2s1 U736 ( .Q(n1158), .DIN1(n1566), .DIN2(N87) );
    hi1s1 U737 ( .Q(n727), .DIN(n713) );
    nnd2s1 U738 ( .Q(n1157), .DIN1(n727), .DIN2(N97) );
    hi1s1 U739 ( .Q(n1567), .DIN(n715) );
    nnd2s1 U740 ( .Q(n1162), .DIN1(n1567), .DIN2(N107) );
    hi1s1 U741 ( .Q(n1568), .DIN(n717) );
    nnd2s1 U742 ( .Q(n1161), .DIN1(n1568), .DIN2(N116) );
    hi1s1 U743 ( .Q(n1569), .DIN(n722) );
    nor2s1 U744 ( .Q(n1165), .DIN1(n722), .DIN2(n617) );
    nor2s1 U745 ( .Q(n962), .DIN1(n643), .DIN2(n960) );
    hi1s1 U746 ( .Q(n719), .DIN(n961) );
    nor2s1 U747 ( .Q(n1164), .DIN1(n719), .DIN2(n644) );
    nnd2s1 U748 ( .Q(n1141), .DIN1(N124), .DIN2(n803) );
    nnd2s1 U749 ( .Q(n1140), .DIN1(N159), .DIN2(n1565) );
    nnd2s1 U750 ( .Q(n1144), .DIN1(N150), .DIN2(n961) );
    nnd2s1 U751 ( .Q(n1143), .DIN1(N143), .DIN2(n1569) );
    nnd2s1 U752 ( .Q(n1148), .DIN1(N137), .DIN2(n1566) );
    nnd2s1 U753 ( .Q(n1147), .DIN1(N132), .DIN2(n727) );
    nnd2s1 U754 ( .Q(n1151), .DIN1(N128), .DIN2(n1567) );
    nnd2s1 U755 ( .Q(n1150), .DIN1(N125), .DIN2(n1568) );
    nnd2s1 U756 ( .Q(n560), .DIN1(n1169), .DIN2(n1168) );
    nnd2s1 U757 ( .Q(n1128), .DIN1(N232), .DIN2(n867) );
    hi1s1 U758 ( .Q(n1472), .DIN(n1470) );
    nnd2s1 U759 ( .Q(n875), .DIN1(n1126), .DIN2(n1125) );
    hi1s1 U760 ( .Q(n1478), .DIN(n873) );
    hi1s1 U761 ( .Q(n701), .DIN(n638) );
    nnd2s1 U762 ( .Q(n877), .DIN1(n1474), .DIN2(n1478) );
    nnd2s1 U763 ( .Q(n1464), .DIN1(n1117), .DIN2(n1116) );
    hi1s1 U764 ( .Q(n1122), .DIN(n1136) );
    nnd2s1 U765 ( .Q(n1119), .DIN1(N238), .DIN2(n867) );
    hi1s1 U766 ( .Q(n1570), .DIN(n1463) );
    nnd2s1 U767 ( .Q(n883), .DIN1(n1086), .DIN2(n1084) );
    hi1s1 U768 ( .Q(n1431), .DIN(n881) );
    nnd2s1 U769 ( .Q(n1088), .DIN1(N244), .DIN2(n867) );
    hi1s1 U770 ( .Q(n1425), .DIN(n1423) );
    nnd2s1 U771 ( .Q(n885), .DIN1(n1427), .DIN2(n1431) );
    nnd2s1 U772 ( .Q(n1571), .DIN1(n857), .DIN2(n644) );
    nnd2s1 U773 ( .Q(n902), .DIN1(n1101), .DIN2(n1571) );
    nnd2s1 U774 ( .Q(n1433), .DIN1(N33), .DIN2(n853) );
    hi1s1 U775 ( .Q(n1511), .DIN(n900) );
    hi1s1 U776 ( .Q(n892), .DIN(n890) );
    hi1s1 U777 ( .Q(n1111), .DIN(n897) );
    nnd2s1 U778 ( .Q(n914), .DIN1(n1441), .DIN2(n900) );
    hi1s1 U779 ( .Q(n1110), .DIN(n914) );
    nnd2s1 U780 ( .Q(n915), .DIN1(n1438), .DIN2(n1511) );
    hi1s1 U781 ( .Q(n917), .DIN(n674) );
    nnd2s1 U782 ( .Q(n1100), .DIN1(N257), .DIN2(n893) );
    hi1s1 U783 ( .Q(n1114), .DIN(n903) );
    nnd2s1 U784 ( .Q(n908), .DIN1(n1098), .DIN2(n1097) );
    hi1s1 U785 ( .Q(n1572), .DIN(n906) );
    nnd2s1 U786 ( .Q(n929), .DIN1(n1103), .DIN2(n1102) );
    hi1s1 U787 ( .Q(n1492), .DIN(n919) );
    nnd2s1 U788 ( .Q(n1105), .DIN1(N270), .DIN2(n893) );
    hi1s1 U789 ( .Q(n1112), .DIN(n894) );
    nnd2s1 U790 ( .Q(n913), .DIN1(n1446), .DIN2(n1572) );
    nnd2s1 U791 ( .Q(n1452), .DIN1(n1096), .DIN2(n1095) );
    hi1s1 U792 ( .Q(n1193), .DIN(n1106) );
    nnd2s1 U793 ( .Q(n1093), .DIN1(N264), .DIN2(n893) );
    hi1s1 U794 ( .Q(n1113), .DIN(n909) );
    nnd2s1 U795 ( .Q(n931), .DIN1(n1457), .DIN2(n1492) );
    nnd2s1 U796 ( .Q(n1573), .DIN1(n946), .DIN2(N330) );
    nnd2s1 U797 ( .Q(n927), .DIN1(n1574), .DIN2(n1484) );
    hi1s1 U798 ( .Q(n597), .DIN(n925) );
    nor2s1 U799 ( .Q(n935), .DIN1(n599), .DIN2(n921) );
    nor2s1 U800 ( .Q(n1575), .DIN1(n932), .DIN2(n599) );
    nnd2s1 U801 ( .Q(n1576), .DIN1(n998), .DIN2(n1534) );
    nnd2s1 U802 ( .Q(n1577), .DIN1(n748), .DIN2(n1576) );
    nnd2s1 U803 ( .Q(n1578), .DIN1(n939), .DIN2(n1577) );
    nnd2s1 U804 ( .Q(n1579), .DIN1(n1561), .DIN2(n1578) );
    nnd2s1 U805 ( .Q(n561), .DIN1(n1580), .DIN2(n1579) );
    hi1s1 U806 ( .Q(n1398), .DIN(N5120) );
    nnd2s1 U807 ( .Q(n1182), .DIN1(n803), .DIN2(N294) );
    nor2s1 U808 ( .Q(n1358), .DIN1(n805), .DIN2(n644) );
    hi1s1 U809 ( .Q(n1181), .DIN(n1358) );
    nor2s1 U810 ( .Q(n1186), .DIN1(n722), .DIN2(n631) );
    nnd2s1 U811 ( .Q(n1188), .DIN1(n961), .DIN2(N77) );
    nnd2s1 U812 ( .Q(n1173), .DIN1(N125), .DIN2(n803) );
    nnd2s1 U813 ( .Q(n1172), .DIN1(n1565), .DIN2(N50) );
    nnd2s1 U814 ( .Q(n1191), .DIN1(n1581), .DIN2(n771) );
    nnd2s1 U815 ( .Q(n1192), .DIN1(n788), .DIN2(n571) );
    nnd2s1 U816 ( .Q(n563), .DIN1(n998), .DIN2(n750) );
    hi1s1 U817 ( .Q(n1402), .DIN(N5102) );
    nnd2s1 U818 ( .Q(n1341), .DIN1(n1566), .DIN2(N107) );
    nnd2s1 U819 ( .Q(n1344), .DIN1(n727), .DIN2(N116) );
    nnd2s1 U820 ( .Q(n1343), .DIN1(n1567), .DIN2(N283) );
    nnd2s1 U821 ( .Q(n1348), .DIN1(n1568), .DIN2(N294) );
    nor2s1 U822 ( .Q(n1247), .DIN1(n719), .DIN2(n631) );
    hi1s1 U823 ( .Q(n1347), .DIN(n1247) );
    nnd2s1 U824 ( .Q(n1350), .DIN1(n1565), .DIN2(N77) );
    nnd2s1 U825 ( .Q(n1328), .DIN1(n961), .DIN2(N50) );
    nnd2s1 U826 ( .Q(n1331), .DIN1(N159), .DIN2(n1569) );
    nnd2s1 U827 ( .Q(n1330), .DIN1(N150), .DIN2(n1566) );
    nnd2s1 U828 ( .Q(n1335), .DIN1(N143), .DIN2(n727) );
    nnd2s1 U829 ( .Q(n1334), .DIN1(N137), .DIN2(n1567) );
    nnd2s1 U830 ( .Q(n1337), .DIN1(N132), .DIN2(n1568) );
    nnd2s1 U831 ( .Q(n1354), .DIN1(n1338), .DIN2(n1332) );
    nnd2s1 U832 ( .Q(n1353), .DIN1(n1351), .DIN2(n1345) );
    nnd2s1 U833 ( .Q(n559), .DIN1(n1356), .DIN2(n1355) );
    hi1s1 U834 ( .Q(n1399), .DIN(N5121) );
    nnd2s1 U835 ( .Q(n1373), .DIN1(n1566), .DIN2(N116) );
    nnd2s1 U836 ( .Q(n1376), .DIN1(n727), .DIN2(N283) );
    nnd2s1 U837 ( .Q(n1375), .DIN1(n1567), .DIN2(N294) );
    nnd2s1 U838 ( .Q(n1380), .DIN1(n1568), .DIN2(N303) );
    nor2s1 U839 ( .Q(n1287), .DIN1(n719), .DIN2(n647) );
    hi1s1 U840 ( .Q(n1379), .DIN(n1287) );
    nnd2s1 U841 ( .Q(n1195), .DIN1(n1565), .DIN2(N87) );
    nnd2s1 U842 ( .Q(n1360), .DIN1(n961), .DIN2(N58) );
    nnd2s1 U843 ( .Q(n1363), .DIN1(n1569), .DIN2(N50) );
    nnd2s1 U844 ( .Q(n1362), .DIN1(N159), .DIN2(n1566) );
    nnd2s1 U845 ( .Q(n1367), .DIN1(N150), .DIN2(n727) );
    nnd2s1 U846 ( .Q(n1366), .DIN1(N143), .DIN2(n1567) );
    nnd2s1 U847 ( .Q(n1369), .DIN1(N137), .DIN2(n1568) );
    nnd2s1 U848 ( .Q(n1385), .DIN1(n1370), .DIN2(n1364) );
    nnd2s1 U849 ( .Q(n1384), .DIN1(n1382), .DIN2(n1377) );
    nnd2s1 U850 ( .Q(n568), .DIN1(n1387), .DIN2(n1386) );
    nnd2s1 U851 ( .Q(n569), .DIN1(n1582), .DIN2(n1538) );
    hi1s1 U852 ( .Q(n1404), .DIN(N4944) );
    nnd2s1 U853 ( .Q(n973), .DIN1(n808), .DIN2(n968) );
    hi1s1 U854 ( .Q(n595), .DIN(n972) );
    hi1s1 U855 ( .Q(n971), .DIN(n969) );
    nnd2s1 U856 ( .Q(n1202), .DIN1(N322), .DIN2(n803) );
    nnd2s1 U857 ( .Q(n1201), .DIN1(n961), .DIN2(N116) );
    nnd2s1 U858 ( .Q(n1208), .DIN1(n1565), .DIN2(N107) );
    hi1s1 U859 ( .Q(n846), .DIN(n974) );
    nnd2s1 U860 ( .Q(n984), .DIN1(n1505), .DIN2(n1583) );
    nnd2s1 U861 ( .Q(n985), .DIN1(n1502), .DIN2(n1584) );
    hi1s1 U862 ( .Q(n1508), .DIN(n983) );
    nnd2s1 U863 ( .Q(n1585), .DIN1(n1509), .DIN2(n628) );
    nnd2s1 U864 ( .Q(n1210), .DIN1(n975), .DIN2(n1585) );
    nnd2s1 U865 ( .Q(n1211), .DIN1(n976), .DIN2(n759) );
    nnd2s1 U866 ( .Q(n565), .DIN1(n1057), .DIN2(n750) );
    hi1s1 U867 ( .Q(n1401), .DIN(N5078) );
    nnd2s1 U868 ( .Q(n1230), .DIN1(n1569), .DIN2(N116) );
    nnd2s1 U869 ( .Q(n1233), .DIN1(n1566), .DIN2(N283) );
    nnd2s1 U870 ( .Q(n1232), .DIN1(n727), .DIN2(N294) );
    nnd2s1 U871 ( .Q(n1237), .DIN1(n1567), .DIN2(N303) );
    nnd2s1 U872 ( .Q(n1236), .DIN1(N311), .DIN2(n1568) );
    nnd2s1 U873 ( .Q(n1239), .DIN1(n1565), .DIN2(N97) );
    nnd2s1 U874 ( .Q(n1217), .DIN1(N137), .DIN2(n803) );
    nnd2s1 U875 ( .Q(n1220), .DIN1(n1569), .DIN2(N58) );
    nnd2s1 U876 ( .Q(n1219), .DIN1(n1566), .DIN2(N50) );
    nnd2s1 U877 ( .Q(n1224), .DIN1(N159), .DIN2(n727) );
    nnd2s1 U878 ( .Q(n1223), .DIN1(N150), .DIN2(n1567) );
    nnd2s1 U879 ( .Q(n1226), .DIN1(N143), .DIN2(n1568) );
    nnd2s1 U880 ( .Q(n987), .DIN1(n1522), .DIN2(n1586) );
    nnd2s1 U881 ( .Q(n988), .DIN1(n1519), .DIN2(n1587) );
    nnd2s1 U882 ( .Q(n1243), .DIN1(n1227), .DIN2(n1221) );
    nnd2s1 U883 ( .Q(n1242), .DIN1(n1240), .DIN2(n1234) );
    nnd2s1 U884 ( .Q(n587), .DIN1(n1245), .DIN2(n1244) );
    nnd2s1 U885 ( .Q(n1588), .DIN1(n1496), .DIN2(n1057) );
    nnd2s1 U886 ( .Q(n1589), .DIN1(n810), .DIN2(n1588) );
    nnd2s1 U887 ( .Q(n1590), .DIN1(n939), .DIN2(n1589) );
    nnd2s1 U888 ( .Q(n1591), .DIN1(n1561), .DIN2(n1590) );
    nnd2s1 U889 ( .Q(n588), .DIN1(n1515), .DIN2(n1591) );
    hi1s1 U890 ( .Q(n1408), .DIN(N5045) );
    hi1s1 U891 ( .Q(n1273), .DIN(n979) );
    nnd2s1 U892 ( .Q(n1262), .DIN1(n961), .DIN2(N283) );
    nnd2s1 U893 ( .Q(n1265), .DIN1(n1569), .DIN2(N294) );
    nnd2s1 U894 ( .Q(n1264), .DIN1(n1566), .DIN2(N303) );
    nnd2s1 U895 ( .Q(n1269), .DIN1(N311), .DIN2(n727) );
    nnd2s1 U896 ( .Q(n1268), .DIN1(N317), .DIN2(n1567) );
    nnd2s1 U897 ( .Q(n1271), .DIN1(N322), .DIN2(n1568) );
    nnd2s1 U898 ( .Q(n1251), .DIN1(N150), .DIN2(n803) );
    nnd2s1 U899 ( .Q(n1250), .DIN1(n1566), .DIN2(N68) );
    nnd2s1 U900 ( .Q(n1255), .DIN1(n727), .DIN2(N58) );
    nnd2s1 U901 ( .Q(n1254), .DIN1(n1567), .DIN2(N50) );
    nnd2s1 U902 ( .Q(n1257), .DIN1(N159), .DIN2(n1568) );
    nnd2s1 U903 ( .Q(n1282), .DIN1(n1258), .DIN2(n1252) );
    nnd2s1 U904 ( .Q(n1281), .DIN1(n1272), .DIN2(n1266) );
    nnd2s1 U905 ( .Q(n567), .DIN1(n1284), .DIN2(n1283) );
    hi1s1 U906 ( .Q(n1405), .DIN(N5047) );
    nnd2s1 U907 ( .Q(n603), .DIN1(n655), .DIN2(n647) );
    nnd2s1 U908 ( .Q(n1082), .DIN1(n1313), .DIN2(n1592) );
    nnd2s1 U909 ( .Q(n1083), .DIN1(n1531), .DIN2(n1528) );
    hi1s1 U910 ( .Q(n1593), .DIN(n850) );
    nnd2s1 U911 ( .Q(n1302), .DIN1(n961), .DIN2(N294) );
    nnd2s1 U912 ( .Q(n1305), .DIN1(n1569), .DIN2(N303) );
    nnd2s1 U913 ( .Q(n1304), .DIN1(N311), .DIN2(n1566) );
    nnd2s1 U914 ( .Q(n1309), .DIN1(N317), .DIN2(n727) );
    nnd2s1 U915 ( .Q(n1308), .DIN1(N322), .DIN2(n1567) );
    nnd2s1 U916 ( .Q(n1311), .DIN1(N326), .DIN2(n1568) );
    nnd2s1 U917 ( .Q(n1291), .DIN1(N159), .DIN2(n803) );
    nnd2s1 U918 ( .Q(n1290), .DIN1(n1566), .DIN2(N77) );
    nnd2s1 U919 ( .Q(n1295), .DIN1(n727), .DIN2(N68) );
    nnd2s1 U920 ( .Q(n1294), .DIN1(n1567), .DIN2(N58) );
    nnd2s1 U921 ( .Q(n1297), .DIN1(n1568), .DIN2(N50) );
    nnd2s1 U922 ( .Q(n1316), .DIN1(n1298), .DIN2(n1292) );
    nnd2s1 U923 ( .Q(n1315), .DIN1(n1312), .DIN2(n1306) );
    nnd2s1 U924 ( .Q(n591), .DIN1(n1318), .DIN2(n1317) );
    nnd2s1 U925 ( .Q(n1582), .DIN1(n1561), .DIN2(n708) );
    nnd2s1 U926 ( .Q(n592), .DIN1(n1285), .DIN2(n1582) );
    hi1s1 U927 ( .Q(n1407), .DIN(N4815) );
    nnd2s1 U928 ( .Q(n1547), .DIN1(n1544), .DIN2(N350) );
    nnd2s1 U929 ( .Q(n1546), .DIN1(N5120), .DIN2(n1594) );
    nor2s1 U930 ( .Q(n1544), .DIN1(n886), .DIN2(N343) );
    hi1s1 U931 ( .Q(n1409), .DIN(N5192) );
    nnd2s1 U932 ( .Q(n1553), .DIN1(N1), .DIN2(n852) );
    nnd2s1 U933 ( .Q(n590), .DIN1(n1410), .DIN2(N1) );
    nnd2s1 U934 ( .Q(n598), .DIN1(n924), .DIN2(n922) );
    nnd2s1 U935 ( .Q(n1595), .DIN1(n1152), .DIN2(n1145) );
    nnd2s1 U936 ( .Q(n1596), .DIN1(n1166), .DIN2(n1159) );
    hi1s1 U937 ( .Q(n1597), .DIN(n855) );
    hi1s1 U938 ( .Q(n637), .DIN(n887) );
    nnd2s1 U939 ( .Q(n594), .DIN1(n1593), .DIN2(n939) );
    nor2s1 U940 ( .Q(n992), .DIN1(n884), .DIN2(n1430) );
    nnd2s1 U941 ( .Q(n1598), .DIN1(n1430), .DIN2(n884) );
    hi1s1 U942 ( .Q(n757), .DIN(n936) );
    nnd2s1 U943 ( .Q(n1041), .DIN1(n1038), .DIN2(n892) );
    nnd2s1 U944 ( .Q(n1040), .DIN1(n890), .DIN2(N274) );
    nnd2s1 U945 ( .Q(n1037), .DIN1(n1034), .DIN2(N107) );
    nnd2s1 U946 ( .Q(n1036), .DIN1(n609), .DIN2(n655) );
    nnd2s1 U947 ( .Q(n1599), .DIN1(N169), .DIN2(n909) );
    nnd2s1 U948 ( .Q(n1600), .DIN1(n1113), .DIN2(N179) );
    nnd2s1 U949 ( .Q(n978), .DIN1(n1600), .DIN2(n1599) );
    nnd2s1 U950 ( .Q(n1601), .DIN1(n1113), .DIN2(n871) );
    nnd2s1 U951 ( .Q(n1602), .DIN1(n909), .DIN2(n872) );
    nnd2s1 U952 ( .Q(n1603), .DIN1(n1602), .DIN2(n1601) );
    nnd2s1 U953 ( .Q(n1033), .DIN1(n1193), .DIN2(n1603) );
    nnd2s1 U954 ( .Q(n1604), .DIN1(n1045), .DIN2(n876) );
    nnd2s1 U955 ( .Q(n1605), .DIN1(n1042), .DIN2(N179) );
    nnd2s1 U956 ( .Q(n1606), .DIN1(n1605), .DIN2(n1604) );
    nnd2s1 U957 ( .Q(n1607), .DIN1(n1414), .DIN2(n923) );
    nnd2s1 U958 ( .Q(n1608), .DIN1(n1606), .DIN2(n798) );
    nnd2s1 U959 ( .Q(n933), .DIN1(n1608), .DIN2(n1607) );
    nnd2s1 U960 ( .Q(n1609), .DIN1(N169), .DIN2(n1463) );
    nnd2s1 U961 ( .Q(n1610), .DIN1(n1570), .DIN2(N179) );
    nnd2s1 U962 ( .Q(n945), .DIN1(n1610), .DIN2(n1609) );
    nnd2s1 U963 ( .Q(n1611), .DIN1(n1570), .DIN2(n871) );
    nnd2s1 U964 ( .Q(n1612), .DIN1(n1463), .DIN2(n872) );
    nnd2s1 U965 ( .Q(n1613), .DIN1(n1612), .DIN2(n1611) );
    nnd2s1 U966 ( .Q(n1049), .DIN1(n1122), .DIN2(n1613) );
    hi1s1 U967 ( .Q(n879), .DIN(n1048) );
    nnd2s1 U968 ( .Q(n1614), .DIN1(n1465), .DIN2(n879) );
    nor2s1 U969 ( .Q(n989), .DIN1(n879), .DIN2(n1465) );
    nnd2s1 U970 ( .Q(n1615), .DIN1(n1466), .DIN2(n695) );
    nor2s1 U971 ( .Q(n994), .DIN1(n695), .DIN2(n1466) );
    hi1s1 U972 ( .Q(n1534), .DIN(n993) );
    nnd2s1 U973 ( .Q(n1053), .DIN1(n1050), .DIN2(N68) );
    nnd2s1 U974 ( .Q(n1052), .DIN1(n609), .DIN2(n644) );
    nor2s1 U975 ( .Q(n997), .DIN1(n698), .DIN2(n1477) );
    nnd2s1 U976 ( .Q(n1616), .DIN1(n1477), .DIN2(n698) );
    hi1s1 U977 ( .Q(n1138), .DIN(n571) );
    nnd2s1 U978 ( .Q(n1617), .DIN1(n1479), .DIN2(n571) );
    nor2s1 U979 ( .Q(n999), .DIN1(n571), .DIN2(n1479) );
    nnd2s1 U980 ( .Q(n1618), .DIN1(N169), .DIN2(n1480) );
    nnd2s1 U981 ( .Q(n1619), .DIN1(n1564), .DIN2(N179) );
    nnd2s1 U982 ( .Q(n1574), .DIN1(n1619), .DIN2(n1618) );
    nnd2s1 U983 ( .Q(n1620), .DIN1(n1564), .DIN2(n871) );
    nnd2s1 U984 ( .Q(n1621), .DIN1(n1480), .DIN2(n872) );
    nnd2s1 U985 ( .Q(n1622), .DIN1(n1621), .DIN2(n1620) );
    nnd2s1 U986 ( .Q(n1054), .DIN1(n1563), .DIN2(n1622) );
    nor2s1 U987 ( .Q(n1002), .DIN1(n1486), .DIN2(n703) );
    nnd2s1 U988 ( .Q(n1623), .DIN1(n703), .DIN2(n1486) );
    nnd2s1 U989 ( .Q(n1624), .DIN1(n1487), .DIN2(n627) );
    nor2s1 U990 ( .Q(n1625), .DIN1(n627), .DIN2(n1487) );
    nnd2s1 U991 ( .Q(n1580), .DIN1(n1626), .DIN2(n1624) );
    nnd2s1 U992 ( .Q(n1627), .DIN1(n1595), .DIN2(n856) );
    nnd2s1 U993 ( .Q(n1628), .DIN1(N33), .DIN2(n1596) );
    nnd2s1 U994 ( .Q(n1629), .DIN1(n1628), .DIN2(n1627) );
    nnd2s1 U995 ( .Q(n1056), .DIN1(n1629), .DIN2(n866) );
    nnd2s1 U996 ( .Q(n1055), .DIN1(N50), .DIN2(N41) );
    nnd2s1 U997 ( .Q(n1004), .DIN1(n1489), .DIN2(n998) );
    nor2s1 U998 ( .Q(n1630), .DIN1(n998), .DIN2(n1489) );
    nnd2s1 U999 ( .Q(n1390), .DIN1(N5102), .DIN2(n1398) );
    nnd2s1 U1000 ( .Q(n1389), .DIN1(N5120), .DIN2(n1402) );
    nnd2s1 U1001 ( .Q(n1007), .DIN1(n1107), .DIN2(n1490) );
    nor2s1 U1002 ( .Q(n1631), .DIN1(n1490), .DIN2(n1107) );
    hi1s1 U1003 ( .Q(n759), .DIN(n1005) );
    nor2s1 U1004 ( .Q(n1632), .DIN1(n930), .DIN2(n1491) );
    nnd2s1 U1005 ( .Q(n1008), .DIN1(n1491), .DIN2(n930) );
    nor2s1 U1006 ( .Q(n1633), .DIN1(n1493), .DIN2(n1032) );
    nnd2s1 U1007 ( .Q(n1010), .DIN1(n1032), .DIN2(n1493) );
    hi1s1 U1008 ( .Q(n808), .DIN(n576) );
    nnd2s1 U1009 ( .Q(n1634), .DIN1(n759), .DIN2(n1635) );
    nnd2s1 U1010 ( .Q(n1636), .DIN1(n1005), .DIN2(n596) );
    nnd2s1 U1011 ( .Q(n1637), .DIN1(n1636), .DIN2(n1634) );
    nnd2s1 U1012 ( .Q(n1059), .DIN1(n759), .DIN2(n972) );
    nnd2s1 U1013 ( .Q(n1058), .DIN1(n1637), .DIN2(n595) );
    nnd2s1 U1014 ( .Q(n1638), .DIN1(n1494), .DIN2(n808) );
    nor2s1 U1015 ( .Q(n1013), .DIN1(n808), .DIN2(n1494) );
    hi1s1 U1016 ( .Q(n1496), .DIN(n1012) );
    nnd2s1 U1017 ( .Q(n1639), .DIN1(N97), .DIN2(n631) );
    nnd2s1 U1018 ( .Q(n1640), .DIN1(N87), .DIN2(n647) );
    nnd2s1 U1019 ( .Q(n1584), .DIN1(n1640), .DIN2(n1639) );
    nnd2s1 U1020 ( .Q(n1641), .DIN1(N116), .DIN2(n655) );
    nnd2s1 U1021 ( .Q(n1642), .DIN1(N107), .DIN2(n664) );
    nnd2s1 U1022 ( .Q(n1583), .DIN1(n1642), .DIN2(n1641) );
    nor2s1 U1023 ( .Q(n1643), .DIN1(n674), .DIN2(n1510) );
    nnd2s1 U1024 ( .Q(n1015), .DIN1(n1510), .DIN2(n674) );
    nnd2s1 U1025 ( .Q(n1644), .DIN1(N257), .DIN2(n671) );
    nnd2s1 U1026 ( .Q(n1645), .DIN1(N250), .DIN2(n680) );
    nnd2s1 U1027 ( .Q(n1587), .DIN1(n1645), .DIN2(n1644) );
    nnd2s1 U1028 ( .Q(n1646), .DIN1(N270), .DIN2(n684) );
    nnd2s1 U1029 ( .Q(n1647), .DIN1(N264), .DIN2(n836) );
    nnd2s1 U1030 ( .Q(n1586), .DIN1(n1647), .DIN2(n1646) );
    nnd2s1 U1031 ( .Q(n1061), .DIN1(n846), .DIN2(n631) );
    nnd2s1 U1032 ( .Q(n1060), .DIN1(n974), .DIN2(n986) );
    nnd2s1 U1033 ( .Q(n1321), .DIN1(N5045), .DIN2(n1401) );
    nnd2s1 U1034 ( .Q(n1320), .DIN1(N5078), .DIN2(n1408) );
    nnd2s1 U1035 ( .Q(n1276), .DIN1(N244), .DIN2(n657) );
    nnd2s1 U1036 ( .Q(n1275), .DIN1(N238), .DIN2(n666) );
    nnd2s1 U1037 ( .Q(n1279), .DIN1(N232), .DIN2(n633) );
    nnd2s1 U1038 ( .Q(n1278), .DIN1(N226), .DIN2(n649) );
    nnd2s1 U1039 ( .Q(n1648), .DIN1(n1274), .DIN2(n1649) );
    nor2s1 U1040 ( .Q(n1018), .DIN1(n1649), .DIN2(n1274) );
    nnd2s1 U1041 ( .Q(n1063), .DIN1(n1017), .DIN2(N45) );
    nnd2s1 U1042 ( .Q(n1062), .DIN1(n840), .DIN2(n851) );
    nnd2s1 U1043 ( .Q(n1066), .DIN1(n1064), .DIN2(n628) );
    nnd2s1 U1044 ( .Q(n1065), .DIN1(n788), .DIN2(n979) );
    nnd2s1 U1045 ( .Q(n1650), .DIN1(N58), .DIN2(n773) );
    nnd2s1 U1046 ( .Q(n1651), .DIN1(N50), .DIN2(n771) );
    nnd2s1 U1047 ( .Q(n1592), .DIN1(n1651), .DIN2(n1650) );
    nnd2s1 U1048 ( .Q(n1068), .DIN1(N45), .DIN2(n1081) );
    nnd2s1 U1049 ( .Q(n1067), .DIN1(n1593), .DIN2(n851) );
    nnd2s1 U1050 ( .Q(n1071), .DIN1(n1069), .DIN2(n628) );
    nnd2s1 U1051 ( .Q(n1070), .DIN1(n788), .DIN2(N1947) );
    nnd2s1 U1052 ( .Q(n1324), .DIN1(N4815), .DIN2(n1405) );
    nnd2s1 U1053 ( .Q(n1323), .DIN1(N5047), .DIN2(n1407) );
    nnd2s1 U1054 ( .Q(n1652), .DIN1(n1319), .DIN2(n1653) );
    nor2s1 U1055 ( .Q(n1021), .DIN1(n1653), .DIN2(n1319) );
    hi1s1 U1056 ( .Q(n1654), .DIN(n1020) );
    nnd2s1 U1057 ( .Q(n1025), .DIN1(N4944), .DIN2(n1399) );
    nnd2s1 U1058 ( .Q(n1024), .DIN1(N5121), .DIN2(n1404) );
    hi1s1 U1059 ( .Q(n1655), .DIN(n1023) );
    nnd2s1 U1060 ( .Q(n1656), .DIN1(n1543), .DIN2(n1545) );
    nor2s1 U1061 ( .Q(n1392), .DIN1(n1545), .DIN2(n1543) );
    nnd2s1 U1062 ( .Q(n1396), .DIN1(n1654), .DIN2(n1655) );
    nnd2s1 U1063 ( .Q(n1395), .DIN1(n1023), .DIN2(n1020) );
    nor2s1 U1064 ( .Q(n1657), .DIN1(n1391), .DIN2(n1394) );
    nnd2s1 U1065 ( .Q(n1026), .DIN1(n1394), .DIN2(n1391) );
    nnd2s1 U1066 ( .Q(n1075), .DIN1(n1072), .DIN2(n644) );
    nnd2s1 U1067 ( .Q(n1074), .DIN1(N68), .DIN2(n773) );
    nnd2s1 U1068 ( .Q(n1658), .DIN1(n946), .DIN2(n1548) );
    nor2s1 U1069 ( .Q(n1659), .DIN1(n1548), .DIN2(n946) );
    nnd2s1 U1070 ( .Q(n1550), .DIN1(n1660), .DIN2(n1658) );
    nor2s1 U1071 ( .Q(n1661), .DIN1(n949), .DIN2(n934) );
    nnd2s1 U1072 ( .Q(n1412), .DIN1(n934), .DIN2(n949) );
    nor2s1 U1073 ( .Q(n1662), .DIN1(n1549), .DIN2(n1411) );
    nnd2s1 U1074 ( .Q(n1663), .DIN1(n1411), .DIN2(n1549) );
    nnd2s1 U1075 ( .Q(n1552), .DIN1(n1663), .DIN2(n1664) );
    nnd2s1 U1076 ( .Q(n1665), .DIN1(N97), .DIN2(n655) );
    nnd2s1 U1077 ( .Q(n1666), .DIN1(N107), .DIN2(n647) );
    nnd2s1 U1078 ( .Q(n1555), .DIN1(n1666), .DIN2(n1665) );
    nnd2s1 U1079 ( .Q(n1029), .DIN1(n1508), .DIN2(n1081) );
    nor2s1 U1080 ( .Q(n1667), .DIN1(n1081), .DIN2(n1508) );
    nnd2s1 U1081 ( .Q(n1031), .DIN1(n1017), .DIN2(n1668) );
    nor2s1 U1082 ( .Q(n1669), .DIN1(n1017), .DIN2(n1668) );
    nnd2s1 U1083 ( .Q(n1080), .DIN1(n1077), .DIN2(n855) );
    nnd2s1 U1084 ( .Q(n1079), .DIN1(n1076), .DIN2(n1597) );
    hi1s1 U1085 ( .Q(n1009), .DIN(n1632) );
    hi1s1 U1086 ( .Q(n1499), .DIN(n1498) );
    hi1s1 U1087 ( .Q(n1167), .DIN(n1163) );
    hi1s1 U1088 ( .Q(n1393), .DIN(n1656) );
    hi1s1 U1089 ( .Q(n1027), .DIN(n1657) );
    hi1s1 U1090 ( .Q(n1660), .DIN(n1659) );
    hi1s1 U1091 ( .Q(n1215), .DIN(n1350) );
    hi1s1 U1092 ( .Q(n1207), .DIN(n1206) );
    hi1s1 U1093 ( .Q(n1189), .DIN(n1187) );
    hi1s1 U1094 ( .Q(n1664), .DIN(n1662) );
    hi1s1 U1095 ( .Q(n1421), .DIN(n863) );
    hi1s1 U1096 ( .Q(n1085), .DIN(n859) );
    hi1s1 U1097 ( .Q(n1516), .DIN(n1514) );
    hi1s1 U1098 ( .Q(n599), .DIN(n924) );
    hi1s1 U1099 ( .Q(n1467), .DIN(n1115) );
    hi1s1 U1100 ( .Q(n810), .DIN(n970) );
    hi1s1 U1101 ( .Q(n1001), .DIN(n1623) );
    hi1s1 U1102 ( .Q(n1626), .DIN(n1625) );
    hi1s1 U1103 ( .Q(n1003), .DIN(n1630) );
    hi1s1 U1104 ( .Q(n1107), .DIN(n912) );
    hi1s1 U1105 ( .Q(n1649), .DIN(n1277) );
    hi1s1 U1106 ( .Q(n793), .DIN(n976) );
    hi1s1 U1107 ( .Q(n1653), .DIN(n1322) );
    hi1s1 U1108 ( .Q(n1488), .DIN(n1573) );
    hi1s1 U1109 ( .Q(n748), .DIN(n937) );
    hi1s1 U1110 ( .Q(n1540), .DIN(n1388) );
    hi1s1 U1111 ( .Q(n1413), .DIN(n1661) );
    hi1s1 U1112 ( .Q(n1668), .DIN(n986) );
    hi1s1 U1113 ( .Q(n990), .DIN(n1614) );
    hi1s1 U1114 ( .Q(n991), .DIN(n1598) );
    hi1s1 U1115 ( .Q(n995), .DIN(n1615) );
    hi1s1 U1116 ( .Q(n938), .DIN(n1575) );
    hi1s1 U1117 ( .Q(n1011), .DIN(n1633) );
    hi1s1 U1118 ( .Q(n1014), .DIN(n1638) );
    hi1s1 U1119 ( .Q(n1019), .DIN(n1648) );
    hi1s1 U1120 ( .Q(n1260), .DIN(n802) );
    hi1s1 U1121 ( .Q(n1300), .DIN(n816) );
    hi1s1 U1122 ( .Q(n1006), .DIN(n1631) );
    hi1s1 U1123 ( .Q(n1635), .DIN(n596) );
    hi1s1 U1124 ( .Q(n1016), .DIN(n1643) );
    hi1s1 U1125 ( .Q(n1022), .DIN(n1652) );
    hi1s1 U1126 ( .Q(n996), .DIN(n1616) );
    hi1s1 U1127 ( .Q( tempn1000 ), .DIN(n1617) );
    hi1s1 U1128 ( .Q(n1177), .DIN(n726) );
    hi1s1 U1129 ( .Q(n1581), .DIN(n622) );
    hi1s1 U1130 ( .Q(n1542), .DIN(n1394) );
    hi1s1 U1131 ( .Q(n1594), .DIN(n1544) );
    hi1s1 U1132 ( .Q(n600), .DIN(n1414) );
    hi1s1 U1133 ( .Q(n1028), .DIN(n1667) );
    hi1s1 U1134 ( .Q(n1030), .DIN(n1669) );
  and4s1 troj51_0U1 ( .DIN1(n864), .DIN2(n644), .DIN3(troj51_0n1), .DIN4(troj51_0n2), .Q(        Trigger_en51_0) );
  and4s1 troj51_0U2 ( .DIN1(n1377), .DIN2(n1188), .DIN3(troj51_0n3), .DIN4(n1118), .Q(troj51_0n2) );
  nor2s1 troj51_0U3 ( .DIN1(n603), .DIN2(troj51_0n4), .Q(troj51_0n3) );
  i1s1 troj51_0U4 ( .DIN(n1042), .Q(troj51_0n4) );
  and3s1 troj51_0U5 ( .DIN1(n1513), .DIN2(n1506), .DIN3(n1554), .Q(troj51_0n1) );
    xor2s1 trojan51_0  (.DIN1(tempn1000), .DIN2(Trigger_en51_0), .Q(n1000) );

endmodule

