//****************************************************************
// TRIT-ASIC Generated Trojans.  The design generated below is for academic use only.
// Please cite the following if using the benchmark provided:
// J. Cruz, Y. Huang, P. Mishra, S. Bhunia, 
// "An Automated Configurable Trojan Insertion Framework for Dynamic Trust Benchmarks", DATE, 2018
//****************************************************************

module s38417( GND, VDD, CLK, RST, g1249, g1943, g2637, g3212, g3213, g3214, 
		g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, 
		g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, 
		g51, g563, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, 
		g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090, g4200, 
		g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, 
		g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
		g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
		g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
		g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
		g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
		g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
		g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
		g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275);

	input GND, VDD, CLK, RST, g1249, g1943, g2637, g3212, g3213, g3214, g3215,
         g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225,
         g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51,
         g563;

	output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275;

	wire n5361, n7281, n7280, n10033, n10032, g2962, n15168, g2934, n15169, n10081, 
		n10084, n7247, n10065, n5369, n10066, n14868, n14891, n15502, n14915, n7283, 
		n10082, n10083, n9956, n9955, n5370, n10034, n10089, n5304, n9972, n5591, 
		n5356, n9960, n5589, n5354, n9965, n5590, n9963, n5362, n9962, n9952, 
		n10070, n10068, n10072, n5366, n10071, n5353, n9958, n5357, n9957, n9951, 
		n10040, n10038, n10042, n5365, n10041, n9977, n5592, n9975, n5364, n9974, 
		n9954, n10012, n10011, n10014, n5368, n10013, n5355, n9970, n5363, n9969, 
		n9953, n9990, n9989, n9992, n5367, n9991, g2256, g1562, g868, g180, 
		n10051, n10062, n5372, n10061, n10060, n5371, n10059, n9967, n10085, n10086, 
		n10087, n5377, n10088, n10029, n10028, n5374, n10027, n10026, n5373, n10025, 
		n10001, n10007, n10006, n10005, n5378, n10004, g286, n10016, g536, n7441, 
		n7440, n5401, n5434, n7433, n7439, n5436, n7424, n7434, g284, n10017, 
		g534, n5358, n9861, n5662, n9862, n5642, g454, n10020, g531, n10030, 
		n5376, n5498, n5329, g452, n10021, g530, n5497, n5328, g450, n10022, 
		g529, n7286, n5496, n5327, g1139, n9999, g1216, n5493, n5324, g1137, 
		n10000, g1215, n7285, n5492, n5323, g2527, n10049, g2604, n7284, n5485, 
		n5316, g288, n10015, g537, n7445, n5413, n7446, n5435, n7442, n7444, 
		n5442, n7435, n7443, g282, n10018, g533, n5499, n5330, g280, n10019, 
		g532, n9859, n5661, n9860, n5641, n10031, n5678, n7397, n7398, n9978, 
		n5604, n7390, n7393, n10023, n5632, n5381, n7631, n5552, n5342, n7635, 
		n9837, n5660, n7456, n5424, g558, n7272, n9884, n5718, n9885, n5587, 
		n9985, n5588, n7313, n7314, n10024, n5673, n9839, n5634, n7627, n5553, 
		n5343, n7622, n7341, n7342, n9835, n5658, n7462, n5425, g549, n5383, 
		n5307, n5384, n7379, n7380, n7473, n7474, n9841, n5630, n9836, n5659, 
		n7458, n5426, g543, g544, n15417, n9924, n5579, n9927, n5585, n9983, 
		n5569, n7651, n9848, n5736, n9849, n5692, n7649, n9850, n5734, n9851, 
		n5690, n7650, n9852, n5733, n9853, n5689, n7469, n7470, n9840, n5631, 
		n7655, n9846, n5732, n9847, n5688, n7657, n5527, n9856, n5713, n7654, 
		n9843, n5731, n9844, n5687, n7471, n7472, n9842, n5629, n7332, n7334, 
		n7652, n5529, n9858, n5716, n7656, n5528, n9857, n5715, n7621, n5526, 
		n9845, n5714, n7653, n9854, n5735, n9855, n5691, g471, g568, n15652, 
		g468, g566, g567, g465, g574, n9834, g528, g535, g542, g376, 
		g382, n15068, g373, g380, n15069, g361, g367, n15071, g358, g365, 
		n15073, g391, g397, n15064, g388, g395, n15065, g387, g394, g357, 
		g364, g372, g379, g346, g352, n15066, g343, g350, n15067, g342, 
		g349, g461, g572, n15638, g458, g570, g571, g455, g564, n9838, 
		g513, g523, g524, n15426, n5394, g975, n9993, g1223, n7437, n5412, 
		n7438, n5433, n7431, n7436, n5441, n7423, n7432, g973, n9994, g1222, 
		n7430, n7429, n5400, n5432, n7421, n7428, n5440, n7412, n7422, g971, 
		n9995, g1220, n5306, n9827, n5657, n9828, n5640, g969, n9996, g1219, 
		n5495, n5326, g967, n9997, g1218, n9825, n5656, n9826, n5639, g1141, 
		n9998, g1217, n10008, n5375, n5494, n5325, n9973, n5603, n7387, n7389, 
		n10002, n5670, n7630, n9808, n5633, n7584, n5332, n7634, n5524, n9806, 
		n5655, n7454, n5421, g1244, n7640, n5313, n9950, n5717, n7583, n10009, 
		n5677, n7395, n7396, n7339, n7340, n10003, n5671, n7626, n9809, n5672, 
		n5333, n7620, n5525, n9804, n5653, n7461, n5422, g1235, n9906, n5582, 
		n5308, n5309, n7378, n7377, n7468, n9811, n5664, n7467, n9805, n5654, 
		n7457, n5423, g1229, n14876, n9923, n9916, n5578, n7666, n5311, n7333, 
		n7643, n5397, n9817, n5712, n7648, n5537, n9822, n5705, n7645, n9813, 
		n5728, n9814, n5685, n7464, n9810, n5665, n7463, n7642, n5540, n9820, 
		n5707, n7646, n5536, n9816, n5706, n7466, n9812, n5663, n7465, n7331, 
		n7644, n5538, n9824, n5711, n7647, n5539, n9823, n5710, n7618, n5535, 
		n9815, n5709, n7619, n5541, n9821, n5708, n7641, n9818, n5729, n9819, 
		n5686, g1158, g1254, n15647, g1155, g1252, g1253, g1152, g1260, n9803, 
		g1214, g1221, g1228, g985, n5568, g1041, g1029, g1036, g1063, g1069, 
		n15058, g1067, n15059, g1071, g1059, g1066, g1048, g1054, n15061, g1052, 
		n15063, g1056, g1044, g1051, g1078, g1084, n15054, g1082, n15055, g1085, 
		g1074, g1081, g1033, g1039, n15056, g1037, n15057, g1148, g1258, n15631, 
		g1145, g1256, g1257, g1142, g1250, n9807, g1199, g1209, g1210, g1831, 
		n10080, g1909, n5488, n5319, g2363, n10043, g2611, n7414, n5410, n7415, 
		n5428, n7407, n7413, n5438, n7402, n7408, g2361, n10044, g2610, n7406, 
		n7405, n5398, n5427, n7400, n7404, n5437, n7399, n7401, g2359, n10045, 
		g2608, n5359, n9909, n5647, n9910, n5636, g2357, n10046, g2607, n7287, 
		n5487, n5318, g2355, n10047, g2606, n5305, n9907, n5646, n9908, n5635, 
		g2529, n10048, g2605, n10063, n5379, n5486, n5317, g2525, n10050, g2603, 
		n5484, n5315, n10064, n5675, n7388, n7391, n7382, n7381, n7674, n5521, 
		n9896, n5694, n7670, n5395, n9897, n5698, n7672, n9901, n5721, n9902, 
		n5680, n7668, n9898, n5720, n9899, n5679, n7572, n7571, n9892, n5611, 
		n7675, n5523, n9904, n5696, n7669, n5522, n9900, n5695, n7676, n5519, 
		n9903, n5693, n7673, n5331, n5547, n7667, n9895, n5738, n5542, n7574, 
		n7573, n9894, n5609, n9880, n5644, n7453, n5417, g2617, n14885, n7327, 
		n7328, n7576, n7575, n9893, n5610, n7671, n5520, n9905, n5697, g2546, 
		g2642, n15635, g2543, g2640, g2641, g2540, g2648, n9878, g2602, g2609, 
		g2616, g2451, g2457, n15038, g2448, g2455, n15039, g2436, g2442, n15041, 
		g2433, g2440, n15043, g2466, g2472, n15034, g2463, g2470, n15035, g2462, 
		g2469, g2432, g2439, g2447, g2454, g2421, g2427, n15036, g2418, g2425, 
		n15037, g2417, g2424, g2536, g2646, n15627, g2533, g2644, g2645, g2530, 
		g2638, n9882, g2587, g2597, g2598, n14920, n9961, n5601, n7383, n7384, 
		n10052, n5612, n5380, n7628, n5548, n5338, n7617, n9881, n5645, n7451, 
		n5415, g2632, n9984, n5737, n9931, n5586, n5314, n7310, n7309, n10058, 
		n5666, n9889, n5667, n7624, n5549, n5339, n7677, n7336, n7335, n9879, 
		n5643, n7459, n5416, g2623, n9890, n5575, n5386, n9891, n5576, g1669, 
		n10073, g1917, n7426, n5411, n7427, n5430, n7419, n7425, n5439, n7411, 
		n7420, g1667, n10074, g1916, n7418, n7417, n5399, n5429, n7409, n7416, 
		n5431, n7403, n7410, g1665, n10075, g1914, n9796, n5652, n9797, n5638, 
		g1663, n10076, g1913, n5491, n5322, g1661, n10077, g1912, n5360, n9794, 
		n5651, n9795, n5637, g1835, n10078, g1911, n5490, n5321, g1833, n10079, 
		g1910, n5489, n5320, n9968, n5602, n7385, n7386, n5562, n9792, n5620, 
		n7629, n5550, n5340, n7633, n9929, n5650, n7452, n5418, g1938, n5500, 
		n9932, n5580, n5389, n7312, n7311, n9987, n5676, n7392, n7394, n7338, 
		n7337, n9986, n5668, n9793, n5669, n7625, n5551, n5341, n7623, n9926, 
		n5648, n7460, n5419, g1929, n5385, n5310, n9981, n5581, n7376, n7375, 
		n7582, n7581, n9935, n5618, n7681, n5396, n9939, n5704, n7679, n9943, 
		n5725, n9944, n5683, n7578, n7577, n9933, n5619, n7686, n5532, n9949, 
		n5702, n7678, n5531, n9947, n5701, n7683, n9940, n5726, n9941, n5684, 
		n7680, n5534, n9942, n5700, n7685, n9945, n5724, n9946, n5682, n7687, 
		n5533, n9948, n5699, n7684, n9937, n5723, n9938, n5681, n7580, n7579, 
		n9934, n5617, n7329, n7330, n7682, n5530, n9936, n5703, g1852, g1948, 
		n15642, g1849, g1946, g1947, g1846, g1954, n9925, g1908, g1915, g1922, 
		g1757, g1763, n15048, g1754, g1761, n15049, g1742, g1748, n15051, g1739, 
		g1746, n15053, g1772, g1778, n15044, g1769, g1776, n15045, g1768, g1775, 
		g1738, g1745, g1753, g1760, g1727, g1733, n15046, g1724, g1731, n15047, 
		g1723, g1730, g1842, g1952, n15629, g1839, g1950, g1951, g1836, g1944, 
		n9930, g1893, g1903, g1904, g1679, n9966, n5674, n7632, n9928, n5649, 
		n7455, n5420, g1923, n14880, n9922, n5387, n9915, n5577, n5388, n9913, 
		n9982, n5583, n9912, n5584, n5312, n9888, n9887, n10055, n5483, n9979, 
		n9980, n5382, n10054, n5352, n15211, g3194, n10057, n10053, n15214, g3198, 
		n15217, n15213, n10056, n5739, g3125, n15212, n5567, g2878, g2365, DFF_1503_D, 
		n9863, n9872, g2873, g977, DFF_803_D, n9865, n9866, g2857, g290, DFF_453_D, 
		n9868, n9869, g2877, g1671, DFF_1153_D, n9864, n9914, n5406, n9798, n5623, 
		n9799, n5597, n5407, n9800, n5624, n9801, n5598, n5556, n5346, n7663, 
		n15150, n5509, n7359, n7360, n5511, n7361, n7362, n5510, n7365, n7366, 
		n5512, n5555, n5345, n7662, n9988, n5621, n7449, n5392, n5564, n9802, 
		n5727, n7638, n7363, n7364, n9867, n5572, n7534, n5458, n5408, n9829, 
		n5627, n9830, n5599, n5409, n9831, n5628, n9832, n5600, n5558, n5348, 
		n7665, n15423, n9976, n5518, n7549, n7551, n7560, n7562, n7564, n7566, 
		n7557, n7553, n7555, n7568, n7318, n7548, n7550, n7559, n7561, n7563, 
		n7565, n7556, n7552, n7554, n7567, n5336, n5463, n5466, n5472, n5469, 
		n5470, n5467, n5465, n10036, n5626, n5464, n5471, n5545, n9971, n5517, 
		n7525, n7527, n7536, n7538, n7540, n7542, n7533, n7529, n7531, n7544, 
		n7317, n7524, n7526, n7535, n7537, n7539, n7541, n7532, n7528, n7530, 
		n7543, n5335, n5453, n5456, n5462, n5459, n5460, n5457, n5455, n10035, 
		n5622, n5454, n5461, n7523, n7546, n7545, n5544, g3061, g3060, g3059, 
		g3058, g3057, g3056, g3055, g3053, g3052, n5513, n7367, n7368, n5515, 
		n7369, n7370, n5514, n7373, n7374, n5516, n5557, n5347, n7664, n10010, 
		n5625, n7450, n5393, n5565, n9833, n5730, n7639, n7371, n7372, n9870, 
		n5573, n7558, n5468, n7547, n7570, n7569, g3050, g3048, g3044, g3046, 
		g3045, g3043, g3049, g3051, g3047, n5402, n9873, n5607, n9874, n5593, 
		n5403, n9875, n5608, n9876, n5594, n5561, n5351, n7659, g2581, n5501, 
		n7343, n7344, n5503, n7345, n7346, n5502, n7349, n7350, n5504, n5560, 
		n5350, n7658, n10037, n5605, n7447, n5390, n5566, n9877, n5719, n7636, 
		n7347, n7348, n9871, n5570, n7486, n5448, n5404, n9917, n5615, n9918, 
		n5595, n5405, n9919, n5616, n9920, n5596, n5559, n5349, n7661, n9911, 
		n5571, n7510, n5478, n15018, n9964, n7501, n7503, n7512, n7514, n7516, 
		n7518, n7509, n7505, n7507, n7520, n7316, n7500, n7502, n7511, n7513, 
		n7515, n7517, n7508, n7504, n7506, n7519, n5337, n5473, n5476, n5482, 
		n5479, n5480, n5477, n5475, n10069, n5614, n5474, n5481, n5546, g3068, 
		g3066, n9959, n5574, n7477, n7479, n7488, n7490, n7492, n7494, n7485, 
		n7481, n7483, n7496, n7315, n7476, n7478, n7487, n7489, n7491, n7493, 
		n7484, n7480, n7482, n7495, n5334, n5443, n5446, n5452, n5450, n5449, 
		n5447, n5445, n10039, n5606, n5444, n5451, n7475, n7498, n7497, n5543, 
		g3078, g3076, g3077, g2997, g2990, g3075, g3074, g3071, g3073, g3072, 
		n15173, n5505, n7351, n7352, n5507, n7353, n7354, n5506, n7357, n7358, 
		n5508, n5554, n5344, n7660, n5563, n9921, n5722, n7637, n10067, n5613, 
		n7448, n5391, n7499, n7522, n7521, g3064, g3062, g3065, g3063, g3069, 
		g3070, g3083, g3067, n15172, n7355, n7356, n9883, n15165, n5414, n15162, 
		g3128, n9886, n7602, n7597, n7604, n7608, n7600, n7606, n7325, n7715, 
		n7735, n7740, n7323, n7736, n7734, n7739, n7737, n7713, n7732, n7324, 
		n7714, n7733, n7738, g2950, n7613, n7612, n7616, n7615, n7610, n7609, 
		n7614, n7322, n7611, g354, g384, g369, g398, g2429, g2459, g2444, 
		g2473, g1735, g1765, g1750, g1779, n7745, n7744, n7742, n7741, n7743, 
		n7725, n7731, n7730, n7594, n7242, g1060, g1045, g1075, g1030, n7278, 
		n7276, n7275, n7277, n7729, n7728, n7726, n7727, n7288, n7294, n7289, 
		n7723, n7724, n7255, n7587, n7291, n7603, n7595, n7601, n7596, n7607, 
		n7599, n7605, n7598, n7709, n7307, n7710, n7308, n7712, n7306, n7711, 
		n7305, n7321, n7588, n7722, n7269, n7241, n7270, n7292, n7293, n7261, 
		n7221, n7704, n7700, n7701, n7703, n7258, n7260, n7257, n7259, n7716, 
		n7589, n7326, n7290, n7696, n7699, n7697, n7702, n7304, n7698, n7593, 
		n7243, n7233, n7223, n7222, n7590, n7591, n7254, g1186, g1880, n7303, 
		n7268, n7244, n7273, n7274, n7299, n7302, n7301, g3080, n7320, n7707, 
		n7708, n7706, n7705, n7585, n7592, n7720, n7717, n7718, n7719, n7232, 
		n7240, n7252, n7251, n7586, n7234, g499, g2574, n7226, n7224, n7225, 
		n7227, n7279, n7721, n7249, n7319, n7235, n7250, n7246, n7282, n7248, 
		n7267, n7245, n7271, n7300, n7690, n7296, n7689, n7295, n7688, n7691, 
		n7265, n7298, n7297, n7239, n7237, n7236, n7238, n7692, n7695, n7694, 
		n7693, n7262, n7229, n7230, n7231, n7264, n7266, n7263, n7782, n7256, 
		n7780, n7784, n7228, n7775, n5740, n5742, n5746, n5750, n5743, n5744, 
		n5749, n5747, n5748, n5753, n5754, n5745, n5752, n5751, n5741, n5755, 
		n5757, n5756, n5758, n5762, n5760, n5759, n5761, n5763, n5764, n5765, 
		n89, n5766, n88, n5769, n87, n5770, n86, n5771, n85, n5772, 
		n84, n5773, n83, n5774, n82, n5775, n81, n5776, n80, n5777, 
		n79, n5778, n78, n5779, n77, n5780, n76, n5781, n75, n5782, 
		n74, n5783, n73, n5784, n72, n5785, n5768, n5767, n69, n67, 
		n66, n65, n64, n63, n62, n61, n60, n57, n56, n55, 
		n54, n5303, n5302, n5799, n5300, n53, n5299, n5805, n5297, n5296, 
		n5810, n5294, n5293, n5815, n5291, n5290, n5289, n5288, n5287, n5286, 
		n5285, n5284, n5283, n5282, n5281, n5280, n5279, n5278, n5277, n5276, 
		n5275, n5274, n5854, n5273, n5856, n5272, n5271, n5859, n5270, n5862, 
		n5861, n5269, n5860, n5866, n5268, n5870, n5869, n5873, n5868, n5864, 
		n5863, n5865, n5872, n5267, n5875, n5877, n5266, n5879, n5265, n5880, 
		n5878, n5264, n5882, n5263, n5883, n5881, n5262, n5885, n5884, n5261, 
		n5876, n5887, n5260, n5259, n5886, n5258, n5257, n5256, n5255, n5897, 
		n5254, n5901, n5253, n5898, n5909, n5911, n5908, n5915, n5918, n5917, 
		n5916, n5923, n5922, n5921, n5914, n5929, n5928, n5927, n5913, n5912, 
		n5252, n5251, n5250, n5936, n5249, n5891, n5248, n5939, n5301, n5910, 
		n5247, n5941, n5803, n5895, n5246, n5946, n5245, n5947, n5244, n5243, 
		n5948, n5242, n5949, n5241, n5240, n5950, n5239, n5951, n5238, n5237, 
		n5952, n5236, n5953, n5235, n5234, n5954, n5233, n5955, n5232, n5231, 
		n5956, n5230, n5957, n5229, n5228, n5958, n5227, n5959, n5226, n5225, 
		n5224, n5223, n5222, n5962, n5221, n5963, n5220, n5219, n5899, n5964, 
		n5896, n5890, n5218, n5902, n5966, n5900, n5892, n5217, n5905, n5903, 
		n5894, n5967, n5216, n5969, n5215, n5970, n5214, n5973, n5972, n5971, 
		n5213, n5975, n5212, n5976, n5974, n5211, n5978, n5210, n5977, n5802, 
		n5933, n5209, n5979, n5800, n5208, n5893, n5801, n5980, n5965, n5207, 
		n5968, n5206, n5937, n5205, n5985, n5786, n5204, n5203, n5202, n5988, 
		n5991, n5201, n5200, n52, n5199, n5997, n5995, n5998, n6000, n6003, 
		n5198, n5197, n5196, n6007, n6006, n6008, n6002, n6011, n6013, n6012, 
		n6010, n6020, n6024, n6028, n6019, n6035, n6036, n6037, n6034, n6009, 
		n6038, n6001, n6040, n6031, n6039, n6014, n6046, n6044, n6049, n6051, 
		n6052, n6050, n6048, n6055, n6043, n6058, n6060, n6027, n6059, n6016, 
		n6026, n6029, n6057, n6017, n6062, n6056, n6033, n6047, n6063, n6022, 
		n6064, n5195, n5194, n5193, n6065, n6005, n6068, n6067, n5192, n5191, 
		n5990, n5989, n5190, n6070, n6004, n6073, n6072, n5993, n58, n5992, 
		n5189, n6078, n5188, n6081, n5187, n6075, n6023, n5186, n6086, n5185, 
		n6087, n5184, n6085, n6090, n6025, n6088, n5183, n6092, n5182, n6093, 
		n5181, n6091, n6089, n6084, n6042, n5180, n6095, n6077, n6076, n5179, 
		n6097, n6080, n6079, n5178, n6083, n6094, n6099, n6021, n6102, n6100, 
		n6103, n6030, n6018, n6054, n6032, n6061, n6104, n6041, n6105, n6015, 
		n6053, n6106, n6082, n5177, n5176, n5175, n5174, n6111, n5173, n5172, 
		n5171, n6114, n5170, n5169, n6109, n5168, n6116, n6110, n5167, n6112, 
		n5166, n5165, n5164, n5163, n5162, n5161, n6117, n5160, n5987, n5986, 
		n5159, n6045, n5158, n5157, n5156, n5155, n5154, n5153, n5152, n5151, 
		n5150, n6120, n6126, n6125, n6124, n6123, n6132, n6119, n6137, n6136, 
		n6135, n6134, n6143, n6142, n6141, n5149, n6148, n6147, n5148, n5147, 
		n5146, n6155, n6154, n5145, n6160, n6159, n5144, n6162, n6156, n6153, 
		n6165, n5143, n6170, n5142, n6173, n5141, n6176, n6175, n6172, n6177, 
		n6169, n6180, n6179, n6183, n5140, n5139, n6192, n5138, n6190, n6194, 
		n6196, n6197, n6200, n6202, n6205, n6201, n6199, n6181, n5137, n5136, 
		n6209, n5135, n6208, n6210, n6212, n6213, n6216, n6217, n6218, n6215, 
		n6221, n6223, n6220, n6222, n6186, n6229, n6230, n6228, n6225, n5134, 
		n5133, n6242, n5132, n6241, n6244, n5131, n6248, n6247, n5130, n6251, 
		n6250, n5129, n6252, n6249, n6255, n6246, n6258, n5128, n5127, n5126, 
		n6260, n6115, n6262, n6256, n6266, n6253, n6254, n6267, n6269, n6268, 
		n6263, n6270, n6261, n5125, n5124, n5123, n6271, n6257, n6275, n6274, 
		n6273, n6259, n6280, n6272, n5122, n6284, n6283, n5121, n6287, n6286, 
		n5120, n6288, n6285, n5119, n5118, n5117, n6292, n6294, n6296, n6291, 
		n6293, n5116, n6188, n6157, n6152, n5115, n6191, n6149, n6158, n5114, 
		n6193, n6164, n6161, n6300, n6302, n6304, n6282, n6290, n6306, n6295, 
		n6307, n6168, n6303, n6309, n6298, n6305, n6308, n6299, n6312, n6289, 
		n6151, n6107, n6313, n6297, n6314, n6301, n5113, n5112, n6315, n6317, 
		n5111, n6320, n6318, n6319, n5110, n6322, n5109, n6321, n5108, n6325, 
		n6324, n6323, n5107, n6327, n5106, n6326, n6329, n6328, n5105, n6330, 
		n5104, n6333, n6332, n6331, n5103, n6316, n6335, n6334, n5102, n6338, 
		n5101, n5100, n6340, n6346, n6351, n6353, n51, n5099, n5098, n5097, 
		n6357, n6361, n6362, n6352, n6364, n6367, n6366, n5096, n5095, n5094, 
		n6370, n6371, n6372, n6373, n6374, n5093, n5092, n5091, n6376, n6377, 
		n6378, n6365, n6380, n5090, n5089, n5088, n6382, n6383, n6385, n6379, 
		n6386, n5087, n5086, n5085, n6389, n6390, n6391, n6387, n5084, n6395, 
		n5083, n5082, n6396, n6397, n6398, n6394, n6393, n6399, n5081, n5080, 
		n5079, n6403, n6404, n6406, n6359, n6405, n6401, n6409, n5078, n5077, 
		n5076, n6411, n6350, n6360, n6412, n6413, n6414, n5075, n6341, n6339, 
		n5074, n6342, n6343, n5073, n6345, n6416, n6417, n6418, n6349, n6347, 
		n6422, n6424, n6423, n6219, n6426, n6171, n6174, n6425, n6185, n6239, 
		n6431, n6430, n6428, n6432, n6227, n6237, n6236, n6238, n6429, n6427, 
		n6232, n6224, n6437, n6436, n6434, n6235, n6438, n6226, n6233, n6234, 
		n6435, n6433, n6231, n6113, n6182, n6184, n6421, n6206, n6441, n6420, 
		n6384, n6408, n6419, n6195, n6167, n6443, n6163, n6178, n6166, n6445, 
		n6449, n6450, n6448, n6453, n6447, n6456, n6446, n6204, n6214, n6440, 
		n6460, n6459, n6463, n6458, n6466, n6444, n6472, n6473, n6471, n6475, 
		n6470, n6477, n6469, n6481, n6482, n6480, n6485, n6487, n6474, n6457, 
		n6478, n6486, n6489, n6476, n6488, n6483, n6484, n6492, n6491, n6479, 
		n6496, n6490, n6122, n6498, n6442, n6499, n6138, n6363, n6500, n6356, 
		n6139, n6407, n6501, n6410, n6133, n6502, n6497, n6146, n6504, n6381, 
		n6503, n6128, n6439, n6505, n6415, n6129, n6368, n6506, n6369, n6144, 
		n6507, n6375, n6145, n6508, n6388, n6392, n6354, n6243, n6211, n6140, 
		n6400, n6509, n6402, n6127, n6510, n6344, n5072, n5071, n6515, n5070, 
		n6513, n6276, n6521, n5828, n5826, n5824, n5821, n6520, n5836, n5834, 
		n5830, n6518, n5069, n6523, n5068, n5067, n5066, n6526, n5065, n5064, 
		n5063, n6511, n6512, n5062, n6462, n6514, n6516, n5061, n6461, n6517, 
		n6528, n5832, n6519, n5060, n5059, n6451, n5058, n6531, n6310, n6348, 
		n6536, n6527, n6452, n5057, n5056, n6454, n5055, n6537, n6311, n6358, 
		n6538, n6524, n6277, n6455, n5054, n6495, n5053, n5052, n6539, n5051, 
		n6493, n5050, n5049, n6540, n5048, n5047, n5046, n6541, n5045, n5044, 
		n5043, n6542, n5042, n6494, n5041, n5040, n6543, n5039, n5038, n5037, 
		n6544, n5036, n5035, n6467, n5034, n6468, n6525, n5033, n6530, n6336, 
		n5032, n6464, n6532, n6533, n5031, n6465, n6534, n6535, n6522, n5030, 
		n5029, n5028, n5027, n6553, n5026, n6557, n5025, n6554, n6565, n6567, 
		n6564, n6571, n6574, n6573, n6572, n6579, n6578, n6577, n6570, n6585, 
		n6584, n6583, n6569, n6568, n5024, n5023, n5022, n6591, n5021, n6547, 
		n5020, n6594, n5298, n6566, n5019, n6596, n5809, n6551, n5018, n6601, 
		n5017, n6602, n5016, n5015, n6603, n5014, n6604, n5013, n5012, n6605, 
		n5011, n6606, n5010, n5009, n6607, n5008, n6608, n5007, n5006, n6609, 
		n5005, n6610, n5004, n5003, n6611, n5002, n6612, n5001, n5000, n6613, 
		n50, n4999, n6615, n4998, n4997, n4996, n4995, n4994, n6618, n4993, 
		n6619, n4992, n4991, n6555, n6620, n6552, n6546, n4990, n6558, n6622, 
		n6556, n6548, n4989, n6561, n6559, n6550, n6623, n4988, n6625, n4987, 
		n6626, n4986, n6629, n6628, n6627, n4985, n6631, n4984, n6632, n6630, 
		n4983, n6634, n4982, n6633, n5808, n6635, n4981, n6636, n5806, n4980, 
		n6549, n5807, n6637, n6621, n4979, n6624, n4978, n6592, n4977, n4976, 
		n4975, n4974, n4973, n4972, n6643, n6646, n4971, n4970, n4969, n6651, 
		n6650, n6652, n6654, n4968, n4967, n4966, n6660, n6659, n6661, n6664, 
		n6657, n6670, n6668, n6676, n6677, n6666, n6685, n6687, n6688, n6663, 
		n6658, n6655, n6691, n6681, n6690, n6665, n6697, n6695, n6700, n6702, 
		n6703, n6701, n6699, n6669, n6694, n6708, n6678, n6711, n6710, n6673, 
		n6706, n6709, n6679, n6707, n6682, n6698, n6713, n6674, n6714, n4965, 
		n4964, n4963, n6715, n6656, n6718, n6717, n4962, n4961, n6645, n6644, 
		n4960, n6720, n6689, n6723, n6722, n6648, n6647, n4959, n6728, n4958, 
		n6731, n4957, n6725, n6675, n4956, n6736, n4955, n6737, n4954, n6735, 
		n6683, n6686, n6738, n4953, n6741, n4952, n6742, n4951, n6740, n6739, 
		n6734, n6693, n4950, n6744, n6727, n6726, n4949, n6745, n6730, n6729, 
		n4948, n6733, n6743, n6746, n6667, n6749, n6747, n6750, n6680, n6671, 
		n6705, n6672, n6712, n6751, n6692, n6752, n6684, n6704, n6753, n6732, 
		n6640, n6756, n6595, n6649, n6599, n6754, n6757, n4947, n4946, n4945, 
		n4944, n4943, n6764, n4942, n4941, n4940, n6768, n4939, n4938, n6761, 
		n4937, n6770, n6763, n4936, n6766, n4935, n4934, n4933, n4932, n4931, 
		n4930, n4929, n6642, n6641, n4928, n6696, n4927, n4926, n4925, n4924, 
		n4923, n4922, n4921, n4920, n4919, n6150, n6772, n4918, n4917, n4916, 
		n6779, n6778, n4915, n6784, n6783, n4914, n6787, n6780, n6777, n6790, 
		n4913, n6795, n4912, n6798, n4911, n6801, n6800, n6797, n6802, n6794, 
		n6805, n6804, n6808, n4910, n4909, n6817, n4908, n6815, n6819, n6821, 
		n6822, n6825, n6827, n6830, n6826, n6824, n6806, n4907, n4906, n6834, 
		n4905, n6833, n6835, n6837, n6838, n6842, n6843, n6844, n6840, n6846, 
		n6848, n6811, n6853, n6854, n6852, n6849, n4904, n4903, n6866, n4902, 
		n6865, n6868, n4901, n6872, n6871, n4900, n6875, n6874, n49, n4899, 
		n6877, n6873, n6880, n6870, n6883, n4898, n4897, n4896, n6885, n6887, 
		n6881, n6889, n6878, n6879, n6890, n6892, n6769, n6891, n6894, n6895, 
		n6886, n4895, n4894, n4893, n6896, n6884, n6898, n6893, n6882, n6901, 
		n6900, n6899, n6897, n4892, n6908, n6907, n4891, n6911, n6910, n4890, 
		n6912, n6909, n4889, n4888, n4887, n6916, n6918, n6920, n6915, n6917, 
		n4886, n6813, n6781, n6776, n4885, n6816, n6785, n6782, n4884, n6818, 
		n6789, n6786, n6924, n6926, n6928, n6906, n6914, n6930, n6919, n6931, 
		n6793, n6927, n6933, n6922, n6929, n6932, n6923, n6936, n6913, n6775, 
		n6759, n6937, n6921, n6938, n6925, n4883, n4882, n6940, n6942, n4881, 
		n6945, n6944, n6943, n4880, n6947, n4879, n6946, n4878, n6950, n6949, 
		n6948, n4877, n6952, n4876, n6951, n6953, n4875, n6955, n6954, n6957, 
		n4874, n6958, n6956, n4873, n6941, n6960, n6959, n4872, n4871, n4870, 
		n6964, n6970, n6975, n6978, n4869, n4868, n4867, n6982, n6983, n6986, 
		n6984, n6977, n6990, n6993, n6992, n4866, n4865, n4864, n6998, n6999, 
		n7000, n7001, n7002, n4863, n4862, n4861, n7004, n7005, n7006, n6991, 
		n7008, n4860, n4859, n4858, n7011, n7012, n7013, n7007, n7014, n4857, 
		n4856, n4855, n7018, n7019, n7020, n7015, n4854, n4853, n4852, n7027, 
		n7028, n7030, n7025, n7031, n4851, n4850, n4849, n7036, n7037, n7039, 
		n6987, n7038, n7023, n7033, n7042, n4848, n4847, n4846, n7045, n6974, 
		n7046, n7047, n7048, n4845, n6965, n6963, n4844, n6966, n6967, n4843, 
		n6969, n7051, n7052, n7053, n6973, n6971, n7057, n7059, n7058, n6845, 
		n7061, n6796, n6799, n7060, n6810, n6863, n7066, n7065, n7063, n6855, 
		n6857, n7064, n7067, n6850, n6859, n7062, n6858, n6847, n7071, n7070, 
		n7068, n6860, n6856, n6862, n6861, n7069, n6851, n7072, n6767, n6807, 
		n7056, n6831, n7074, n6869, n7055, n6985, n7041, n7054, n6820, n6792, 
		n7077, n6788, n6803, n6791, n7079, n7083, n7084, n7082, n7087, n7081, 
		n7090, n7080, n6829, n6841, n7073, n7094, n7093, n7097, n7092, n7100, 
		n7078, n7106, n7107, n7105, n7109, n7104, n7111, n7103, n7115, n7116, 
		n7114, n7120, n7122, n7108, n7091, n7112, n7121, n7124, n7110, n7123, 
		n7117, n7119, n7127, n7126, n7113, n7132, n7125, n7076, n7134, n7022, 
		n6980, n6867, n6968, n4842, n4841, n7139, n4840, n7137, n6902, n7145, 
		n5844, n5842, n5840, n5838, n7144, n5852, n5848, n5846, n7142, n4839, 
		n7147, n4838, n4837, n4836, n7150, n4835, n4834, n4833, n7135, n7136, 
		n4832, n7096, n7138, n7140, n4831, n7095, n7141, n7152, n5850, n7143, 
		n4830, n4829, n7085, n4828, n7154, n6934, n6972, n7159, n7151, n7086, 
		n4827, n4826, n7088, n4825, n7160, n6935, n6988, n7161, n7148, n7089, 
		n4824, n7130, n4823, n4822, n7162, n4821, n7129, n4820, n4819, n7163, 
		n4818, n7128, n4817, n4816, n7164, n5, n4815, n4814, n4813, n7165, 
		n6, n4812, n7131, n4811, n4810, n7166, n7, n4809, n7118, n4808, 
		n4807, n7167, n8, n4806, n4805, n7101, n4804, n7149, n9, n7102, 
		n4803, n7153, n6961, n4802, n7098, n7155, n7156, n4801, n7099, n7157, 
		n7158, n7146, n4800, n48, n4799, n4798, n4797, n7176, n4796, n7180, 
		n4795, n7177, n7188, n7190, n7187, n7194, n7197, n7196, n7195, n7202, 
		n7201, n7200, n7193, n7208, n7207, n7206, n7192, n7191, n4794, n4793, 
		n4792, n7215, n4791, n7170, n4790, n7218, n5295, n7189, n4789, n7220, 
		n5814, n7174, n4788, n7749, n4787, n7750, n4786, n4785, n7751, n4784, 
		n7752, n4783, n4782, n7753, n4781, n7754, n4780, n4779, n7755, n4778, 
		n7756, n4777, n4776, n7757, n4775, n7758, n4774, n4773, n7759, n4772, 
		n7760, n4771, n4770, n7761, n4769, n7762, n4768, n4767, n4766, n4765, 
		n4764, n7765, n4763, n7766, n4762, n4761, n7178, n7767, n7175, n7169, 
		n4760, n7181, n7769, n7179, n7171, n4759, n7184, n7182, n7173, n7770, 
		n4758, n7772, n4757, n7773, n4756, n7777, n7776, n7774, n4755, n7779, 
		n4754, n7781, n7778, n4753, n7785, n4752, n7783, n5813, n7212, n4751, 
		n7786, n5811, n4750, n7172, n5812, n7787, n7768, n4749, n7771, n4748, 
		n7216, n4747, n4746, n4745, n4744, n4743, n4742, n7793, n7796, n4741, 
		n4740, n4739, n7801, n7800, n7802, n7804, n4738, n4737, n4736, n7810, 
		n7809, n7811, n7814, n7807, n7820, n7818, n7826, n7827, n7816, n7835, 
		n7837, n7838, n7813, n7808, n7805, n7841, n7831, n7840, n7815, n7847, 
		n7845, n7850, n7852, n7853, n7851, n7849, n7819, n7844, n7858, n7828, 
		n7861, n7860, n7823, n7856, n7859, n7829, n7857, n7832, n7848, n7863, 
		n7824, n7864, n4735, n4734, n4733, n7865, n7806, n7868, n7867, n4732, 
		n4731, n7795, n7794, n4730, n7870, n7839, n7873, n7872, n7798, n7797, 
		n4729, n7878, n4728, n7881, n4727, n7875, n7825, n4726, n7886, n4725, 
		n7887, n4724, n7885, n7833, n7836, n7888, n4723, n7891, n4722, n7892, 
		n4721, n7890, n7889, n7884, n7843, n4720, n7894, n7877, n7876, n4719, 
		n7895, n7880, n7879, n4718, n7883, n7893, n7896, n7817, n7899, n7897, 
		n7900, n7830, n7821, n7855, n7822, n7862, n7901, n7842, n7902, n7834, 
		n7854, n7903, n7882, n7790, n7905, n7219, n7799, n7747, n7904, n7906, 
		n4717, n4716, n4715, n4714, n7912, n4713, n4712, n4711, n7916, n4710, 
		n4709, n7909, n4708, n7918, n7911, n4707, n7914, n4706, n4705, n4704, 
		n4703, n4702, n4701, n4700, n7792, n7791, n4699, n7846, n4698, n4697, 
		n4696, n4695, n4694, n4693, n4692, n4691, n4690, n6773, n7920, n4689, 
		n4688, n4687, n7926, n7925, n4686, n7931, n4685, n7935, n7934, n7924, 
		n7928, n7938, n4684, n7941, n4683, n7946, n7945, n4682, n7948, n7943, 
		n7940, n7950, n7952, n7954, n7951, n4681, n4680, n4679, n7960, n7966, 
		n7968, n7969, n7972, n7974, n7977, n7973, n7971, n7959, n7965, n4678, 
		n4677, n4676, n7979, n7982, n7984, n7985, n7989, n7990, n7988, n7994, 
		n7993, n7995, n7957, n8001, n8002, n8000, n7981, n4675, n4674, n4673, 
		n8011, n8015, n8013, n4672, n8020, n8019, n4671, n8023, n8021, n8024, 
		n8022, n4670, n8018, n8030, n8028, n4669, n4668, n8035, n4667, n8034, 
		n7917, n8036, n8025, n8033, n8027, n8026, n8038, n8040, n8039, n8037, 
		n8041, n4666, n4665, n4664, n8042, n8029, n8046, n8045, n8044, n8031, 
		n8051, n8043, n4663, n8053, n4662, n8056, n4661, n8059, n8058, n8055, 
		n4660, n4659, n8063, n4658, n8062, n8064, n8066, n8061, n4657, n7961, 
		n7944, n7923, n4656, n7963, n7947, n7929, n4655, n7964, n7936, n7933, 
		n8070, n8072, n8074, n8052, n8060, n8076, n8065, n8077, n7953, n8073, 
		n8079, n8068, n8075, n8078, n8069, n8082, n8054, n8057, n7922, n7907, 
		n8083, n8067, n8084, n8071, n4654, n4653, n8085, n8087, n4652, n8090, 
		n8089, n8088, n4651, n8092, n4650, n8091, n4649, n8095, n8094, n8093, 
		n4648, n8097, n4647, n8096, n8098, n4646, n8100, n8099, n8102, n4645, 
		n8103, n8101, n4644, n8086, n8105, n8104, n4643, n4642, n4641, n8109, 
		n8115, n8121, n8122, n4640, n4639, n4638, n8126, n8127, n8129, n8131, 
		n8130, n8123, n8136, n4637, n4636, n4635, n8139, n8140, n8142, n8143, 
		n8135, n8144, n4634, n4633, n4632, n8147, n8148, n8150, n8145, n4631, 
		n4630, n4629, n8155, n8156, n8158, n8160, n8151, n8152, n4628, n4627, 
		n4626, n8165, n8166, n8168, n8162, n8170, n4625, n4624, n4623, n8173, 
		n8174, n8169, n8176, n4622, n4621, n4620, n8179, n8180, n8183, n8181, 
		n8175, n8189, n4619, n4618, n4617, n8191, n8119, n8184, n8192, n8193, 
		n8195, n4616, n8108, n8110, n4615, n8111, n8112, n4614, n8114, n8197, 
		n8199, n8201, n8118, n8116, n8205, n8207, n8206, n7992, n8209, n7942, 
		n7949, n8208, n7956, n7991, n7997, n8210, n8215, n8214, n8212, n8216, 
		n7999, n8009, n8008, n8010, n8213, n8159, n8211, n8004, n7996, n8219, 
		n8222, n8221, n8224, n8220, n8003, n8226, n8005, n8225, n8006, n8223, 
		n7998, n8007, n7915, n8017, n7955, n8204, n7978, n8230, n8203, n8137, 
		n8128, n7967, n7939, n8233, n7930, n7937, n8235, n8239, n8240, n8238, 
		n8243, n8237, n8246, n8236, n7976, n7987, n8229, n8250, n8249, n8254, 
		n8248, n8257, n8234, n8263, n8264, n8262, n8267, n8261, n8269, n8260, 
		n8273, n8274, n8272, n8277, n8279, n8265, n8247, n8270, n8278, n8281, 
		n8268, n8280, n8275, n8276, n8284, n8283, n8271, n8289, n8282, n8188, 
		n8202, n8232, n8291, n8120, n8014, n7983, n8113, n4613, n4612, n8296, 
		n4611, n8294, n8047, n8302, n8149, n8200, n8253, n8301, n8182, n8167, 
		n8141, n8266, n8299, n4610, n8304, n4609, n4608, n4607, n8307, n4606, 
		n4605, n4604, n8292, n8293, n4603, n8252, n8295, n8297, n4602, n8251, 
		n8298, n8309, n8157, n8300, n4601, n4600, n8241, n46, n4599, n8311, 
		n8080, n8117, n8316, n8308, n8242, n4598, n4597, n8244, n4596, n8317, 
		n8081, n8227, n8318, n8305, n8245, n4595, n8286, n4594, n4593, n8319, 
		n4592, n8287, n4591, n4590, n8320, n4589, n4588, n4587, n8321, n4586, 
		n8285, n4585, n4584, n8322, n4583, n8288, n4582, n4581, n8323, n4580, 
		n4579, n4578, n8324, n4577, n4576, n8255, n4575, n8256, n8306, n4574, 
		n8310, n8106, n4573, n8258, n8312, n8313, n4572, n8259, n8314, n8315, 
		n8303, n4571, n4570, n4569, n4568, n8333, n4567, n8337, n4566, n8334, 
		n8345, n8347, n8344, n8351, n8354, n8353, n8352, n8359, n8358, n8357, 
		n8350, n8365, n8364, n8363, n8349, n8348, n4565, n4564, n4563, n8372, 
		n4562, n8327, n4561, n8375, n5292, n8346, n4560, n8377, n5819, n8331, 
		n4559, n8382, n4558, n8383, n4557, n4556, n8384, n4555, n8385, n4554, 
		n4553, n8386, n4552, n8387, n4551, n4550, n8388, n4549, n8389, n4548, 
		n4547, n8390, n4546, n8391, n4545, n4544, n8392, n4543, n8393, n4542, 
		n4541, n8394, n4540, n8395, n4539, n4538, n4537, n4536, n4535, n8398, 
		n4534, n8399, n4533, n4532, n8335, n8400, n8332, n8326, n4531, n8338, 
		n8402, n8336, n8328, n4530, n8341, n8339, n8330, n8403, n4529, n8405, 
		n4528, n8406, n4527, n8409, n8408, n8407, n4526, n8411, n4525, n8412, 
		n8410, n4524, n8414, n4523, n8413, n5818, n8369, n4522, n8415, n5816, 
		n4521, n8329, n5817, n8416, n8401, n4520, n8404, n4519, n8373, n4518, 
		n4517, n4516, n4515, n4514, n4513, n8422, n8425, n4512, n4511, n4510, 
		n8430, n8429, n8431, n8433, n4509, n4508, n4507, n8439, n8438, n8440, 
		n8443, n8436, n8449, n8447, n8455, n8456, n8445, n8464, n8466, n8467, 
		n8442, n8437, n8434, n8470, n8460, n8469, n8444, n8476, n8474, n8479, 
		n8481, n8482, n8480, n8478, n8448, n8473, n8487, n8457, n8490, n8489, 
		n8452, n8485, n8488, n8458, n8486, n8461, n8477, n8492, n8453, n8493, 
		n4506, n4505, n4504, n8494, n8435, n8497, n8496, n4503, n4502, n8424, 
		n8423, n4501, n8499, n8468, n8502, n8501, n8427, n8426, n4500, n8507, 
		n45, n4499, n8510, n4498, n8504, n8454, n4497, n8515, n4496, n8516, 
		n4495, n8514, n8462, n8465, n8517, n5984, n4494, n8520, n4493, n8521, 
		n4492, n8519, n8518, n8513, n8472, n4491, n8523, n8506, n8505, n4490, 
		n8524, n8509, n8508, n4489, n8512, n8522, n8525, n8446, n8528, n8526, 
		n8529, n8459, n8450, n8484, n8451, n8491, n8530, n8471, n8531, n8463, 
		n8483, n8532, n8511, n8419, n8534, n8376, n8428, n8380, n8533, n8535, 
		n4488, n4486, n4485, n8541, n4484, n4483, n4482, n8545, n4481, n4480, 
		n8538, n4479, n8547, n8540, n4478, n8543, n4477, n4476, n4475, n4474, 
		n4473, n4472, n4471, n8421, n6118, n5999, n8549, n5874, n8550, n8551, 
		n8420, n4470, n8475, n4469, n4468, n4467, n4466, n4465, n4464, n4463, 
		n4462, n4461, n8553, n8559, n8558, n8557, n8556, n8564, n8552, n8569, 
		n8568, n8567, n8566, n8575, n8574, n8573, n4460, n7921, n8579, n4459, 
		n4458, n4457, n8584, n8583, n4456, n8589, n8588, n4455, n8592, n8585, 
		n8582, n8595, n4454, n8600, n4453, n8603, n4452, n8606, n8605, n8602, 
		n8607, n8599, n8610, n8609, n8613, n4451, n4450, n8622, n4449, n8620, 
		n8624, n8626, n8627, n8630, n8632, n8635, n8631, n8629, n8611, n4448, 
		n4447, n8639, n4446, n8638, n8640, n8642, n8643, n8646, n8647, n8645, 
		n8651, n8650, n8652, n8616, n8658, n8659, n8657, n4445, n4444, n8670, 
		n4443, n8669, n8672, n4442, n8676, n8675, n4441, n8679, n8678, n4440, 
		n8680, n8677, n8683, n8674, n8686, n4439, n4438, n4437, n8688, n8546, 
		n8690, n8684, n8694, n8681, n8682, n8695, n8697, n8696, n8691, n8698, 
		n8689, n4436, n4435, n4434, n8699, n8685, n8703, n8702, n8701, n8687, 
		n8708, n8700, n4433, n8712, n8711, n4432, n8715, n8714, n4431, n8716, 
		n8713, n4430, n4429, n4428, n8720, n8722, n8724, n8719, n8721, n4427, 
		n8618, n8586, n8581, n4426, n8587, n8621, n8590, n4425, n8623, n8594, 
		n8591, n8728, n8730, n8732, n8710, n8718, n8734, n8723, n8735, n8598, 
		n8731, n8737, n8726, n8733, n8736, n8727, n8740, n8717, n8580, n8536, 
		n8741, n8725, n8742, n8729, n4424, n4423, n8743, n8745, n4422, n8748, 
		n8746, n8747, n4421, n8750, n4420, n8749, n4419, n8753, n8752, n8751, 
		n4418, n8755, n4417, n8754, n8757, n8756, n4416, n8758, n4415, n8761, 
		n8760, n8759, n4414, n8744, n8763, n8762, n4413, n4412, n4411, n8767, 
		n8773, n8778, n8780, n4410, n4409, n4408, n8783, n8784, n8787, n8785, 
		n8779, n8792, n4407, n4406, n4405, n8794, n8795, n8796, n8791, n8799, 
		n4404, n4403, n4402, n8801, n8802, n8804, n8798, n8806, n4401, n4400, 
		n4399, n8808, n8809, n8810, n8805, n8813, n4398, n4397, n4396, n8816, 
		n8817, n8819, n8812, n8821, n4395, n4394, n4393, n8824, n8825, n8820, 
		n8827, n4392, n4391, n4390, n8829, n8830, n8832, n8788, n8831, n8826, 
		n8835, n4389, n4388, n4387, n8838, n8777, n8839, n8834, n8840, n4386, 
		n8766, n8768, n4385, n8770, n91, n8769, n4384, n8772, n90, n8842, 
		n8844, n8846, n8776, n8774, n8850, n8852, n8851, n8649, n8854, n8601, 
		n8604, n8853, n8615, n8648, n8654, n8855, n8860, n8859, n8666, n8857, 
		n8661, n8862, n8665, n8861, n8656, n8667, n8858, n8856, n8653, n8863, 
		n8868, n8867, n8865, n8664, n8663, n8662, n8866, n8814, n8869, n8655, 
		n8864, n8660, n8544, n8612, n8614, n8849, n8636, n8872, n8848, n8781, 
		n8786, n8625, n8597, n8874, n8593, n8608, n8596, n8876, n8880, n8881, 
		n8879, n8884, n8878, n8887, n8877, n8634, n8644, n8871, n8891, n8890, 
		n8895, n8889, n8898, n8875, n8904, n8905, n8903, n8908, n8902, n8910, 
		n8901, n8914, n8915, n8913, n8918, n8920, n8906, n8888, n8911, n8919, 
		n8922, n8909, n8921, n8916, n8917, n8925, n8924, n8912, n8930, n8923, 
		n8841, n8847, n8873, n8932, n8560, n8570, n8671, n8641, n8555, n8933, 
		n8822, n8934, n8823, n8565, n8935, n8765, n8790, n8936, n8782, n8931, 
		n8578, n8938, n8807, n8937, n8561, n8939, n8843, n8562, n8940, n8793, 
		n8576, n8941, n8800, n8577, n8942, n8815, n8572, n8833, n8943, n8828, 
		n8571, n8836, n8944, n8837, n8706, n8771, n8707, n4383, n4382, n8949, 
		n4381, n8947, n8704, n8955, n8803, n8845, n8894, n8954, n8870, n8818, 
		n8797, n8907, n8952, n4380, n8957, n4379, n4378, n4377, n8960, n4376, 
		n4375, n4374, n8945, n8946, n4373, n8893, n8948, n8950, n4372, n8892, 
		n8951, n8962, n8811, n8953, n6529, n4371, n4370, n8882, n4369, n8965, 
		n8738, n8775, n8970, n8961, n8883, n4368, n4367, n8885, n4366, n8971, 
		n8739, n8789, n8972, n8958, n8705, n8886, n4365, n8927, n4364, n4363, 
		n8973, n99, n4362, n8926, n4361, n4360, n8974, n98, n4359, n4358, 
		n4357, n8975, n97, n4356, n8929, n4355, n4354, n8976, n96, n4353, 
		n8928, n4352, n4351, n8977, n95, n4350, n4349, n4348, n8978, n94, 
		n4347, n4346, n8896, n4345, n8959, n93, n8897, n4344, n8964, n8764, 
		n4343, n8899, n8966, n8967, n4342, n8900, n8968, n8969, n8956, n92, 
		n4341, n4340, n4339, n4338, n4337, n4336, n4335, n4334, n4333, n4332, 
		n4331, n4330, n4329, n4328, n4327, n4326, n4325, n4324, n4323, n4322, 
		n4321, n4320, n4319, n8989, n4318, n4317, n4316, n4315, n4314, n6758, 
		n4313, n8994, n4312, n8996, n4311, n4310, n4309, n4308, n8997, n4487, 
		n4307, n4306, n4305, n9000, n4304, n4303, n4302, n9001, n4301, n4300, 
		n9003, n43, n4299, n9002, n4298, n8999, n8981, n4297, n8983, n8991, 
		n4296, n8985, n9004, n8992, n4295, n8982, n4294, n4293, n4292, n4291, 
		n4290, n4289, n4288, n4287, n4286, n4285, n4284, n4283, n4282, n4281, 
		n4280, n4279, n4278, n4277, n9006, n4276, n9008, n4275, n9010, n4274, 
		n9013, n9012, n4273, n9011, n9016, n9015, n9014, n9018, n4272, n9020, 
		n9021, n9022, n9017, n4271, n9023, n9025, n4270, n9027, n4269, n9028, 
		n9026, n4268, n9030, n4267, n9031, n9029, n4266, n9024, n9033, n4265, 
		n4264, n4263, n5796, n4262, n5797, n4261, n5798, n4260, n5804, n4259, 
		n5996, n4258, n6355, n4257, n9037, n6614, n4256, n9038, n6876, n4255, 
		n4254, n4253, n4252, n4251, n4250, n4249, n9045, n4248, n9047, n4247, 
		n4246, n4245, n4244, n9065, n4243, n4242, n9068, n4241, n9060, n4240, 
		n9062, n9072, n4239, n4238, n4237, n4236, n4235, n4234, n4233, n9075, 
		n4232, n9077, n4231, n5888, n4230, n4229, n4228, n9036, n9092, n9094, 
		n4227, n9039, n9098, n9100, n9099, n4226, n9040, n9093, n4225, n9091, 
		n9042, n9041, n9108, n9104, n9096, n9110, n9095, n9111, n9112, n9109, 
		n9105, n9101, n9113, n9107, n9102, n9114, n6265, n4224, n9044, n9117, 
		n9119, n4223, n9049, n9123, n9125, n9124, n4222, n9052, n9118, n4221, 
		n9116, n9056, n9055, n9135, n9129, n9121, n9137, n9120, n9138, n9139, 
		n9136, n9130, n9126, n9140, n9134, n9127, n9141, n6888, n4220, n9059, 
		n9144, n4219, n9064, n9149, n9151, n9150, n4218, n9067, n9145, n4217, 
		n9143, n9071, n9070, n9160, n9156, n9152, n9146, n9163, n9147, n9165, 
		n9161, n9154, n9153, n9167, n9159, n9169, n7927, n9168, n4216, n9074, 
		n9172, n9174, n4215, n9079, n9178, n9180, n9179, n4214, n9082, n9173, 
		n4213, n9171, n9086, n9085, n9188, n9184, n9176, n9190, n9175, n9191, 
		n9192, n9189, n9185, n9181, n9193, n5983, n9187, n9182, n9194, n8693, 
		n4212, n4211, n4210, n4209, n8984, n4208, n4207, n4206, n4205, n4204, 
		n4203, n9196, n9195, n9201, n9198, n9200, n9199, n9206, n9208, n9207, 
		n9205, n9214, n9213, n4202, n9220, n9204, n9222, n9219, n9210, n4201, 
		n9229, n9203, n9230, n9228, n9211, n9233, n4200, n9235, n9216, n9223, 
		n9237, n42, n4199, n9240, n9215, n9231, n9241, n4198, n9243, n9209, 
		n4197, n9244, n9218, n9246, n4196, n9245, n9249, n47, n8980, n9236, 
		n9248, n9212, n9227, n9224, n9226, n9234, n4195, n9252, n9202, n9217, 
		n9247, n9239, n9254, n9232, n9225, n9242, n9251, n9253, n9256, n9257, 
		n9221, n9197, n9255, n5982, n9250, n9259, n9238, n9263, n5925, n9264, 
		n5920, n9265, n5932, n9266, n9262, n5924, n9269, n5945, n5960, n5961, 
		n9268, n5926, n9270, n9267, n5889, n9261, n5919, n9272, n9271, n9273, 
		n5906, n5938, n5907, n5931, n9274, n9260, n5934, n9275, n5930, n9276, 
		n5935, n9277, n5904, n5942, n5943, n4194, n9279, n9278, n9284, n9283, 
		n9282, n9288, n9290, n9289, n9287, n9296, n9295, n4193, n9302, n9286, 
		n9304, n9301, n9291, n4192, n9312, n9285, n9313, n9311, n9298, n9316, 
		n4191, n9318, n9300, n9305, n9320, n4190, n9324, n9294, n4189, n9325, 
		n9299, n9327, n4188, n9326, n9330, n9329, n9292, n9310, n9306, n9309, 
		n6662, n9332, n4187, n9333, n9293, n9328, n9334, n9323, n9335, n9331, 
		n9336, n6560, n4186, n9338, n9337, n9343, n9340, n9342, n9341, n9348, 
		n9350, n9349, n9347, n9356, n9355, n4185, n9362, n9346, n9364, n9361, 
		n9352, n4184, n9371, n9345, n9372, n9370, n9353, n9375, n4183, n9377, 
		n9358, n9365, n9379, n4182, n9382, n9357, n9373, n9383, n4181, n9385, 
		n9351, n4180, n9386, n9360, n9388, n4179, n9387, n9391, n44, n8987, 
		n9378, n9393, n9390, n9354, n9369, n9366, n9368, n7812, n9395, n9376, 
		n4178, n9396, n9344, n9359, n9389, n9397, n9374, n7803, n9398, n9384, 
		n9363, n9339, n7788, n9400, n9367, n7919, n9381, n9394, n9399, n9392, 
		n9402, n9380, n9406, n7204, n9407, n7199, n9408, n7211, n9409, n9405, 
		n7203, n9412, n7748, n7763, n7764, n9411, n7205, n9413, n9410, n7168, 
		n9404, n7198, n9415, n9414, n9416, n7185, n7217, n7186, n7210, n9417, 
		n9403, n7213, n9418, n7209, n9419, n7214, n9420, n7183, n7253, n7746, 
		n4177, n9422, n6098, n9421, n9427, n9426, n9425, n9431, n9433, n9432, 
		n9430, n9439, n9438, n4176, n9445, n9429, n9447, n9444, n9434, n4175, 
		n9455, n9428, n9456, n9454, n9436, n9459, n4174, n9461, n9441, n9448, 
		n9463, n4173, n9466, n9440, n9457, n9467, n4172, n9469, n9437, n4171, 
		n9470, n9443, n9472, n4170, n9471, n9475, n9462, n9474, n9435, n9453, 
		n9449, n9452, n8441, n9478, n9460, n4169, n9479, n9451, n9424, n9442, 
		n9481, n9458, n8432, n9482, n9468, n9446, n9423, n8417, n9480, n9450, 
		n8548, n9465, n9473, n9484, n9477, n9485, n9483, n9476, n9486, n9464, 
		n9490, n8361, n9491, n8356, n9492, n8368, n9493, n9489, n8360, n9496, 
		n8381, n8396, n8397, n9495, n8362, n9497, n9494, n8325, n9488, n8355, 
		n9499, n9498, n9500, n8342, n8374, n8343, n8367, n9501, n9487, n8370, 
		n9502, n8366, n9503, n8371, n9504, n8340, n8378, n8379, n4168, n4167, 
		n4166, n4165, n4164, n4163, n4162, n4161, n4160, n7075, n9507, n7133, 
		n7021, n9508, n6996, n7049, n9506, n9510, n7043, n9511, n7044, n9509, 
		n9514, n7040, n9515, n7050, n9513, n7016, n9516, n7017, n9512, n6976, 
		n9517, n6962, n9505, n9521, n7024, n7029, n9522, n7026, n9520, n7034, 
		n7032, n9523, n7035, n9519, n6979, n6989, n9524, n6981, n9518, n9527, 
		n7009, n9528, n7010, n9526, n6994, n9529, n6997, n9525, n6995, n9530, 
		n7003, n6903, n4159, n4158, n4157, n4156, n4155, n8231, n9533, n8290, 
		n8163, n9534, n8133, n9532, n9538, n8171, n8217, n9539, n8172, n9537, 
		n8196, n8187, n9540, n8198, n9536, n8134, n9541, n8138, n9535, n9542, 
		n8218, n9543, n8107, n6131, n9531, n9547, n8124, n8132, n9548, n8125, 
		n9546, n8186, n8194, n9549, n8190, n9545, n8185, n8177, n9550, n8178, 
		n9544, n9553, n8228, n9554, n8146, n9552, n8161, n9555, n8164, n9551, 
		n8153, n9556, n8154, n8048, n4154, n4153, n4152, n4151, n4150, n4149, 
		n9319, n9303, n9557, n9308, n9280, n9558, n9297, n9314, n9322, n9560, 
		n9561, n9315, n9321, n9565, n6581, n9566, n6576, n9567, n6589, n9568, 
		n9564, n6580, n9571, n6600, n6616, n6617, n9570, n6582, n9572, n9569, 
		n6545, n9563, n6575, n9574, n9573, n9575, n6562, n6593, n6563, n6587, 
		n9576, n9562, n6588, n9577, n6586, n9578, n6590, n9579, n6597, n6598, 
		n6653, n9580, n9307, n9559, n6638, n9317, n9281, n9581, n6771, n4148, 
		n6096, n5994, n9583, n9582, n5981, n5944, n9584, n5940, n9585, n6755, 
		n9586, n4147, n4146, n4145, n4144, n4143, n4142, n4141, n4140, n4139, 
		n4138, n4137, n4136, n4135, n4134, n4133, n4132, n4130, n4129, n4128, 
		n4127, n4126, n4125, n4124, n4123, n4122, n4121, n4120, n4119, n4118, 
		n4117, n4116, n4115, n4114, n4113, n4112, n4111, n4110, n4109, n4108, 
		n4107, n4106, n4105, n4104, n4103, n4102, n4101, n4100, n41, n4099, 
		n4098, n4097, n4096, n9588, n9587, n68, n59, n6071, n9088, n9589, 
		n9089, n9590, n4095, n5789, n4094, n5790, n4093, n9592, n6121, n5791, 
		n4092, n6108, n5792, n4091, n5787, n5793, n4090, n6130, n6245, n6187, 
		n9593, n6240, n6203, n9594, n6207, n6198, n9595, n6189, n6264, n5788, 
		n5794, n4089, n4088, n4087, n9132, n6839, n4086, n6760, n4085, n4084, 
		n9600, n9133, n6812, n9603, n6864, n6809, n6823, n9604, n6814, n6836, 
		n6828, n9605, n6832, n4083, n4082, n4081, n9607, n7986, n4080, n7908, 
		n4079, n4078, n9158, n8016, n7958, n9613, n8012, n7975, n9614, n7980, 
		n7970, n9615, n7962, n4077, n4076, n4075, n9617, n8554, n4074, n8537, 
		n4073, n4072, n8563, n8673, n8617, n9623, n8668, n8633, n9624, n8637, 
		n8628, n9625, n8619, n4071, n5795, n4070, n4069, n5839, n4068, n5841, 
		n4067, n5843, n4066, n4065, n4064, n5849, n4063, n4062, n5853, n4061, 
		n9626, n9007, n9640, n9642, n9641, n9639, n9644, n9643, n4060, n5823, 
		n4059, n5825, n4058, n5827, n4057, n5829, n4056, n5831, n4055, n5833, 
		n4054, n5835, n4053, n5837, n4052, n9627, n9009, n9655, n9657, n5845, 
		n9656, n5851, n9654, n9659, n5847, n9658, n9638, n5822, n4051, n4050, 
		n4049, n9591, n9660, n4048, n4047, n5871, n70, n5867, n4046, n9662, 
		n4045, n9663, n4044, n9664, n4043, n6069, n9665, n4042, n6074, n9666, 
		n6101, n4041, n9667, n4040, n9668, n4039, n9669, n4038, n6719, n9670, 
		n4037, n6724, n9671, n6748, n4036, n8963, n9672, n6337, n9673, n4035, 
		n9674, n4034, n9675, n4033, n9676, n4032, n7869, n9677, n4031, n7874, 
		n9678, n7898, n4030, n9679, n4029, n9680, n4028, n9681, n4027, n8498, 
		n9682, n4026, n8503, n9683, n8527, n4025, n9684, n5855, n9687, n9689, 
		n9688, n9686, n9691, n9690, n4024, n9692, n9685, n5857, n9694, n9696, 
		n9695, n9693, n9698, n9697, n4023, n4022, n4021, n4020, n4019, n4018, 
		n4017, n4016, n4015, n4014, n4013, n4012, n4011, n4010, n4009, n4008, 
		n4007, n4006, n4005, n4004, n4003, n4002, n4001, n4000, n40, n4, 
		n3999, n3998, n3997, n3996, n3995, n3994, n3993, n3992, n3991, n3990, 
		n3989, n9090, n3988, n9097, n3987, n9103, n3986, n9106, n3985, n3984, 
		n3983, n9115, n3982, n9122, n3981, n9128, n3980, n9131, n3979, n3978, 
		n3977, n9142, n3976, n9148, n3975, n9155, n3974, n9157, n3973, n3972, 
		n3971, n3970, n9170, n3969, n9177, n3968, n9183, n3967, n9186, n3966, 
		n3965, n3964, n3963, n3962, n3961, n7932, n3960, n6281, n3959, n6939, 
		n3958, n8709, n3957, n5820, n9005, n39, n38, n37, n6278, n36, 
		n6279, n35, n8988, n34, n8990, n9258, n9699, n6066, n8993, n9700, 
		n33, n6639, n32, n8986, n31, n8995, n9401, n9701, n9702, n8998, 
		n9703, n3, n9661, n29, n6762, n28, n6765, n27, n9596, n26, 
		n9597, n25, n9598, n24, n9599, n23, n9601, n22, n9602, n21, 
		n6721, n20, n6716, n19, n9043, n18, n9046, n172, n6774, n171, 
		n170, n6904, n17, n9048, n169, n6905, n168, n9628, n167, n7789, 
		n166, n9629, n165, n9630, n164, n9631, n163, n9632, n162, n7910, 
		n161, n7913, n160, n9606, n16, n9050, n159, n9608, n158, n9609, 
		n157, n9633, n156, n9610, n155, n9611, n154, n9612, n153, n7871, 
		n152, n7866, n151, n9634, n150, n9635, n15, n9051, n149, n9636, 
		n148, n9637, n147, n9645, n146, n9058, n145, n9061, n144, n9063, 
		n143, n9164, n142, n9066, n141, n9162, n140, n9069, n14, n9053, 
		n139, n9166, n138, n8032, n137, n9646, n136, n9647, n135, n9648, 
		n134, n9649, n133, n132, n131, n130, n13, n9054, n129, n128, 
		n127, n9650, n126, n125, n124, n8049, n123, n8050, n122, n9704, 
		n9034, n9019, n9707, n9706, n9035, n4131, n9708, n9032, n9705, n121, 
		n9651, n120, n9652, n12, n9057, n119, n8418, n118, n8539, n117, 
		n8542, n116, n9616, n115, n9618, n114, n9619, n113, n9620, n112, 
		n9621, n111, n9622, n110, n8500, n11, n9653, n109, n8495, n108, 
		n9073, n107, n9076, n106, n9078, n105, n9080, n104, n9081, n103, 
		n9083, n102, n9084, n101, n9087, n100, n8692, n10, n8979, n9712, 
		n9714, n9716, n9719, n9720, n9711, n9710, n9730, n9734, n9733, n9732, 
		n9729, n9741, n9728, n9746, n9744, n9727, n9709, n9751, n9756, n9759, 
		n9760, n9755, n9763, n9754, n9765, n9753, n9768, n9772, n9773, n9725, 
		n9774, n9761, n9715, n9758, n9735, n9757, n9736, n9771, n9781, n9743, 
		n9742, n9739, n9762, n9723, n9770, n9782, n9766, n9740, n9749, n9779, 
		n9764, n9748, n9780, n9738, n9745, n9776, n9769, n9784, n9750, n9767, 
		n9747, n9778, n9717, n9737, n9783, n9787, n9786, n9788, n9789, n9721, 
		n9722, n9785, n9775, n9731, n9752, n9791, n9724, n9718, n9726, n9790, 
		n9777, n9713, n5858, troj6_0_n1, troj6_0_n2, tempn4402, Trigger_en_6_0;

	dfxbp_1 DFF_0_Q_reg( .D(n3), .CLK(CLK), .Q_N(n5361) );
	dfxtp_1 DFF_31_Q_reg( .D(n4288), .CLK(CLK), .Q(n7281) );
	dfxtp_1 DFF_28_Q_reg( .D(n4286), .CLK(CLK), .Q(n7280) );
	dfxtp_1 DFF_1611_Q_reg( .D(n70), .CLK(CLK), .Q(g5388) );
	dfxbp_1 DFF_1612_Q_reg( .D(n5272), .CLK(CLK), .Q(n10033) );
	dfxtp_1 DFF_17_Q_reg( .D(n3), .CLK(CLK), .Q(g8021) );
	dfxbp_1 DFF_18_Q_reg( .D(n4278), .CLK(CLK), .Q(n10032) );
	dfxtp_1 DFF_29_Q_reg( .D(n4051), .CLK(CLK), .Q(g2962) );
	dfxbp_1 DFF_16_Q_reg( .D(n4277), .CLK(CLK), .Q_N(n15168) );
	dfxtp_1 DFF_20_Q_reg( .D(n4050), .CLK(CLK), .Q(g2934) );
	dfxbp_1 DFF_15_Q_reg( .D(n4276), .CLK(CLK), .Q_N(n15169) );
	dfxbp_1 DFF_4_Q_reg( .D(n122), .CLK(CLK), .Q(n10081) );
	dfxbp_1 DFF_6_Q_reg( .D(n4267), .CLK(CLK), .Q(n10084) );
	dfxtp_1 DFF_10_Q_reg( .D(n4271), .CLK(CLK), .Q(n7247) );
	dfxbp_1 DFF_12_Q_reg( .D(n4273), .CLK(CLK), .Q(n10065), .Q_N(n5369) );
	dfxbp_1 DFF_14_Q_reg( .D(n4275), .CLK(CLK), .Q(n10066) );
	dfxbp_1 DFF_1_Q_reg( .D(n4264), .CLK(CLK), .Q_N(n14868) );
	dfxbp_1 DFF_2_Q_reg( .D(n4265), .CLK(CLK), .Q_N(n14891) );
	dfxbp_1 DFF_1561_Q_reg( .D(n5259), .CLK(CLK), .Q_N(n15502) );
	dfxbp_1 DFF_1562_Q_reg( .D(n5260), .CLK(CLK), .Q_N(n14915) );
	dfxtp_1 DFF_1601_Q_reg( .D(n5262), .CLK(CLK), .Q(n7283) );
	dfxbp_1 DFF_1602_Q_reg( .D(n5263), .CLK(CLK), .Q(n10082) );
	dfxbp_1 DFF_1605_Q_reg( .D(n5266), .CLK(CLK), .Q(n10083) );
	dfxbp_1 DFF_1607_Q_reg( .D(n5268), .CLK(CLK), .Q(n9956) );
	dfxbp_1 DFF_1608_Q_reg( .D(n5269), .CLK(CLK), .Q(n9955), .Q_N(n5370) );
	dfxbp_1 DFF_1610_Q_reg( .D(n5271), .CLK(CLK), .Q(n10034) );
	dfxbp_1 DFF_94_Q_reg( .D(n4295), .CLK(CLK), .Q(n10089), .Q_N(n5304) );
	dfxbp_1 DFF_709_Q_reg( .D(n4700), .CLK(CLK), .Q(n9972), .Q_N(n5591) );
	dfxtp_1 DFF_353_Q_reg( .D(n4231), .CLK(CLK), .Q(g5629) );
	dfxbp_1 DFF_355_Q_reg( .D(n4470), .CLK(CLK), .Q_N(n5356) );
	dfxbp_1 DFF_1409_Q_reg( .D(n5160), .CLK(CLK), .Q(n9960), .Q_N(n5589) );
	dfxtp_1 DFF_1053_Q_reg( .D(n4231), .CLK(CLK), .Q(g5695) );
	dfxbp_1 DFF_1055_Q_reg( .D(n4928), .CLK(CLK), .Q_N(n5354) );
	dfxbp_1 DFF_1059_Q_reg( .D(n4929), .CLK(CLK), .Q(n9965), .Q_N(n5590) );
	dfxbp_1 DFF_1157_Q_reg( .D(n4978), .CLK(CLK), .Q(n9963), .Q_N(n5362) );
	dfxbp_1 DFF_1159_Q_reg( .D(n4980), .CLK(CLK), .Q(n9962) );
	dfxbp_1 DFF_1161_Q_reg( .D(n5299), .CLK(CLK), .Q(n9952) );
	dfxbp_1 DFF_1163_Q_reg( .D(n4983), .CLK(CLK), .Q(n10070) );
	dfxbp_1 DFF_1165_Q_reg( .D(n4985), .CLK(CLK), .Q(n10068) );
	dfxbp_1 DFF_1167_Q_reg( .D(n4987), .CLK(CLK), .Q(n10072), .Q_N(n5366) );
	dfxbp_1 DFF_1168_Q_reg( .D(n4988), .CLK(CLK), .Q(n10071) );
	dfxtp_1 DFF_1403_Q_reg( .D(n4231), .CLK(CLK), .Q(g5747) );
	dfxbp_1 DFF_1405_Q_reg( .D(n5159), .CLK(CLK), .Q_N(n5353) );
	dfxbp_1 DFF_1507_Q_reg( .D(n5206), .CLK(CLK), .Q(n9958), .Q_N(n5357) );
	dfxbp_1 DFF_1509_Q_reg( .D(n5208), .CLK(CLK), .Q(n9957) );
	dfxbp_1 DFF_1511_Q_reg( .D(n5302), .CLK(CLK), .Q(n9951) );
	dfxbp_1 DFF_1513_Q_reg( .D(n5211), .CLK(CLK), .Q(n10040) );
	dfxbp_1 DFF_1515_Q_reg( .D(n5213), .CLK(CLK), .Q(n10038) );
	dfxbp_1 DFF_1517_Q_reg( .D(n5215), .CLK(CLK), .Q(n10042), .Q_N(n5365) );
	dfxbp_1 DFF_1518_Q_reg( .D(n5216), .CLK(CLK), .Q(n10041) );
	dfxbp_1 DFF_359_Q_reg( .D(n4471), .CLK(CLK), .Q(n9977), .Q_N(n5592) );
	dfxbp_1 DFF_457_Q_reg( .D(n4519), .CLK(CLK), .Q(n9975), .Q_N(n5364) );
	dfxbp_1 DFF_459_Q_reg( .D(n4521), .CLK(CLK), .Q(n9974) );
	dfxbp_1 DFF_461_Q_reg( .D(n5293), .CLK(CLK), .Q(n9954) );
	dfxbp_1 DFF_463_Q_reg( .D(n4524), .CLK(CLK), .Q(n10012) );
	dfxbp_1 DFF_465_Q_reg( .D(n4526), .CLK(CLK), .Q(n10011) );
	dfxbp_1 DFF_467_Q_reg( .D(n4528), .CLK(CLK), .Q(n10014), .Q_N(n5368) );
	dfxbp_1 DFF_468_Q_reg( .D(n4529), .CLK(CLK), .Q(n10013) );
	dfxtp_1 DFF_703_Q_reg( .D(n4231), .CLK(CLK), .Q(g5657) );
	dfxbp_1 DFF_705_Q_reg( .D(n4699), .CLK(CLK), .Q_N(n5355) );
	dfxbp_1 DFF_807_Q_reg( .D(n4748), .CLK(CLK), .Q(n9970), .Q_N(n5363) );
	dfxbp_1 DFF_809_Q_reg( .D(n4750), .CLK(CLK), .Q(n9969) );
	dfxbp_1 DFF_811_Q_reg( .D(n5296), .CLK(CLK), .Q(n9953) );
	dfxbp_1 DFF_813_Q_reg( .D(n4753), .CLK(CLK), .Q(n9990) );
	dfxbp_1 DFF_815_Q_reg( .D(n4755), .CLK(CLK), .Q(n9989) );
	dfxbp_1 DFF_817_Q_reg( .D(n4757), .CLK(CLK), .Q(n9992), .Q_N(n5367) );
	dfxbp_1 DFF_818_Q_reg( .D(n4758), .CLK(CLK), .Q(n9991) );
	dfxtp_1 DFF_1296_Q_reg( .D(n4036), .CLK(CLK), .Q(g2256) );
	dfxtp_1 DFF_946_Q_reg( .D(n4036), .CLK(CLK), .Q(g1562) );
	dfxtp_1 DFF_596_Q_reg( .D(n4036), .CLK(CLK), .Q(g868) );
	dfxtp_1 DFF_246_Q_reg( .D(n4036), .CLK(CLK), .Q(g180) );
	dfxtp_1 DFF_1297_Q_reg( .D(n3965), .CLK(CLK), .Q(g5637) );
	dfxtp_1 DFF_947_Q_reg( .D(n3964), .CLK(CLK), .Q(g5612) );
	dfxtp_1 DFF_597_Q_reg( .D(n3963), .CLK(CLK), .Q(g5595) );
	dfxtp_1 DFF_247_Q_reg( .D(n3962), .CLK(CLK), .Q(g5549) );
	dfxbp_1 DFF_1286_Q_reg( .D(n5103), .CLK(CLK), .Q(n10051) );
	dfxbp_1 DFF_1288_Q_reg( .D(n5105), .CLK(CLK), .Q(n10062), .Q_N(n5372) );
	dfxbp_1 DFF_1290_Q_reg( .D(n5107), .CLK(CLK), .Q(n10061) );
	dfxbp_1 DFF_1292_Q_reg( .D(n5109), .CLK(CLK), .Q(n10060), .Q_N(n5371) );
	dfxbp_1 DFF_1295_Q_reg( .D(n5112), .CLK(CLK), .Q(n10059) );
	dfxbp_1 DFF_936_Q_reg( .D(n4873), .CLK(CLK), .Q(n9967) );
	dfxbp_1 DFF_938_Q_reg( .D(n4875), .CLK(CLK), .Q(n10085) );
	dfxbp_1 DFF_940_Q_reg( .D(n4877), .CLK(CLK), .Q(n10086) );
	dfxbp_1 DFF_942_Q_reg( .D(n4879), .CLK(CLK), .Q(n10087), .Q_N(n5377) );
	dfxbp_1 DFF_945_Q_reg( .D(n4882), .CLK(CLK), .Q(n10088) );
	dfxbp_1 DFF_236_Q_reg( .D(n4414), .CLK(CLK), .Q(n10029) );
	dfxbp_1 DFF_238_Q_reg( .D(n4416), .CLK(CLK), .Q(n10028), .Q_N(n5374) );
	dfxbp_1 DFF_240_Q_reg( .D(n4418), .CLK(CLK), .Q(n10027) );
	dfxbp_1 DFF_242_Q_reg( .D(n4420), .CLK(CLK), .Q(n10026), .Q_N(n5373) );
	dfxbp_1 DFF_245_Q_reg( .D(n4423), .CLK(CLK), .Q(n10025) );
	dfxbp_1 DFF_586_Q_reg( .D(n4644), .CLK(CLK), .Q(n10001) );
	dfxbp_1 DFF_588_Q_reg( .D(n4646), .CLK(CLK), .Q(n10007) );
	dfxbp_1 DFF_590_Q_reg( .D(n4648), .CLK(CLK), .Q(n10006) );
	dfxbp_1 DFF_592_Q_reg( .D(n4650), .CLK(CLK), .Q(n10005), .Q_N(n5378) );
	dfxbp_1 DFF_595_Q_reg( .D(n4653), .CLK(CLK), .Q(n10004) );
	dfxtp_1 DFF_77_Q_reg( .D(n4068), .CLK(CLK), .Q(g4200) );
	dfxtp_1 DFF_310_Q_reg( .D(n93), .CLK(CLK), .Q(g286) );
	dfxbp_1 DFF_311_Q_reg( .D(n3998), .CLK(CLK), .Q(n10016) );
	dfxtp_1 DFF_450_Q_reg( .D(n4105), .CLK(CLK), .Q(g536) );
	dfxtp_1 DFF_199_Q_reg( .D(n4377), .CLK(CLK), .Q(n7441) );
	dfxtp_1 DFF_198_Q_reg( .D(n4376), .CLK(CLK), .Q(n7440) );
	dfxbp_1 DFF_197_Q_reg( .D(n4375), .CLK(CLK), .Q_N(n5401) );
	dfxbp_1 DFF_193_Q_reg( .D(n4371), .CLK(CLK), .Q_N(n5434) );
	dfxtp_1 DFF_192_Q_reg( .D(n4370), .CLK(CLK), .Q(n7433) );
	dfxtp_1 DFF_191_Q_reg( .D(n4369), .CLK(CLK), .Q(n7439) );
	dfxbp_1 DFF_169_Q_reg( .D(n4347), .CLK(CLK), .Q_N(n5436) );
	dfxtp_1 DFF_168_Q_reg( .D(n4346), .CLK(CLK), .Q(n7424) );
	dfxtp_1 DFF_167_Q_reg( .D(n4345), .CLK(CLK), .Q(n7434) );
	dfxtp_1 DFF_75_Q_reg( .D(n4067), .CLK(CLK), .Q(g3993) );
	dfxtp_1 DFF_308_Q_reg( .D(n94), .CLK(CLK), .Q(g284) );
	dfxbp_1 DFF_309_Q_reg( .D(n3997), .CLK(CLK), .Q(n10017) );
	dfxtp_1 DFF_449_Q_reg( .D(n4104), .CLK(CLK), .Q(g534) );
	dfxbp_1 DFF_172_Q_reg( .D(n4350), .CLK(CLK), .Q_N(n5358) );
	dfxbp_1 DFF_171_Q_reg( .D(n4349), .CLK(CLK), .Q(n9861), .Q_N(n5662) );
	dfxbp_1 DFF_170_Q_reg( .D(n4348), .CLK(CLK), .Q(n9862), .Q_N(n5642) );
	dfxtp_1 DFF_69_Q_reg( .D(n4064), .CLK(CLK), .Q(g4321) );
	dfxtp_1 DFF_302_Q_reg( .D(n97), .CLK(CLK), .Q(g454) );
	dfxbp_1 DFF_303_Q_reg( .D(n3994), .CLK(CLK), .Q(n10020) );
	dfxtp_1 DFF_446_Q_reg( .D(n4101), .CLK(CLK), .Q(g531) );
	dfxbp_1 DFF_181_Q_reg( .D(n4359), .CLK(CLK), .Q(n10030), .Q_N(n5376) );
	dfxbp_1 DFF_180_Q_reg( .D(n4358), .CLK(CLK), .Q_N(n5498) );
	dfxbp_1 DFF_179_Q_reg( .D(n4357), .CLK(CLK), .Q_N(n5329) );
	dfxtp_1 DFF_67_Q_reg( .D(n4063), .CLK(CLK), .Q(g4088) );
	dfxtp_1 DFF_300_Q_reg( .D(n98), .CLK(CLK), .Q(g452) );
	dfxbp_1 DFF_301_Q_reg( .D(n3993), .CLK(CLK), .Q(n10021) );
	dfxtp_1 DFF_445_Q_reg( .D(n4100), .CLK(CLK), .Q(g530) );
	dfxbp_1 DFF_183_Q_reg( .D(n4361), .CLK(CLK), .Q_N(n5497) );
	dfxbp_1 DFF_182_Q_reg( .D(n4360), .CLK(CLK), .Q_N(n5328) );
	dfxtp_1 DFF_65_Q_reg( .D(n4062), .CLK(CLK), .Q(g8249) );
	dfxtp_1 DFF_298_Q_reg( .D(n99), .CLK(CLK), .Q(g450) );
	dfxbp_1 DFF_299_Q_reg( .D(n3992), .CLK(CLK), .Q(n10022) );
	dfxtp_1 DFF_444_Q_reg( .D(n4099), .CLK(CLK), .Q(g529) );
	dfxtp_1 DFF_187_Q_reg( .D(n4365), .CLK(CLK), .Q(n7286) );
	dfxbp_1 DFF_186_Q_reg( .D(n4364), .CLK(CLK), .Q_N(n5496) );
	dfxbp_1 DFF_185_Q_reg( .D(n4363), .CLK(CLK), .Q_N(n5327) );
	dfxtp_1 DFF_49_Q_reg( .D(n4054), .CLK(CLK), .Q(g4090) );
	dfxtp_1 DFF_650_Q_reg( .D(n132), .CLK(CLK), .Q(g1139) );
	dfxbp_1 DFF_651_Q_reg( .D(n4001), .CLK(CLK), .Q(n9999) );
	dfxtp_1 DFF_795_Q_reg( .D(n4108), .CLK(CLK), .Q(g1216) );
	dfxbp_1 DFF_533_Q_reg( .D(n4591), .CLK(CLK), .Q_N(n5493) );
	dfxbp_1 DFF_532_Q_reg( .D(n4590), .CLK(CLK), .Q_N(n5324) );
	dfxtp_1 DFF_47_Q_reg( .D(n4053), .CLK(CLK), .Q(g8251) );
	dfxtp_1 DFF_648_Q_reg( .D(n133), .CLK(CLK), .Q(g1137) );
	dfxbp_1 DFF_649_Q_reg( .D(n4000), .CLK(CLK), .Q(n10000) );
	dfxtp_1 DFF_794_Q_reg( .D(n4107), .CLK(CLK), .Q(g1215) );
	dfxtp_1 DFF_537_Q_reg( .D(n4595), .CLK(CLK), .Q(n7285) );
	dfxbp_1 DFF_536_Q_reg( .D(n4594), .CLK(CLK), .Q_N(n5492) );
	dfxbp_1 DFF_535_Q_reg( .D(n4593), .CLK(CLK), .Q_N(n5323) );
	dfxtp_1 DFF_1350_Q_reg( .D(n45), .CLK(CLK), .Q(g2527) );
	dfxbp_1 DFF_1351_Q_reg( .D(n4017), .CLK(CLK), .Q(n10049) );
	dfxtp_1 DFF_1495_Q_reg( .D(n4124), .CLK(CLK), .Q(g2604) );
	dfxtp_1 DFF_1234_Q_reg( .D(n5051), .CLK(CLK), .Q(n7284) );
	dfxbp_1 DFF_1233_Q_reg( .D(n5050), .CLK(CLK), .Q_N(n5485) );
	dfxbp_1 DFF_1232_Q_reg( .D(n5049), .CLK(CLK), .Q_N(n5316) );
	dfxtp_1 DFF_79_Q_reg( .D(n4069), .CLK(CLK), .Q(g4450) );
	dfxtp_1 DFF_312_Q_reg( .D(n92), .CLK(CLK), .Q(g288) );
	dfxbp_1 DFF_313_Q_reg( .D(n3999), .CLK(CLK), .Q(n10015) );
	dfxtp_1 DFF_451_Q_reg( .D(n4106), .CLK(CLK), .Q(g537) );
	dfxtp_1 DFF_202_Q_reg( .D(n4380), .CLK(CLK), .Q(n7445) );
	dfxbp_1 DFF_201_Q_reg( .D(n4379), .CLK(CLK), .Q_N(n5413) );
	dfxtp_1 DFF_200_Q_reg( .D(n4378), .CLK(CLK), .Q(n7446) );
	dfxbp_1 DFF_190_Q_reg( .D(n4368), .CLK(CLK), .Q_N(n5435) );
	dfxtp_1 DFF_189_Q_reg( .D(n4367), .CLK(CLK), .Q(n7442) );
	dfxtp_1 DFF_188_Q_reg( .D(n4366), .CLK(CLK), .Q(n7444) );
	dfxbp_1 DFF_166_Q_reg( .D(n4344), .CLK(CLK), .Q_N(n5442) );
	dfxtp_1 DFF_165_Q_reg( .D(n4343), .CLK(CLK), .Q(n7435) );
	dfxtp_1 DFF_164_Q_reg( .D(n4342), .CLK(CLK), .Q(n7443) );
	dfxtp_1 DFF_73_Q_reg( .D(n4066), .CLK(CLK), .Q(g8175) );
	dfxtp_1 DFF_306_Q_reg( .D(n95), .CLK(CLK), .Q(g282) );
	dfxbp_1 DFF_307_Q_reg( .D(n3996), .CLK(CLK), .Q(n10018) );
	dfxtp_1 DFF_448_Q_reg( .D(n4103), .CLK(CLK), .Q(g533) );
	dfxbp_1 DFF_174_Q_reg( .D(n4352), .CLK(CLK), .Q_N(n5499) );
	dfxbp_1 DFF_173_Q_reg( .D(n4351), .CLK(CLK), .Q_N(n5330) );
	dfxtp_1 DFF_71_Q_reg( .D(n4065), .CLK(CLK), .Q(g8023) );
	dfxtp_1 DFF_304_Q_reg( .D(n96), .CLK(CLK), .Q(g280) );
	dfxbp_1 DFF_305_Q_reg( .D(n3995), .CLK(CLK), .Q(n10019) );
	dfxtp_1 DFF_447_Q_reg( .D(n4102), .CLK(CLK), .Q(g532) );
	dfxbp_1 DFF_177_Q_reg( .D(n4355), .CLK(CLK), .Q(n9859), .Q_N(n5661) );
	dfxbp_1 DFF_176_Q_reg( .D(n4354), .CLK(CLK), .Q(n9860), .Q_N(n5641) );
	dfxbp_1 DFF_196_Q_reg( .D(n4374), .CLK(CLK), .Q(n10031), .Q_N(n5678) );
	dfxtp_1 DFF_195_Q_reg( .D(n4373), .CLK(CLK), .Q(n7397) );
	dfxtp_1 DFF_194_Q_reg( .D(n4372), .CLK(CLK), .Q(n7398) );
	dfxbp_1 DFF_205_Q_reg( .D(n4383), .CLK(CLK), .Q(n9978), .Q_N(n5604) );
	dfxtp_1 DFF_204_Q_reg( .D(n4382), .CLK(CLK), .Q(n7390) );
	dfxtp_1 DFF_203_Q_reg( .D(n4381), .CLK(CLK), .Q(n7393) );
	dfxbp_1 DFF_276_Q_reg( .D(n4436), .CLK(CLK), .Q(n10023), .Q_N(n5632) );
	dfxbp_1 DFF_275_Q_reg( .D(n4435), .CLK(CLK), .Q_N(n5381) );
	dfxtp_1 DFF_274_Q_reg( .D(n4434), .CLK(CLK), .Q(n7631) );
	dfxbp_1 DFF_279_Q_reg( .D(n4439), .CLK(CLK), .Q_N(n5552) );
	dfxbp_1 DFF_278_Q_reg( .D(n4438), .CLK(CLK), .Q_N(n5342) );
	dfxtp_1 DFF_277_Q_reg( .D(n4437), .CLK(CLK), .Q(n7635) );
	dfxbp_1 DFF_382_Q_reg( .D(n4480), .CLK(CLK), .Q(n9837), .Q_N(n5660) );
	dfxtp_1 DFF_381_Q_reg( .D(n4479), .CLK(CLK), .Q(n7456) );
	dfxbp_1 DFF_380_Q_reg( .D(n4478), .CLK(CLK), .Q_N(n5424) );
	dfxtp_1 DFF_403_Q_reg( .D(n4030), .CLK(CLK), .Q(g558) );
	dfxtp_1 DFF_404_Q_reg( .D(n4488), .CLK(CLK), .Q(n7272) );
	dfxbp_1 DFF_97_Q_reg( .D(n4298), .CLK(CLK), .Q(n9884), .Q_N(n5718) );
	dfxbp_1 DFF_96_Q_reg( .D(n4297), .CLK(CLK), .Q(n9885), .Q_N(n5587) );
	dfxbp_1 DFF_95_Q_reg( .D(n4296), .CLK(CLK), .Q(n9985), .Q_N(n5588) );
	dfxtp_1 DFF_282_Q_reg( .D(n4442), .CLK(CLK), .Q(n7313) );
	dfxtp_1 DFF_281_Q_reg( .D(n4441), .CLK(CLK), .Q(n7314) );
	dfxbp_1 DFF_267_Q_reg( .D(n4427), .CLK(CLK), .Q(n10024), .Q_N(n5673) );
	dfxbp_1 DFF_266_Q_reg( .D(n4426), .CLK(CLK), .Q(n9839), .Q_N(n5634) );
	dfxtp_1 DFF_265_Q_reg( .D(n4425), .CLK(CLK), .Q(n7627) );
	dfxbp_1 DFF_270_Q_reg( .D(n4430), .CLK(CLK), .Q_N(n5553) );
	dfxbp_1 DFF_269_Q_reg( .D(n4429), .CLK(CLK), .Q_N(n5343) );
	dfxtp_1 DFF_268_Q_reg( .D(n4428), .CLK(CLK), .Q(n7622) );
	dfxtp_1 DFF_273_Q_reg( .D(n4433), .CLK(CLK), .Q(n7341) );
	dfxtp_1 DFF_272_Q_reg( .D(n4432), .CLK(CLK), .Q(n7342) );
	dfxbp_1 DFF_391_Q_reg( .D(n4486), .CLK(CLK), .Q(n9835), .Q_N(n5658) );
	dfxtp_1 DFF_390_Q_reg( .D(n4485), .CLK(CLK), .Q(n7462) );
	dfxbp_1 DFF_389_Q_reg( .D(n4484), .CLK(CLK), .Q_N(n5425) );
	dfxtp_1 DFF_401_Q_reg( .D(n4029), .CLK(CLK), .Q(g549) );
	dfxbp_1 DFF_121_Q_reg( .D(n4322), .CLK(CLK), .Q_N(n5383) );
	dfxbp_1 DFF_120_Q_reg( .D(n4321), .CLK(CLK), .Q_N(n5307) );
	dfxbp_1 DFF_119_Q_reg( .D(n4320), .CLK(CLK), .Q_N(n5384) );
	dfxtp_1 DFF_297_Q_reg( .D(n4457), .CLK(CLK), .Q(n7379) );
	dfxtp_1 DFF_296_Q_reg( .D(n4456), .CLK(CLK), .Q(n7380) );
	dfxtp_1 DFF_288_Q_reg( .D(n4448), .CLK(CLK), .Q(n7473) );
	dfxtp_1 DFF_287_Q_reg( .D(n4447), .CLK(CLK), .Q(n7474) );
	dfxbp_1 DFF_286_Q_reg( .D(n4446), .CLK(CLK), .Q(n9841), .Q_N(n5630) );
	dfxbp_1 DFF_388_Q_reg( .D(n4483), .CLK(CLK), .Q(n9836), .Q_N(n5659) );
	dfxtp_1 DFF_387_Q_reg( .D(n4482), .CLK(CLK), .Q(n7458) );
	dfxbp_1 DFF_386_Q_reg( .D(n4481), .CLK(CLK), .Q_N(n5426) );
	dfxtp_1 DFF_398_Q_reg( .D(n4028), .CLK(CLK), .Q(g543) );
	dfxtp_1 DFF_399_Q_reg( .D(n4154), .CLK(CLK), .Q(g544) );
	dfxbp_1 DFF_400_Q_reg( .D(n4487), .CLK(CLK), .Q_N(n15417) );
	dfxbp_1 DFF_109_Q_reg( .D(n4310), .CLK(CLK), .Q(n9924), .Q_N(n5579) );
	dfxbp_1 DFF_108_Q_reg( .D(n4309), .CLK(CLK), .Q(n9927), .Q_N(n5585) );
	dfxbp_1 DFF_107_Q_reg( .D(n4308), .CLK(CLK), .Q(n9983), .Q_N(n5569) );
	dfxtp_1 DFF_208_Q_reg( .D(n4386), .CLK(CLK), .Q(n7651) );
	dfxbp_1 DFF_207_Q_reg( .D(n4385), .CLK(CLK), .Q(n9848), .Q_N(n5736) );
	dfxbp_1 DFF_206_Q_reg( .D(n4384), .CLK(CLK), .Q(n9849), .Q_N(n5692) );
	dfxtp_1 DFF_223_Q_reg( .D(n4401), .CLK(CLK), .Q(n7649) );
	dfxbp_1 DFF_222_Q_reg( .D(n4400), .CLK(CLK), .Q(n9850), .Q_N(n5734) );
	dfxbp_1 DFF_221_Q_reg( .D(n4399), .CLK(CLK), .Q(n9851), .Q_N(n5690) );
	dfxtp_1 DFF_226_Q_reg( .D(n4404), .CLK(CLK), .Q(n7650) );
	dfxbp_1 DFF_225_Q_reg( .D(n4403), .CLK(CLK), .Q(n9852), .Q_N(n5733) );
	dfxbp_1 DFF_224_Q_reg( .D(n4402), .CLK(CLK), .Q(n9853), .Q_N(n5689) );
	dfxtp_1 DFF_285_Q_reg( .D(n4445), .CLK(CLK), .Q(n7469) );
	dfxtp_1 DFF_284_Q_reg( .D(n4444), .CLK(CLK), .Q(n7470) );
	dfxbp_1 DFF_283_Q_reg( .D(n4443), .CLK(CLK), .Q(n9840), .Q_N(n5631) );
	dfxtp_1 DFF_229_Q_reg( .D(n4407), .CLK(CLK), .Q(n7655) );
	dfxbp_1 DFF_228_Q_reg( .D(n4406), .CLK(CLK), .Q(n9846), .Q_N(n5732) );
	dfxbp_1 DFF_227_Q_reg( .D(n4405), .CLK(CLK), .Q(n9847), .Q_N(n5688) );
	dfxtp_1 DFF_232_Q_reg( .D(n4410), .CLK(CLK), .Q(n7657) );
	dfxbp_1 DFF_231_Q_reg( .D(n4409), .CLK(CLK), .Q_N(n5527) );
	dfxbp_1 DFF_230_Q_reg( .D(n4408), .CLK(CLK), .Q(n9856), .Q_N(n5713) );
	dfxtp_1 DFF_235_Q_reg( .D(n4413), .CLK(CLK), .Q(n7654) );
	dfxbp_1 DFF_234_Q_reg( .D(n4412), .CLK(CLK), .Q(n9843), .Q_N(n5731) );
	dfxbp_1 DFF_233_Q_reg( .D(n4411), .CLK(CLK), .Q(n9844), .Q_N(n5687) );
	dfxtp_1 DFF_291_Q_reg( .D(n4451), .CLK(CLK), .Q(n7471) );
	dfxtp_1 DFF_290_Q_reg( .D(n4450), .CLK(CLK), .Q(n7472) );
	dfxbp_1 DFF_289_Q_reg( .D(n4449), .CLK(CLK), .Q(n9842), .Q_N(n5629) );
	dfxtp_1 DFF_294_Q_reg( .D(n4454), .CLK(CLK), .Q(n7332) );
	dfxtp_1 DFF_293_Q_reg( .D(n4453), .CLK(CLK), .Q(n7334) );
	dfxtp_1 DFF_211_Q_reg( .D(n4389), .CLK(CLK), .Q(n7652) );
	dfxbp_1 DFF_210_Q_reg( .D(n4388), .CLK(CLK), .Q_N(n5529) );
	dfxbp_1 DFF_209_Q_reg( .D(n4387), .CLK(CLK), .Q(n9858), .Q_N(n5716) );
	dfxtp_1 DFF_214_Q_reg( .D(n4392), .CLK(CLK), .Q(n7656) );
	dfxbp_1 DFF_213_Q_reg( .D(n4391), .CLK(CLK), .Q_N(n5528) );
	dfxbp_1 DFF_212_Q_reg( .D(n4390), .CLK(CLK), .Q(n9857), .Q_N(n5715) );
	dfxtp_1 DFF_217_Q_reg( .D(n4395), .CLK(CLK), .Q(n7621) );
	dfxbp_1 DFF_216_Q_reg( .D(n4394), .CLK(CLK), .Q_N(n5526) );
	dfxbp_1 DFF_215_Q_reg( .D(n4393), .CLK(CLK), .Q(n9845), .Q_N(n5714) );
	dfxtp_1 DFF_220_Q_reg( .D(n4398), .CLK(CLK), .Q(n7653) );
	dfxbp_1 DFF_219_Q_reg( .D(n4397), .CLK(CLK), .Q(n9854), .Q_N(n5735) );
	dfxbp_1 DFF_218_Q_reg( .D(n4396), .CLK(CLK), .Q(n9855), .Q_N(n5691) );
	dfxtp_1 DFF_394_Q_reg( .D(n4077), .CLK(CLK), .Q(g471) );
	dfxtp_1 DFF_375_Q_reg( .D(n116), .CLK(CLK), .Q(g568) );
	dfxbp_1 DFF_376_Q_reg( .D(n4477), .CLK(CLK), .Q_N(n15652) );
	dfxtp_1 DFF_393_Q_reg( .D(n4076), .CLK(CLK), .Q(g468) );
	dfxtp_1 DFF_373_Q_reg( .D(n115), .CLK(CLK), .Q(g566) );
	dfxtp_1 DFF_374_Q_reg( .D(n4153), .CLK(CLK), .Q(g567) );
	dfxtp_1 DFF_392_Q_reg( .D(n4075), .CLK(CLK), .Q(g465) );
	dfxtp_1 DFF_371_Q_reg( .D(n114), .CLK(CLK), .Q(g574) );
	dfxbp_1 DFF_372_Q_reg( .D(n4476), .CLK(CLK), .Q(n9834) );
	dfxtp_1 DFF_395_Q_reg( .D(n4027), .CLK(CLK), .Q(g528) );
	dfxtp_1 DFF_396_Q_reg( .D(n3972), .CLK(CLK), .Q(g535) );
	dfxtp_1 DFF_397_Q_reg( .D(n4135), .CLK(CLK), .Q(g542) );
	dfxtp_1 DFF_261_Q_reg( .D(n4237), .CLK(CLK), .Q(g376) );
	dfxtp_1 DFF_345_Q_reg( .D(n106), .CLK(CLK), .Q(g382) );
	dfxbp_1 DFF_346_Q_reg( .D(n4467), .CLK(CLK), .Q_N(n15068) );
	dfxtp_1 DFF_260_Q_reg( .D(n4236), .CLK(CLK), .Q(g373) );
	dfxtp_1 DFF_343_Q_reg( .D(n105), .CLK(CLK), .Q(g380) );
	dfxbp_1 DFF_344_Q_reg( .D(n4466), .CLK(CLK), .Q_N(n15069) );
	dfxtp_1 DFF_258_Q_reg( .D(n4235), .CLK(CLK), .Q(g361) );
	dfxtp_1 DFF_339_Q_reg( .D(n104), .CLK(CLK), .Q(g367) );
	dfxbp_1 DFF_340_Q_reg( .D(n4465), .CLK(CLK), .Q_N(n15071) );
	dfxtp_1 DFF_257_Q_reg( .D(n4234), .CLK(CLK), .Q(g358) );
	dfxtp_1 DFF_337_Q_reg( .D(n103), .CLK(CLK), .Q(g365) );
	dfxbp_1 DFF_338_Q_reg( .D(n4464), .CLK(CLK), .Q_N(n15073) );
	dfxtp_1 DFF_264_Q_reg( .D(n4239), .CLK(CLK), .Q(g391) );
	dfxtp_1 DFF_351_Q_reg( .D(n108), .CLK(CLK), .Q(g397) );
	dfxbp_1 DFF_352_Q_reg( .D(n4469), .CLK(CLK), .Q_N(n15064) );
	dfxtp_1 DFF_263_Q_reg( .D(n4238), .CLK(CLK), .Q(g388) );
	dfxtp_1 DFF_349_Q_reg( .D(n107), .CLK(CLK), .Q(g395) );
	dfxbp_1 DFF_350_Q_reg( .D(n4468), .CLK(CLK), .Q_N(n15065) );
	dfxtp_1 DFF_347_Q_reg( .D(n3970), .CLK(CLK), .Q(g387) );
	dfxtp_1 DFF_348_Q_reg( .D(n4152), .CLK(CLK), .Q(g394) );
	dfxtp_1 DFF_335_Q_reg( .D(n3968), .CLK(CLK), .Q(g357) );
	dfxtp_1 DFF_336_Q_reg( .D(n4132), .CLK(CLK), .Q(g364) );
	dfxtp_1 DFF_341_Q_reg( .D(n3969), .CLK(CLK), .Q(g372) );
	dfxtp_1 DFF_342_Q_reg( .D(n4151), .CLK(CLK), .Q(g379) );
	dfxtp_1 DFF_255_Q_reg( .D(n4233), .CLK(CLK), .Q(g346) );
	dfxtp_1 DFF_333_Q_reg( .D(n102), .CLK(CLK), .Q(g352) );
	dfxbp_1 DFF_334_Q_reg( .D(n4463), .CLK(CLK), .Q_N(n15066) );
	dfxtp_1 DFF_254_Q_reg( .D(n4232), .CLK(CLK), .Q(g343) );
	dfxtp_1 DFF_331_Q_reg( .D(n101), .CLK(CLK), .Q(g350) );
	dfxbp_1 DFF_332_Q_reg( .D(n4462), .CLK(CLK), .Q_N(n15067) );
	dfxtp_1 DFF_329_Q_reg( .D(n3967), .CLK(CLK), .Q(g342) );
	dfxtp_1 DFF_330_Q_reg( .D(n4150), .CLK(CLK), .Q(g349) );
	dfxtp_1 DFF_385_Q_reg( .D(n4074), .CLK(CLK), .Q(g461) );
	dfxtp_1 DFF_369_Q_reg( .D(n113), .CLK(CLK), .Q(g572) );
	dfxbp_1 DFF_370_Q_reg( .D(n4475), .CLK(CLK), .Q_N(n15638) );
	dfxtp_1 DFF_384_Q_reg( .D(n4073), .CLK(CLK), .Q(g458) );
	dfxtp_1 DFF_367_Q_reg( .D(n112), .CLK(CLK), .Q(g570) );
	dfxtp_1 DFF_368_Q_reg( .D(n4134), .CLK(CLK), .Q(g571) );
	dfxtp_1 DFF_383_Q_reg( .D(n4072), .CLK(CLK), .Q(g455) );
	dfxtp_1 DFF_365_Q_reg( .D(n111), .CLK(CLK), .Q(g564) );
	dfxbp_1 DFF_366_Q_reg( .D(n4474), .CLK(CLK), .Q(n9838) );
	dfxtp_1 DFF_362_Q_reg( .D(n4026), .CLK(CLK), .Q(g513) );
	dfxtp_1 DFF_363_Q_reg( .D(n3971), .CLK(CLK), .Q(g523) );
	dfxtp_1 DFF_364_Q_reg( .D(n4133), .CLK(CLK), .Q(g524) );
	dfxbp_1 DFF_328_Q_reg( .D(n4461), .CLK(CLK), .Q_N(n15426) );
	dfxbp_1 DFF_317_Q_reg( .D(n4460), .CLK(CLK), .Q_N(n5394) );
	dfxtp_1 DFF_61_Q_reg( .D(n4060), .CLK(CLK), .Q(g7334) );
	dfxtp_1 DFF_662_Q_reg( .D(n125), .CLK(CLK), .Q(g975) );
	dfxbp_1 DFF_663_Q_reg( .D(n4007), .CLK(CLK), .Q(n9993) );
	dfxtp_1 DFF_801_Q_reg( .D(n4114), .CLK(CLK), .Q(g1223) );
	dfxtp_1 DFF_552_Q_reg( .D(n4610), .CLK(CLK), .Q(n7437) );
	dfxbp_1 DFF_551_Q_reg( .D(n4609), .CLK(CLK), .Q_N(n5412) );
	dfxtp_1 DFF_550_Q_reg( .D(n4608), .CLK(CLK), .Q(n7438) );
	dfxbp_1 DFF_540_Q_reg( .D(n4598), .CLK(CLK), .Q_N(n5433) );
	dfxtp_1 DFF_539_Q_reg( .D(n4597), .CLK(CLK), .Q(n7431) );
	dfxtp_1 DFF_538_Q_reg( .D(n4596), .CLK(CLK), .Q(n7436) );
	dfxbp_1 DFF_516_Q_reg( .D(n4574), .CLK(CLK), .Q_N(n5441) );
	dfxtp_1 DFF_515_Q_reg( .D(n4573), .CLK(CLK), .Q(n7423) );
	dfxtp_1 DFF_514_Q_reg( .D(n4572), .CLK(CLK), .Q(n7432) );
	dfxtp_1 DFF_59_Q_reg( .D(n4059), .CLK(CLK), .Q(g6895) );
	dfxtp_1 DFF_660_Q_reg( .D(n126), .CLK(CLK), .Q(g973) );
	dfxbp_1 DFF_661_Q_reg( .D(n4006), .CLK(CLK), .Q(n9994) );
	dfxtp_1 DFF_800_Q_reg( .D(n4113), .CLK(CLK), .Q(g1222) );
	dfxtp_1 DFF_549_Q_reg( .D(n4607), .CLK(CLK), .Q(n7430) );
	dfxtp_1 DFF_548_Q_reg( .D(n4606), .CLK(CLK), .Q(n7429) );
	dfxbp_1 DFF_547_Q_reg( .D(n4605), .CLK(CLK), .Q_N(n5400) );
	dfxbp_1 DFF_543_Q_reg( .D(n4601), .CLK(CLK), .Q_N(n5432) );
	dfxtp_1 DFF_542_Q_reg( .D(n4600), .CLK(CLK), .Q(n7421) );
	dfxtp_1 DFF_541_Q_reg( .D(n4599), .CLK(CLK), .Q(n7428) );
	dfxbp_1 DFF_519_Q_reg( .D(n4577), .CLK(CLK), .Q_N(n5440) );
	dfxtp_1 DFF_518_Q_reg( .D(n4576), .CLK(CLK), .Q(n7412) );
	dfxtp_1 DFF_517_Q_reg( .D(n4575), .CLK(CLK), .Q(n7422) );
	dfxtp_1 DFF_57_Q_reg( .D(n4058), .CLK(CLK), .Q(g6442) );
	dfxtp_1 DFF_658_Q_reg( .D(n128), .CLK(CLK), .Q(g971) );
	dfxbp_1 DFF_659_Q_reg( .D(n4005), .CLK(CLK), .Q(n9995) );
	dfxtp_1 DFF_799_Q_reg( .D(n4112), .CLK(CLK), .Q(g1220) );
	dfxbp_1 DFF_522_Q_reg( .D(n4580), .CLK(CLK), .Q_N(n5306) );
	dfxbp_1 DFF_521_Q_reg( .D(n4579), .CLK(CLK), .Q(n9827), .Q_N(n5657) );
	dfxbp_1 DFF_520_Q_reg( .D(n4578), .CLK(CLK), .Q(n9828), .Q_N(n5640) );
	dfxtp_1 DFF_55_Q_reg( .D(n4057), .CLK(CLK), .Q(g6225) );
	dfxtp_1 DFF_656_Q_reg( .D(n129), .CLK(CLK), .Q(g969) );
	dfxbp_1 DFF_657_Q_reg( .D(n4004), .CLK(CLK), .Q(n9996) );
	dfxtp_1 DFF_798_Q_reg( .D(n4111), .CLK(CLK), .Q(g1219) );
	dfxbp_1 DFF_524_Q_reg( .D(n4582), .CLK(CLK), .Q_N(n5495) );
	dfxbp_1 DFF_523_Q_reg( .D(n4581), .CLK(CLK), .Q_N(n5326) );
	dfxtp_1 DFF_53_Q_reg( .D(n4056), .CLK(CLK), .Q(g4590) );
	dfxtp_1 DFF_654_Q_reg( .D(n130), .CLK(CLK), .Q(g967) );
	dfxbp_1 DFF_655_Q_reg( .D(n4003), .CLK(CLK), .Q(n9997) );
	dfxtp_1 DFF_797_Q_reg( .D(n4110), .CLK(CLK), .Q(g1218) );
	dfxbp_1 DFF_527_Q_reg( .D(n4585), .CLK(CLK), .Q(n9825), .Q_N(n5656) );
	dfxbp_1 DFF_526_Q_reg( .D(n4584), .CLK(CLK), .Q(n9826), .Q_N(n5639) );
	dfxtp_1 DFF_51_Q_reg( .D(n4055), .CLK(CLK), .Q(g4323) );
	dfxtp_1 DFF_652_Q_reg( .D(n131), .CLK(CLK), .Q(g1141) );
	dfxbp_1 DFF_653_Q_reg( .D(n4002), .CLK(CLK), .Q(n9998) );
	dfxtp_1 DFF_796_Q_reg( .D(n4109), .CLK(CLK), .Q(g1217) );
	dfxbp_1 DFF_531_Q_reg( .D(n4589), .CLK(CLK), .Q(n10008), .Q_N(n5375) );
	dfxbp_1 DFF_530_Q_reg( .D(n4588), .CLK(CLK), .Q_N(n5494) );
	dfxbp_1 DFF_529_Q_reg( .D(n4587), .CLK(CLK), .Q_N(n5325) );
	dfxbp_1 DFF_555_Q_reg( .D(n4613), .CLK(CLK), .Q(n9973), .Q_N(n5603) );
	dfxtp_1 DFF_554_Q_reg( .D(n4612), .CLK(CLK), .Q(n7387) );
	dfxtp_1 DFF_553_Q_reg( .D(n4611), .CLK(CLK), .Q(n7389) );
	dfxbp_1 DFF_626_Q_reg( .D(n4666), .CLK(CLK), .Q(n10002), .Q_N(n5670) );
	dfxtp_1 DFF_625_Q_reg( .D(n4665), .CLK(CLK), .Q(n7630) );
	dfxbp_1 DFF_624_Q_reg( .D(n4664), .CLK(CLK), .Q(n9808), .Q_N(n5633) );
	dfxtp_1 DFF_631_Q_reg( .D(n4671), .CLK(CLK), .Q(n7584) );
	dfxbp_1 DFF_629_Q_reg( .D(n4669), .CLK(CLK), .Q_N(n5332) );
	dfxtp_1 DFF_628_Q_reg( .D(n4668), .CLK(CLK), .Q(n7634) );
	dfxbp_1 DFF_627_Q_reg( .D(n4667), .CLK(CLK), .Q_N(n5524) );
	dfxbp_1 DFF_732_Q_reg( .D(n4709), .CLK(CLK), .Q(n9806), .Q_N(n5655) );
	dfxtp_1 DFF_731_Q_reg( .D(n4708), .CLK(CLK), .Q(n7454) );
	dfxbp_1 DFF_730_Q_reg( .D(n4707), .CLK(CLK), .Q_N(n5421) );
	dfxtp_1 DFF_753_Q_reg( .D(n4035), .CLK(CLK), .Q(g1244) );
	dfxtp_1 DFF_99_Q_reg( .D(n4300), .CLK(CLK), .Q(n7640) );
	dfxbp_1 DFF_98_Q_reg( .D(n4299), .CLK(CLK), .Q_N(n5313) );
	dfxbp_1 DFF_100_Q_reg( .D(n4301), .CLK(CLK), .Q(n9950), .Q_N(n5717) );
	dfxtp_1 DFF_632_Q_reg( .D(n4672), .CLK(CLK), .Q(n7583) );
	dfxbp_1 DFF_546_Q_reg( .D(n4604), .CLK(CLK), .Q(n10009), .Q_N(n5677) );
	dfxtp_1 DFF_545_Q_reg( .D(n4603), .CLK(CLK), .Q(n7395) );
	dfxtp_1 DFF_544_Q_reg( .D(n4602), .CLK(CLK), .Q(n7396) );
	dfxtp_1 DFF_621_Q_reg( .D(n4661), .CLK(CLK), .Q(n7339) );
	dfxtp_1 DFF_623_Q_reg( .D(n4663), .CLK(CLK), .Q(n7340) );
	dfxbp_1 DFF_617_Q_reg( .D(n4657), .CLK(CLK), .Q(n10003), .Q_N(n5671) );
	dfxtp_1 DFF_616_Q_reg( .D(n4656), .CLK(CLK), .Q(n7626) );
	dfxbp_1 DFF_615_Q_reg( .D(n4655), .CLK(CLK), .Q(n9809), .Q_N(n5672) );
	dfxbp_1 DFF_620_Q_reg( .D(n4660), .CLK(CLK), .Q_N(n5333) );
	dfxtp_1 DFF_619_Q_reg( .D(n4659), .CLK(CLK), .Q(n7620) );
	dfxbp_1 DFF_618_Q_reg( .D(n4658), .CLK(CLK), .Q_N(n5525) );
	dfxbp_1 DFF_741_Q_reg( .D(n4715), .CLK(CLK), .Q(n9804), .Q_N(n5653) );
	dfxtp_1 DFF_740_Q_reg( .D(n4714), .CLK(CLK), .Q(n7461) );
	dfxbp_1 DFF_739_Q_reg( .D(n4713), .CLK(CLK), .Q_N(n5422) );
	dfxtp_1 DFF_751_Q_reg( .D(n4034), .CLK(CLK), .Q(g1235) );
	dfxbp_1 DFF_124_Q_reg( .D(n4325), .CLK(CLK), .Q(n9906), .Q_N(n5582) );
	dfxbp_1 DFF_123_Q_reg( .D(n4324), .CLK(CLK), .Q_N(n5308) );
	dfxbp_1 DFF_122_Q_reg( .D(n4323), .CLK(CLK), .Q_N(n5309) );
	dfxtp_1 DFF_647_Q_reg( .D(n4687), .CLK(CLK), .Q(n7378) );
	dfxtp_1 DFF_645_Q_reg( .D(n4685), .CLK(CLK), .Q(n7377) );
	dfxtp_1 DFF_638_Q_reg( .D(n4678), .CLK(CLK), .Q(n7468) );
	dfxbp_1 DFF_637_Q_reg( .D(n4677), .CLK(CLK), .Q(n9811), .Q_N(n5664) );
	dfxtp_1 DFF_636_Q_reg( .D(n4676), .CLK(CLK), .Q(n7467) );
	dfxbp_1 DFF_738_Q_reg( .D(n4712), .CLK(CLK), .Q(n9805), .Q_N(n5654) );
	dfxtp_1 DFF_737_Q_reg( .D(n4711), .CLK(CLK), .Q(n7457) );
	dfxbp_1 DFF_736_Q_reg( .D(n4710), .CLK(CLK), .Q_N(n5423) );
	dfxtp_1 DFF_748_Q_reg( .D(n4033), .CLK(CLK), .Q(g1229) );
	dfxbp_1 DFF_749_Q_reg( .D(n4716), .CLK(CLK), .Q_N(n14876) );
	dfxbp_1 DFF_750_Q_reg( .D(n31), .CLK(CLK), .Q(n9923) );
	dfxbp_1 DFF_112_Q_reg( .D(n4313), .CLK(CLK), .Q(n9916), .Q_N(n5578) );
	dfxtp_1 DFF_111_Q_reg( .D(n4312), .CLK(CLK), .Q(n7666) );
	dfxbp_1 DFF_110_Q_reg( .D(n4311), .CLK(CLK), .Q_N(n5311) );
	dfxtp_1 DFF_642_Q_reg( .D(n4682), .CLK(CLK), .Q(n7333) );
	dfxtp_1 DFF_558_Q_reg( .D(n4616), .CLK(CLK), .Q(n7643) );
	dfxbp_1 DFF_557_Q_reg( .D(n4615), .CLK(CLK), .Q_N(n5397) );
	dfxbp_1 DFF_556_Q_reg( .D(n4614), .CLK(CLK), .Q(n9817), .Q_N(n5712) );
	dfxtp_1 DFF_582_Q_reg( .D(n4640), .CLK(CLK), .Q(n7648) );
	dfxbp_1 DFF_581_Q_reg( .D(n4639), .CLK(CLK), .Q_N(n5537) );
	dfxbp_1 DFF_580_Q_reg( .D(n4638), .CLK(CLK), .Q(n9822), .Q_N(n5705) );
	dfxtp_1 DFF_585_Q_reg( .D(n4643), .CLK(CLK), .Q(n7645) );
	dfxbp_1 DFF_584_Q_reg( .D(n4642), .CLK(CLK), .Q(n9813), .Q_N(n5728) );
	dfxbp_1 DFF_583_Q_reg( .D(n4641), .CLK(CLK), .Q(n9814), .Q_N(n5685) );
	dfxtp_1 DFF_635_Q_reg( .D(n4675), .CLK(CLK), .Q(n7464) );
	dfxbp_1 DFF_634_Q_reg( .D(n4674), .CLK(CLK), .Q(n9810), .Q_N(n5665) );
	dfxtp_1 DFF_633_Q_reg( .D(n4673), .CLK(CLK), .Q(n7463) );
	dfxtp_1 DFF_576_Q_reg( .D(n4634), .CLK(CLK), .Q(n7642) );
	dfxbp_1 DFF_575_Q_reg( .D(n4633), .CLK(CLK), .Q_N(n5540) );
	dfxbp_1 DFF_574_Q_reg( .D(n4632), .CLK(CLK), .Q(n9820), .Q_N(n5707) );
	dfxtp_1 DFF_579_Q_reg( .D(n4637), .CLK(CLK), .Q(n7646) );
	dfxbp_1 DFF_578_Q_reg( .D(n4636), .CLK(CLK), .Q_N(n5536) );
	dfxbp_1 DFF_577_Q_reg( .D(n4635), .CLK(CLK), .Q(n9816), .Q_N(n5706) );
	dfxtp_1 DFF_641_Q_reg( .D(n4681), .CLK(CLK), .Q(n7466) );
	dfxbp_1 DFF_640_Q_reg( .D(n4680), .CLK(CLK), .Q(n9812), .Q_N(n5663) );
	dfxtp_1 DFF_639_Q_reg( .D(n4679), .CLK(CLK), .Q(n7465) );
	dfxtp_1 DFF_644_Q_reg( .D(n4684), .CLK(CLK), .Q(n7331) );
	dfxtp_1 DFF_561_Q_reg( .D(n4619), .CLK(CLK), .Q(n7644) );
	dfxbp_1 DFF_560_Q_reg( .D(n4618), .CLK(CLK), .Q_N(n5538) );
	dfxbp_1 DFF_559_Q_reg( .D(n4617), .CLK(CLK), .Q(n9824), .Q_N(n5711) );
	dfxtp_1 DFF_564_Q_reg( .D(n4622), .CLK(CLK), .Q(n7647) );
	dfxbp_1 DFF_563_Q_reg( .D(n4621), .CLK(CLK), .Q_N(n5539) );
	dfxbp_1 DFF_562_Q_reg( .D(n4620), .CLK(CLK), .Q(n9823), .Q_N(n5710) );
	dfxtp_1 DFF_567_Q_reg( .D(n4625), .CLK(CLK), .Q(n7618) );
	dfxbp_1 DFF_566_Q_reg( .D(n4624), .CLK(CLK), .Q_N(n5535) );
	dfxbp_1 DFF_565_Q_reg( .D(n4623), .CLK(CLK), .Q(n9815), .Q_N(n5709) );
	dfxtp_1 DFF_570_Q_reg( .D(n4628), .CLK(CLK), .Q(n7619) );
	dfxbp_1 DFF_569_Q_reg( .D(n4627), .CLK(CLK), .Q_N(n5541) );
	dfxbp_1 DFF_568_Q_reg( .D(n4626), .CLK(CLK), .Q(n9821), .Q_N(n5708) );
	dfxtp_1 DFF_573_Q_reg( .D(n4631), .CLK(CLK), .Q(n7641) );
	dfxbp_1 DFF_572_Q_reg( .D(n4630), .CLK(CLK), .Q(n9818), .Q_N(n5729) );
	dfxbp_1 DFF_571_Q_reg( .D(n4629), .CLK(CLK), .Q(n9819), .Q_N(n5686) );
	dfxtp_1 DFF_744_Q_reg( .D(n4083), .CLK(CLK), .Q(g1158) );
	dfxtp_1 DFF_725_Q_reg( .D(n160), .CLK(CLK), .Q(g1254) );
	dfxbp_1 DFF_726_Q_reg( .D(n4706), .CLK(CLK), .Q_N(n15647) );
	dfxtp_1 DFF_743_Q_reg( .D(n4082), .CLK(CLK), .Q(g1155) );
	dfxtp_1 DFF_723_Q_reg( .D(n159), .CLK(CLK), .Q(g1252) );
	dfxtp_1 DFF_724_Q_reg( .D(n4159), .CLK(CLK), .Q(g1253) );
	dfxtp_1 DFF_742_Q_reg( .D(n4081), .CLK(CLK), .Q(g1152) );
	dfxtp_1 DFF_721_Q_reg( .D(n158), .CLK(CLK), .Q(g1260) );
	dfxbp_1 DFF_722_Q_reg( .D(n4705), .CLK(CLK), .Q(n9803) );
	dfxtp_1 DFF_745_Q_reg( .D(n4032), .CLK(CLK), .Q(g1214) );
	dfxtp_1 DFF_746_Q_reg( .D(n3979), .CLK(CLK), .Q(g1221) );
	dfxtp_1 DFF_747_Q_reg( .D(n4139), .CLK(CLK), .Q(g1228) );
	dfxtp_1 DFF_678_Q_reg( .D(n4155), .CLK(CLK), .Q(g985) );
	dfxbp_1 DFF_667_Q_reg( .D(n4690), .CLK(CLK), .Q_N(n5568) );
	dfxtp_1 DFF_603_Q_reg( .D(n4240), .CLK(CLK), .Q(g1041) );
	dfxtp_1 DFF_679_Q_reg( .D(n139), .CLK(CLK), .Q(g1029) );
	dfxtp_1 DFF_680_Q_reg( .D(n4156), .CLK(CLK), .Q(g1036) );
	dfxtp_1 DFF_611_Q_reg( .D(n4245), .CLK(CLK), .Q(g1063) );
	dfxtp_1 DFF_695_Q_reg( .D(n144), .CLK(CLK), .Q(g1069) );
	dfxbp_1 DFF_696_Q_reg( .D(n4696), .CLK(CLK), .Q_N(n15058) );
	dfxtp_1 DFF_693_Q_reg( .D(n3976), .CLK(CLK), .Q(g1067) );
	dfxbp_1 DFF_694_Q_reg( .D(n4695), .CLK(CLK), .Q_N(n15059) );
	dfxtp_1 DFF_609_Q_reg( .D(n4244), .CLK(CLK), .Q(g1071) );
	dfxtp_1 DFF_691_Q_reg( .D(n143), .CLK(CLK), .Q(g1059) );
	dfxtp_1 DFF_692_Q_reg( .D(n4157), .CLK(CLK), .Q(g1066) );
	dfxtp_1 DFF_608_Q_reg( .D(n4243), .CLK(CLK), .Q(g1048) );
	dfxtp_1 DFF_689_Q_reg( .D(n142), .CLK(CLK), .Q(g1054) );
	dfxbp_1 DFF_690_Q_reg( .D(n4694), .CLK(CLK), .Q_N(n15061) );
	dfxtp_1 DFF_687_Q_reg( .D(n3975), .CLK(CLK), .Q(g1052) );
	dfxbp_1 DFF_688_Q_reg( .D(n4693), .CLK(CLK), .Q_N(n15063) );
	dfxtp_1 DFF_606_Q_reg( .D(n4242), .CLK(CLK), .Q(g1056) );
	dfxtp_1 DFF_685_Q_reg( .D(n141), .CLK(CLK), .Q(g1044) );
	dfxtp_1 DFF_686_Q_reg( .D(n4136), .CLK(CLK), .Q(g1051) );
	dfxtp_1 DFF_614_Q_reg( .D(n4247), .CLK(CLK), .Q(g1078) );
	dfxtp_1 DFF_701_Q_reg( .D(n146), .CLK(CLK), .Q(g1084) );
	dfxbp_1 DFF_702_Q_reg( .D(n4698), .CLK(CLK), .Q_N(n15054) );
	dfxtp_1 DFF_699_Q_reg( .D(n3977), .CLK(CLK), .Q(g1082) );
	dfxbp_1 DFF_700_Q_reg( .D(n4697), .CLK(CLK), .Q_N(n15055) );
	dfxtp_1 DFF_612_Q_reg( .D(n4246), .CLK(CLK), .Q(g1085) );
	dfxtp_1 DFF_697_Q_reg( .D(n145), .CLK(CLK), .Q(g1074) );
	dfxtp_1 DFF_698_Q_reg( .D(n4158), .CLK(CLK), .Q(g1081) );
	dfxtp_1 DFF_605_Q_reg( .D(n4241), .CLK(CLK), .Q(g1033) );
	dfxtp_1 DFF_683_Q_reg( .D(n140), .CLK(CLK), .Q(g1039) );
	dfxbp_1 DFF_684_Q_reg( .D(n4692), .CLK(CLK), .Q_N(n15056) );
	dfxtp_1 DFF_681_Q_reg( .D(n3974), .CLK(CLK), .Q(g1037) );
	dfxbp_1 DFF_682_Q_reg( .D(n4691), .CLK(CLK), .Q_N(n15057) );
	dfxtp_1 DFF_735_Q_reg( .D(n4080), .CLK(CLK), .Q(g1148) );
	dfxtp_1 DFF_719_Q_reg( .D(n156), .CLK(CLK), .Q(g1258) );
	dfxbp_1 DFF_720_Q_reg( .D(n4704), .CLK(CLK), .Q_N(n15631) );
	dfxtp_1 DFF_734_Q_reg( .D(n4079), .CLK(CLK), .Q(g1145) );
	dfxtp_1 DFF_717_Q_reg( .D(n155), .CLK(CLK), .Q(g1256) );
	dfxtp_1 DFF_718_Q_reg( .D(n4138), .CLK(CLK), .Q(g1257) );
	dfxtp_1 DFF_733_Q_reg( .D(n4078), .CLK(CLK), .Q(g1142) );
	dfxtp_1 DFF_715_Q_reg( .D(n154), .CLK(CLK), .Q(g1250) );
	dfxbp_1 DFF_716_Q_reg( .D(n4703), .CLK(CLK), .Q(n9807) );
	dfxtp_1 DFF_712_Q_reg( .D(n4031), .CLK(CLK), .Q(g1199) );
	dfxtp_1 DFF_713_Q_reg( .D(n3978), .CLK(CLK), .Q(g1209) );
	dfxtp_1 DFF_714_Q_reg( .D(n4137), .CLK(CLK), .Q(g1210) );
	dfxtp_1 DFF_998_Q_reg( .D(n171), .CLK(CLK), .Q(g1831) );
	dfxbp_1 DFF_999_Q_reg( .D(n4008), .CLK(CLK), .Q(n10080) );
	dfxtp_1 DFF_1144_Q_reg( .D(n4115), .CLK(CLK), .Q(g1909) );
	dfxbp_1 DFF_886_Q_reg( .D(n4823), .CLK(CLK), .Q_N(n5488) );
	dfxbp_1 DFF_885_Q_reg( .D(n4822), .CLK(CLK), .Q_N(n5319) );
	dfxtp_1 DFF_1362_Q_reg( .D(n38), .CLK(CLK), .Q(g2363) );
	dfxbp_1 DFF_1363_Q_reg( .D(n4023), .CLK(CLK), .Q(n10043) );
	dfxtp_1 DFF_1501_Q_reg( .D(n4130), .CLK(CLK), .Q(g2611) );
	dfxtp_1 DFF_1252_Q_reg( .D(n5069), .CLK(CLK), .Q(n7414) );
	dfxbp_1 DFF_1251_Q_reg( .D(n5068), .CLK(CLK), .Q_N(n5410) );
	dfxtp_1 DFF_1250_Q_reg( .D(n5067), .CLK(CLK), .Q(n7415) );
	dfxbp_1 DFF_1240_Q_reg( .D(n5057), .CLK(CLK), .Q_N(n5428) );
	dfxtp_1 DFF_1239_Q_reg( .D(n5056), .CLK(CLK), .Q(n7407) );
	dfxtp_1 DFF_1238_Q_reg( .D(n5055), .CLK(CLK), .Q(n7413) );
	dfxbp_1 DFF_1216_Q_reg( .D(n5033), .CLK(CLK), .Q_N(n5438) );
	dfxtp_1 DFF_1215_Q_reg( .D(n5032), .CLK(CLK), .Q(n7402) );
	dfxtp_1 DFF_1214_Q_reg( .D(n5031), .CLK(CLK), .Q(n7408) );
	dfxtp_1 DFF_1360_Q_reg( .D(n39), .CLK(CLK), .Q(g2361) );
	dfxbp_1 DFF_1361_Q_reg( .D(n4022), .CLK(CLK), .Q(n10044) );
	dfxtp_1 DFF_1500_Q_reg( .D(n4129), .CLK(CLK), .Q(g2610) );
	dfxtp_1 DFF_1249_Q_reg( .D(n5066), .CLK(CLK), .Q(n7406) );
	dfxtp_1 DFF_1248_Q_reg( .D(n5065), .CLK(CLK), .Q(n7405) );
	dfxbp_1 DFF_1247_Q_reg( .D(n5064), .CLK(CLK), .Q_N(n5398) );
	dfxbp_1 DFF_1243_Q_reg( .D(n5060), .CLK(CLK), .Q_N(n5427) );
	dfxtp_1 DFF_1242_Q_reg( .D(n5059), .CLK(CLK), .Q(n7400) );
	dfxtp_1 DFF_1241_Q_reg( .D(n5058), .CLK(CLK), .Q(n7404) );
	dfxbp_1 DFF_1219_Q_reg( .D(n5036), .CLK(CLK), .Q_N(n5437) );
	dfxtp_1 DFF_1218_Q_reg( .D(n5035), .CLK(CLK), .Q(n7399) );
	dfxtp_1 DFF_1217_Q_reg( .D(n5034), .CLK(CLK), .Q(n7401) );
	dfxtp_1 DFF_1358_Q_reg( .D(n40), .CLK(CLK), .Q(g2359) );
	dfxbp_1 DFF_1359_Q_reg( .D(n4021), .CLK(CLK), .Q(n10045) );
	dfxtp_1 DFF_1499_Q_reg( .D(n4128), .CLK(CLK), .Q(g2608) );
	dfxbp_1 DFF_1222_Q_reg( .D(n5039), .CLK(CLK), .Q_N(n5359) );
	dfxbp_1 DFF_1221_Q_reg( .D(n5038), .CLK(CLK), .Q(n9909), .Q_N(n5647) );
	dfxbp_1 DFF_1220_Q_reg( .D(n5037), .CLK(CLK), .Q(n9910), .Q_N(n5636) );
	dfxtp_1 DFF_1356_Q_reg( .D(n41), .CLK(CLK), .Q(g2357) );
	dfxbp_1 DFF_1357_Q_reg( .D(n4020), .CLK(CLK), .Q(n10046) );
	dfxtp_1 DFF_1498_Q_reg( .D(n4127), .CLK(CLK), .Q(g2607) );
	dfxtp_1 DFF_1225_Q_reg( .D(n5042), .CLK(CLK), .Q(n7287) );
	dfxbp_1 DFF_1224_Q_reg( .D(n5041), .CLK(CLK), .Q_N(n5487) );
	dfxbp_1 DFF_1223_Q_reg( .D(n5040), .CLK(CLK), .Q_N(n5318) );
	dfxtp_1 DFF_1354_Q_reg( .D(n42), .CLK(CLK), .Q(g2355) );
	dfxbp_1 DFF_1355_Q_reg( .D(n4019), .CLK(CLK), .Q(n10047) );
	dfxtp_1 DFF_1497_Q_reg( .D(n4126), .CLK(CLK), .Q(g2606) );
	dfxbp_1 DFF_1228_Q_reg( .D(n5045), .CLK(CLK), .Q_N(n5305) );
	dfxbp_1 DFF_1227_Q_reg( .D(n5044), .CLK(CLK), .Q(n9907), .Q_N(n5646) );
	dfxbp_1 DFF_1226_Q_reg( .D(n5043), .CLK(CLK), .Q(n9908), .Q_N(n5635) );
	dfxtp_1 DFF_1352_Q_reg( .D(n43), .CLK(CLK), .Q(g2529) );
	dfxbp_1 DFF_1353_Q_reg( .D(n4018), .CLK(CLK), .Q(n10048) );
	dfxtp_1 DFF_1496_Q_reg( .D(n4125), .CLK(CLK), .Q(g2605) );
	dfxbp_1 DFF_1231_Q_reg( .D(n5048), .CLK(CLK), .Q(n10063), .Q_N(n5379) );
	dfxbp_1 DFF_1230_Q_reg( .D(n5047), .CLK(CLK), .Q_N(n5486) );
	dfxbp_1 DFF_1229_Q_reg( .D(n5046), .CLK(CLK), .Q_N(n5317) );
	dfxtp_1 DFF_1348_Q_reg( .D(n46), .CLK(CLK), .Q(g2525) );
	dfxbp_1 DFF_1349_Q_reg( .D(n4016), .CLK(CLK), .Q(n10050) );
	dfxtp_1 DFF_1494_Q_reg( .D(n4123), .CLK(CLK), .Q(g2603) );
	dfxbp_1 DFF_1236_Q_reg( .D(n5053), .CLK(CLK), .Q_N(n5484) );
	dfxbp_1 DFF_1235_Q_reg( .D(n5052), .CLK(CLK), .Q_N(n5315) );
	dfxbp_1 DFF_1246_Q_reg( .D(n5063), .CLK(CLK), .Q(n10064), .Q_N(n5675) );
	dfxtp_1 DFF_1245_Q_reg( .D(n5062), .CLK(CLK), .Q(n7388) );
	dfxtp_1 DFF_1244_Q_reg( .D(n5061), .CLK(CLK), .Q(n7391) );
	dfxtp_1 DFF_1347_Q_reg( .D(n5146), .CLK(CLK), .Q(n7382) );
	dfxtp_1 DFF_1346_Q_reg( .D(n5145), .CLK(CLK), .Q(n7381) );
	dfxtp_1 DFF_1279_Q_reg( .D(n5096), .CLK(CLK), .Q(n7674) );
	dfxbp_1 DFF_1278_Q_reg( .D(n5095), .CLK(CLK), .Q_N(n5521) );
	dfxbp_1 DFF_1277_Q_reg( .D(n5094), .CLK(CLK), .Q(n9896), .Q_N(n5694) );
	dfxtp_1 DFF_1258_Q_reg( .D(n5075), .CLK(CLK), .Q(n7670) );
	dfxbp_1 DFF_1257_Q_reg( .D(n5074), .CLK(CLK), .Q_N(n5395) );
	dfxbp_1 DFF_1256_Q_reg( .D(n5073), .CLK(CLK), .Q(n9897), .Q_N(n5698) );
	dfxtp_1 DFF_1270_Q_reg( .D(n5087), .CLK(CLK), .Q(n7672) );
	dfxbp_1 DFF_1269_Q_reg( .D(n5086), .CLK(CLK), .Q(n9901), .Q_N(n5721) );
	dfxbp_1 DFF_1268_Q_reg( .D(n5085), .CLK(CLK), .Q(n9902), .Q_N(n5680) );
	dfxtp_1 DFF_1273_Q_reg( .D(n5090), .CLK(CLK), .Q(n7668) );
	dfxbp_1 DFF_1272_Q_reg( .D(n5089), .CLK(CLK), .Q(n9898), .Q_N(n5720) );
	dfxbp_1 DFF_1271_Q_reg( .D(n5088), .CLK(CLK), .Q(n9899), .Q_N(n5679) );
	dfxtp_1 DFF_1335_Q_reg( .D(n5134), .CLK(CLK), .Q(n7572) );
	dfxtp_1 DFF_1334_Q_reg( .D(n5133), .CLK(CLK), .Q(n7571) );
	dfxbp_1 DFF_1333_Q_reg( .D(n5132), .CLK(CLK), .Q(n9892), .Q_N(n5611) );
	dfxtp_1 DFF_1264_Q_reg( .D(n5081), .CLK(CLK), .Q(n7675) );
	dfxbp_1 DFF_1263_Q_reg( .D(n5080), .CLK(CLK), .Q_N(n5523) );
	dfxbp_1 DFF_1262_Q_reg( .D(n5079), .CLK(CLK), .Q(n9904), .Q_N(n5696) );
	dfxtp_1 DFF_1276_Q_reg( .D(n5093), .CLK(CLK), .Q(n7669) );
	dfxbp_1 DFF_1275_Q_reg( .D(n5092), .CLK(CLK), .Q_N(n5522) );
	dfxbp_1 DFF_1274_Q_reg( .D(n5091), .CLK(CLK), .Q(n9900), .Q_N(n5695) );
	dfxtp_1 DFF_1282_Q_reg( .D(n5099), .CLK(CLK), .Q(n7676) );
	dfxbp_1 DFF_1281_Q_reg( .D(n5098), .CLK(CLK), .Q_N(n5519) );
	dfxbp_1 DFF_1280_Q_reg( .D(n5097), .CLK(CLK), .Q(n9903), .Q_N(n5693) );
	dfxtp_1 DFF_1285_Q_reg( .D(n5102), .CLK(CLK), .Q(n7673) );
	dfxbp_1 DFF_1284_Q_reg( .D(n5101), .CLK(CLK), .Q_N(n5331) );
	dfxbp_1 DFF_1283_Q_reg( .D(n5100), .CLK(CLK), .Q_N(n5547) );
	dfxtp_1 DFF_1267_Q_reg( .D(n5084), .CLK(CLK), .Q(n7667) );
	dfxbp_1 DFF_1266_Q_reg( .D(n5083), .CLK(CLK), .Q(n9895), .Q_N(n5738) );
	dfxbp_1 DFF_1265_Q_reg( .D(n5082), .CLK(CLK), .Q_N(n5542) );
	dfxtp_1 DFF_1341_Q_reg( .D(n5140), .CLK(CLK), .Q(n7574) );
	dfxtp_1 DFF_1340_Q_reg( .D(n5139), .CLK(CLK), .Q(n7573) );
	dfxbp_1 DFF_1339_Q_reg( .D(n5138), .CLK(CLK), .Q(n9894), .Q_N(n5609) );
	dfxbp_1 DFF_1438_Q_reg( .D(n5172), .CLK(CLK), .Q(n9880), .Q_N(n5644) );
	dfxtp_1 DFF_1437_Q_reg( .D(n5171), .CLK(CLK), .Q(n7453) );
	dfxbp_1 DFF_1436_Q_reg( .D(n5170), .CLK(CLK), .Q_N(n5417) );
	dfxtp_1 DFF_1448_Q_reg( .D(n4044), .CLK(CLK), .Q(g2617) );
	dfxbp_1 DFF_1449_Q_reg( .D(n5176), .CLK(CLK), .Q_N(n14885) );
	dfxtp_1 DFF_1344_Q_reg( .D(n5143), .CLK(CLK), .Q(n7327) );
	dfxtp_1 DFF_1343_Q_reg( .D(n5142), .CLK(CLK), .Q(n7328) );
	dfxtp_1 DFF_1338_Q_reg( .D(n5137), .CLK(CLK), .Q(n7576) );
	dfxtp_1 DFF_1337_Q_reg( .D(n5136), .CLK(CLK), .Q(n7575) );
	dfxbp_1 DFF_1336_Q_reg( .D(n5135), .CLK(CLK), .Q(n9893), .Q_N(n5610) );
	dfxtp_1 DFF_1261_Q_reg( .D(n5078), .CLK(CLK), .Q(n7671) );
	dfxbp_1 DFF_1260_Q_reg( .D(n5077), .CLK(CLK), .Q_N(n5520) );
	dfxbp_1 DFF_1259_Q_reg( .D(n5076), .CLK(CLK), .Q(n9905), .Q_N(n5697) );
	dfxtp_1 DFF_1444_Q_reg( .D(n4095), .CLK(CLK), .Q(g2546) );
	dfxtp_1 DFF_1425_Q_reg( .D(n65), .CLK(CLK), .Q(g2642) );
	dfxbp_1 DFF_1426_Q_reg( .D(n5166), .CLK(CLK), .Q_N(n15635) );
	dfxtp_1 DFF_1443_Q_reg( .D(n4094), .CLK(CLK), .Q(g2543) );
	dfxtp_1 DFF_1423_Q_reg( .D(n64), .CLK(CLK), .Q(g2640) );
	dfxtp_1 DFF_1424_Q_reg( .D(n4168), .CLK(CLK), .Q(g2641) );
	dfxtp_1 DFF_1442_Q_reg( .D(n4093), .CLK(CLK), .Q(g2540) );
	dfxtp_1 DFF_1421_Q_reg( .D(n63), .CLK(CLK), .Q(g2648) );
	dfxbp_1 DFF_1422_Q_reg( .D(n5165), .CLK(CLK), .Q(n9878) );
	dfxtp_1 DFF_1445_Q_reg( .D(n4043), .CLK(CLK), .Q(g2602) );
	dfxtp_1 DFF_1446_Q_reg( .D(n3991), .CLK(CLK), .Q(g2609) );
	dfxtp_1 DFF_1447_Q_reg( .D(n4147), .CLK(CLK), .Q(g2616) );
	dfxtp_1 DFF_1311_Q_reg( .D(n4261), .CLK(CLK), .Q(g2451) );
	dfxtp_1 DFF_1395_Q_reg( .D(n54), .CLK(CLK), .Q(g2457) );
	dfxbp_1 DFF_1396_Q_reg( .D(n5156), .CLK(CLK), .Q_N(n15038) );
	dfxtp_1 DFF_1310_Q_reg( .D(n4260), .CLK(CLK), .Q(g2448) );
	dfxtp_1 DFF_1393_Q_reg( .D(n53), .CLK(CLK), .Q(g2455) );
	dfxbp_1 DFF_1394_Q_reg( .D(n5155), .CLK(CLK), .Q_N(n15039) );
	dfxtp_1 DFF_1308_Q_reg( .D(n4259), .CLK(CLK), .Q(g2436) );
	dfxtp_1 DFF_1389_Q_reg( .D(n52), .CLK(CLK), .Q(g2442) );
	dfxbp_1 DFF_1390_Q_reg( .D(n5154), .CLK(CLK), .Q_N(n15041) );
	dfxtp_1 DFF_1307_Q_reg( .D(n4258), .CLK(CLK), .Q(g2433) );
	dfxtp_1 DFF_1387_Q_reg( .D(n51), .CLK(CLK), .Q(g2440) );
	dfxbp_1 DFF_1388_Q_reg( .D(n5153), .CLK(CLK), .Q_N(n15043) );
	dfxtp_1 DFF_1314_Q_reg( .D(n4263), .CLK(CLK), .Q(g2466) );
	dfxtp_1 DFF_1401_Q_reg( .D(n56), .CLK(CLK), .Q(g2472) );
	dfxbp_1 DFF_1402_Q_reg( .D(n5158), .CLK(CLK), .Q_N(n15034) );
	dfxtp_1 DFF_1313_Q_reg( .D(n4262), .CLK(CLK), .Q(g2463) );
	dfxtp_1 DFF_1399_Q_reg( .D(n55), .CLK(CLK), .Q(g2470) );
	dfxbp_1 DFF_1400_Q_reg( .D(n5157), .CLK(CLK), .Q_N(n15035) );
	dfxtp_1 DFF_1397_Q_reg( .D(n3989), .CLK(CLK), .Q(g2462) );
	dfxtp_1 DFF_1398_Q_reg( .D(n4167), .CLK(CLK), .Q(g2469) );
	dfxtp_1 DFF_1385_Q_reg( .D(n3987), .CLK(CLK), .Q(g2432) );
	dfxtp_1 DFF_1386_Q_reg( .D(n4144), .CLK(CLK), .Q(g2439) );
	dfxtp_1 DFF_1391_Q_reg( .D(n3988), .CLK(CLK), .Q(g2447) );
	dfxtp_1 DFF_1392_Q_reg( .D(n4166), .CLK(CLK), .Q(g2454) );
	dfxtp_1 DFF_1305_Q_reg( .D(n4257), .CLK(CLK), .Q(g2421) );
	dfxtp_1 DFF_1383_Q_reg( .D(n50), .CLK(CLK), .Q(g2427) );
	dfxbp_1 DFF_1384_Q_reg( .D(n5152), .CLK(CLK), .Q_N(n15036) );
	dfxtp_1 DFF_1304_Q_reg( .D(n4256), .CLK(CLK), .Q(g2418) );
	dfxtp_1 DFF_1381_Q_reg( .D(n49), .CLK(CLK), .Q(g2425) );
	dfxbp_1 DFF_1382_Q_reg( .D(n5151), .CLK(CLK), .Q_N(n15037) );
	dfxtp_1 DFF_1379_Q_reg( .D(n3986), .CLK(CLK), .Q(g2417) );
	dfxtp_1 DFF_1380_Q_reg( .D(n4165), .CLK(CLK), .Q(g2424) );
	dfxtp_1 DFF_1435_Q_reg( .D(n4092), .CLK(CLK), .Q(g2536) );
	dfxtp_1 DFF_1419_Q_reg( .D(n62), .CLK(CLK), .Q(g2646) );
	dfxbp_1 DFF_1420_Q_reg( .D(n5164), .CLK(CLK), .Q_N(n15627) );
	dfxtp_1 DFF_1434_Q_reg( .D(n4091), .CLK(CLK), .Q(g2533) );
	dfxtp_1 DFF_1417_Q_reg( .D(n61), .CLK(CLK), .Q(g2644) );
	dfxtp_1 DFF_1418_Q_reg( .D(n4146), .CLK(CLK), .Q(g2645) );
	dfxtp_1 DFF_1433_Q_reg( .D(n4090), .CLK(CLK), .Q(g2530) );
	dfxtp_1 DFF_1415_Q_reg( .D(n60), .CLK(CLK), .Q(g2638) );
	dfxbp_1 DFF_1416_Q_reg( .D(n5163), .CLK(CLK), .Q(n9882) );
	dfxtp_1 DFF_1412_Q_reg( .D(n4042), .CLK(CLK), .Q(g2587) );
	dfxtp_1 DFF_1413_Q_reg( .D(n3990), .CLK(CLK), .Q(g2597) );
	dfxtp_1 DFF_1414_Q_reg( .D(n4145), .CLK(CLK), .Q(g2598) );
	dfxbp_1 DFF_1378_Q_reg( .D(n5150), .CLK(CLK), .Q_N(n14920) );
	dfxbp_1 DFF_1255_Q_reg( .D(n5072), .CLK(CLK), .Q(n9961), .Q_N(n5601) );
	dfxtp_1 DFF_1254_Q_reg( .D(n5071), .CLK(CLK), .Q(n7383) );
	dfxtp_1 DFF_1253_Q_reg( .D(n5070), .CLK(CLK), .Q(n7384) );
	dfxbp_1 DFF_1326_Q_reg( .D(n5125), .CLK(CLK), .Q(n10052), .Q_N(n5612) );
	dfxbp_1 DFF_1325_Q_reg( .D(n5124), .CLK(CLK), .Q_N(n5380) );
	dfxtp_1 DFF_1324_Q_reg( .D(n5123), .CLK(CLK), .Q(n7628) );
	dfxbp_1 DFF_1329_Q_reg( .D(n5128), .CLK(CLK), .Q_N(n5548) );
	dfxbp_1 DFF_1328_Q_reg( .D(n5127), .CLK(CLK), .Q_N(n5338) );
	dfxtp_1 DFF_1327_Q_reg( .D(n5126), .CLK(CLK), .Q(n7617) );
	dfxbp_1 DFF_1432_Q_reg( .D(n5169), .CLK(CLK), .Q(n9881), .Q_N(n5645) );
	dfxtp_1 DFF_1431_Q_reg( .D(n5168), .CLK(CLK), .Q(n7451) );
	dfxbp_1 DFF_1430_Q_reg( .D(n5167), .CLK(CLK), .Q_N(n5415) );
	dfxtp_1 DFF_1453_Q_reg( .D(n4046), .CLK(CLK), .Q(g2632) );
	dfxbp_1 DFF_106_Q_reg( .D(n4307), .CLK(CLK), .Q(n9984), .Q_N(n5737) );
	dfxbp_1 DFF_105_Q_reg( .D(n4306), .CLK(CLK), .Q(n9931), .Q_N(n5586) );
	dfxbp_1 DFF_104_Q_reg( .D(n4305), .CLK(CLK), .Q_N(n5314) );
	dfxtp_1 DFF_1332_Q_reg( .D(n5131), .CLK(CLK), .Q(n7310) );
	dfxtp_1 DFF_1331_Q_reg( .D(n5130), .CLK(CLK), .Q(n7309) );
	dfxbp_1 DFF_1317_Q_reg( .D(n5116), .CLK(CLK), .Q(n10058), .Q_N(n5666) );
	dfxbp_1 DFF_1316_Q_reg( .D(n5115), .CLK(CLK), .Q(n9889), .Q_N(n5667) );
	dfxtp_1 DFF_1315_Q_reg( .D(n5114), .CLK(CLK), .Q(n7624) );
	dfxbp_1 DFF_1320_Q_reg( .D(n5119), .CLK(CLK), .Q_N(n5549) );
	dfxbp_1 DFF_1319_Q_reg( .D(n5118), .CLK(CLK), .Q_N(n5339) );
	dfxtp_1 DFF_1318_Q_reg( .D(n5117), .CLK(CLK), .Q(n7677) );
	dfxtp_1 DFF_1323_Q_reg( .D(n5122), .CLK(CLK), .Q(n7336) );
	dfxtp_1 DFF_1322_Q_reg( .D(n5121), .CLK(CLK), .Q(n7335) );
	dfxbp_1 DFF_1441_Q_reg( .D(n5175), .CLK(CLK), .Q(n9879), .Q_N(n5643) );
	dfxtp_1 DFF_1440_Q_reg( .D(n5174), .CLK(CLK), .Q(n7459) );
	dfxbp_1 DFF_1439_Q_reg( .D(n5173), .CLK(CLK), .Q_N(n5416) );
	dfxtp_1 DFF_1451_Q_reg( .D(n4045), .CLK(CLK), .Q(g2623) );
	dfxbp_1 DFF_130_Q_reg( .D(n4331), .CLK(CLK), .Q(n9890), .Q_N(n5575) );
	dfxbp_1 DFF_129_Q_reg( .D(n4330), .CLK(CLK), .Q_N(n5386) );
	dfxbp_1 DFF_128_Q_reg( .D(n4329), .CLK(CLK), .Q(n9891), .Q_N(n5576) );
	dfxtp_1 DFF_1012_Q_reg( .D(n10), .CLK(CLK), .Q(g1669) );
	dfxbp_1 DFF_1013_Q_reg( .D(n4015), .CLK(CLK), .Q(n10073) );
	dfxtp_1 DFF_1151_Q_reg( .D(n4122), .CLK(CLK), .Q(g1917) );
	dfxtp_1 DFF_902_Q_reg( .D(n4839), .CLK(CLK), .Q(n7426) );
	dfxbp_1 DFF_901_Q_reg( .D(n4838), .CLK(CLK), .Q_N(n5411) );
	dfxtp_1 DFF_900_Q_reg( .D(n4837), .CLK(CLK), .Q(n7427) );
	dfxbp_1 DFF_890_Q_reg( .D(n4827), .CLK(CLK), .Q_N(n5430) );
	dfxtp_1 DFF_889_Q_reg( .D(n4826), .CLK(CLK), .Q(n7419) );
	dfxtp_1 DFF_888_Q_reg( .D(n4825), .CLK(CLK), .Q(n7425) );
	dfxbp_1 DFF_866_Q_reg( .D(n4803), .CLK(CLK), .Q_N(n5439) );
	dfxtp_1 DFF_865_Q_reg( .D(n4802), .CLK(CLK), .Q(n7411) );
	dfxtp_1 DFF_864_Q_reg( .D(n4801), .CLK(CLK), .Q(n7420) );
	dfxtp_1 DFF_1010_Q_reg( .D(n9), .CLK(CLK), .Q(g1667) );
	dfxbp_1 DFF_1011_Q_reg( .D(n4014), .CLK(CLK), .Q(n10074) );
	dfxtp_1 DFF_1150_Q_reg( .D(n4121), .CLK(CLK), .Q(g1916) );
	dfxtp_1 DFF_899_Q_reg( .D(n4836), .CLK(CLK), .Q(n7418) );
	dfxtp_1 DFF_898_Q_reg( .D(n4835), .CLK(CLK), .Q(n7417) );
	dfxbp_1 DFF_897_Q_reg( .D(n4834), .CLK(CLK), .Q_N(n5399) );
	dfxbp_1 DFF_893_Q_reg( .D(n4830), .CLK(CLK), .Q_N(n5429) );
	dfxtp_1 DFF_892_Q_reg( .D(n4829), .CLK(CLK), .Q(n7409) );
	dfxtp_1 DFF_891_Q_reg( .D(n4828), .CLK(CLK), .Q(n7416) );
	dfxbp_1 DFF_869_Q_reg( .D(n4806), .CLK(CLK), .Q_N(n5431) );
	dfxtp_1 DFF_868_Q_reg( .D(n4805), .CLK(CLK), .Q(n7403) );
	dfxtp_1 DFF_867_Q_reg( .D(n4804), .CLK(CLK), .Q(n7410) );
	dfxtp_1 DFF_1008_Q_reg( .D(n8), .CLK(CLK), .Q(g1665) );
	dfxbp_1 DFF_1009_Q_reg( .D(n4013), .CLK(CLK), .Q(n10075) );
	dfxtp_1 DFF_1149_Q_reg( .D(n4120), .CLK(CLK), .Q(g1914) );
	dfxbp_1 DFF_871_Q_reg( .D(n4808), .CLK(CLK), .Q(n9796), .Q_N(n5652) );
	dfxbp_1 DFF_870_Q_reg( .D(n4807), .CLK(CLK), .Q(n9797), .Q_N(n5638) );
	dfxtp_1 DFF_1006_Q_reg( .D(n7), .CLK(CLK), .Q(g1663) );
	dfxbp_1 DFF_1007_Q_reg( .D(n4012), .CLK(CLK), .Q(n10076) );
	dfxtp_1 DFF_1148_Q_reg( .D(n4119), .CLK(CLK), .Q(g1913) );
	dfxbp_1 DFF_874_Q_reg( .D(n4811), .CLK(CLK), .Q_N(n5491) );
	dfxbp_1 DFF_873_Q_reg( .D(n4810), .CLK(CLK), .Q_N(n5322) );
	dfxtp_1 DFF_1004_Q_reg( .D(n6), .CLK(CLK), .Q(g1661) );
	dfxbp_1 DFF_1005_Q_reg( .D(n4011), .CLK(CLK), .Q(n10077) );
	dfxtp_1 DFF_1147_Q_reg( .D(n4118), .CLK(CLK), .Q(g1912) );
	dfxbp_1 DFF_878_Q_reg( .D(n4815), .CLK(CLK), .Q_N(n5360) );
	dfxbp_1 DFF_877_Q_reg( .D(n4814), .CLK(CLK), .Q(n9794), .Q_N(n5651) );
	dfxbp_1 DFF_876_Q_reg( .D(n4813), .CLK(CLK), .Q(n9795), .Q_N(n5637) );
	dfxtp_1 DFF_1002_Q_reg( .D(n5), .CLK(CLK), .Q(g1835) );
	dfxbp_1 DFF_1003_Q_reg( .D(n4010), .CLK(CLK), .Q(n10078) );
	dfxtp_1 DFF_1146_Q_reg( .D(n4117), .CLK(CLK), .Q(g1911) );
	dfxbp_1 DFF_880_Q_reg( .D(n4817), .CLK(CLK), .Q_N(n5490) );
	dfxbp_1 DFF_879_Q_reg( .D(n4816), .CLK(CLK), .Q_N(n5321) );
	dfxtp_1 DFF_1000_Q_reg( .D(n4), .CLK(CLK), .Q(g1833) );
	dfxbp_1 DFF_1001_Q_reg( .D(n4009), .CLK(CLK), .Q(n10079) );
	dfxtp_1 DFF_1145_Q_reg( .D(n4116), .CLK(CLK), .Q(g1910) );
	dfxbp_1 DFF_883_Q_reg( .D(n4820), .CLK(CLK), .Q_N(n5489) );
	dfxbp_1 DFF_882_Q_reg( .D(n4819), .CLK(CLK), .Q_N(n5320) );
	dfxbp_1 DFF_905_Q_reg( .D(n4842), .CLK(CLK), .Q(n9968), .Q_N(n5602) );
	dfxtp_1 DFF_904_Q_reg( .D(n4841), .CLK(CLK), .Q(n7385) );
	dfxtp_1 DFF_903_Q_reg( .D(n4840), .CLK(CLK), .Q(n7386) );
	dfxbp_1 DFF_976_Q_reg( .D(n4895), .CLK(CLK), .Q_N(n5562) );
	dfxbp_1 DFF_975_Q_reg( .D(n4894), .CLK(CLK), .Q(n9792), .Q_N(n5620) );
	dfxtp_1 DFF_974_Q_reg( .D(n4893), .CLK(CLK), .Q(n7629) );
	dfxbp_1 DFF_979_Q_reg( .D(n4898), .CLK(CLK), .Q_N(n5550) );
	dfxbp_1 DFF_978_Q_reg( .D(n4897), .CLK(CLK), .Q_N(n5340) );
	dfxtp_1 DFF_977_Q_reg( .D(n4896), .CLK(CLK), .Q(n7633) );
	dfxbp_1 DFF_1082_Q_reg( .D(n4938), .CLK(CLK), .Q(n9929), .Q_N(n5650) );
	dfxtp_1 DFF_1081_Q_reg( .D(n4937), .CLK(CLK), .Q(n7452) );
	dfxbp_1 DFF_1080_Q_reg( .D(n4936), .CLK(CLK), .Q_N(n5418) );
	dfxtp_1 DFF_1103_Q_reg( .D(n4041), .CLK(CLK), .Q(g1938) );
	dfxbp_1 DFF_103_Q_reg( .D(n4304), .CLK(CLK), .Q_N(n5500) );
	dfxbp_1 DFF_102_Q_reg( .D(n4303), .CLK(CLK), .Q(n9932), .Q_N(n5580) );
	dfxbp_1 DFF_101_Q_reg( .D(n4302), .CLK(CLK), .Q_N(n5389) );
	dfxtp_1 DFF_982_Q_reg( .D(n4901), .CLK(CLK), .Q(n7312) );
	dfxtp_1 DFF_981_Q_reg( .D(n4900), .CLK(CLK), .Q(n7311) );
	dfxbp_1 DFF_896_Q_reg( .D(n4833), .CLK(CLK), .Q(n9987), .Q_N(n5676) );
	dfxtp_1 DFF_895_Q_reg( .D(n4832), .CLK(CLK), .Q(n7392) );
	dfxtp_1 DFF_894_Q_reg( .D(n4831), .CLK(CLK), .Q(n7394) );
	dfxtp_1 DFF_973_Q_reg( .D(n4892), .CLK(CLK), .Q(n7338) );
	dfxtp_1 DFF_972_Q_reg( .D(n4891), .CLK(CLK), .Q(n7337) );
	dfxbp_1 DFF_967_Q_reg( .D(n4886), .CLK(CLK), .Q(n9986), .Q_N(n5668) );
	dfxbp_1 DFF_966_Q_reg( .D(n4885), .CLK(CLK), .Q(n9793), .Q_N(n5669) );
	dfxtp_1 DFF_965_Q_reg( .D(n4884), .CLK(CLK), .Q(n7625) );
	dfxbp_1 DFF_970_Q_reg( .D(n4889), .CLK(CLK), .Q_N(n5551) );
	dfxbp_1 DFF_969_Q_reg( .D(n4888), .CLK(CLK), .Q_N(n5341) );
	dfxtp_1 DFF_968_Q_reg( .D(n4887), .CLK(CLK), .Q(n7623) );
	dfxbp_1 DFF_1091_Q_reg( .D(n4944), .CLK(CLK), .Q(n9926), .Q_N(n5648) );
	dfxtp_1 DFF_1090_Q_reg( .D(n4943), .CLK(CLK), .Q(n7460) );
	dfxbp_1 DFF_1089_Q_reg( .D(n4942), .CLK(CLK), .Q_N(n5419) );
	dfxtp_1 DFF_1101_Q_reg( .D(n4040), .CLK(CLK), .Q(g1929) );
	dfxbp_1 DFF_127_Q_reg( .D(n4328), .CLK(CLK), .Q_N(n5385) );
	dfxbp_1 DFF_126_Q_reg( .D(n4327), .CLK(CLK), .Q_N(n5310) );
	dfxbp_1 DFF_125_Q_reg( .D(n4326), .CLK(CLK), .Q(n9981), .Q_N(n5581) );
	dfxtp_1 DFF_997_Q_reg( .D(n4916), .CLK(CLK), .Q(n7376) );
	dfxtp_1 DFF_996_Q_reg( .D(n4915), .CLK(CLK), .Q(n7375) );
	dfxtp_1 DFF_988_Q_reg( .D(n4907), .CLK(CLK), .Q(n7582) );
	dfxtp_1 DFF_987_Q_reg( .D(n4906), .CLK(CLK), .Q(n7581) );
	dfxbp_1 DFF_986_Q_reg( .D(n4905), .CLK(CLK), .Q(n9935), .Q_N(n5618) );
	dfxtp_1 DFF_908_Q_reg( .D(n4845), .CLK(CLK), .Q(n7681) );
	dfxbp_1 DFF_907_Q_reg( .D(n4844), .CLK(CLK), .Q_N(n5396) );
	dfxbp_1 DFF_906_Q_reg( .D(n4843), .CLK(CLK), .Q(n9939), .Q_N(n5704) );
	dfxtp_1 DFF_923_Q_reg( .D(n4860), .CLK(CLK), .Q(n7679) );
	dfxbp_1 DFF_922_Q_reg( .D(n4859), .CLK(CLK), .Q(n9943), .Q_N(n5725) );
	dfxbp_1 DFF_921_Q_reg( .D(n4858), .CLK(CLK), .Q(n9944), .Q_N(n5683) );
	dfxtp_1 DFF_985_Q_reg( .D(n4904), .CLK(CLK), .Q(n7578) );
	dfxtp_1 DFF_984_Q_reg( .D(n4903), .CLK(CLK), .Q(n7577) );
	dfxbp_1 DFF_983_Q_reg( .D(n4902), .CLK(CLK), .Q(n9933), .Q_N(n5619) );
	dfxtp_1 DFF_914_Q_reg( .D(n4851), .CLK(CLK), .Q(n7686) );
	dfxbp_1 DFF_913_Q_reg( .D(n4850), .CLK(CLK), .Q_N(n5532) );
	dfxbp_1 DFF_912_Q_reg( .D(n4849), .CLK(CLK), .Q(n9949), .Q_N(n5702) );
	dfxtp_1 DFF_917_Q_reg( .D(n4854), .CLK(CLK), .Q(n7678) );
	dfxbp_1 DFF_916_Q_reg( .D(n4853), .CLK(CLK), .Q_N(n5531) );
	dfxbp_1 DFF_915_Q_reg( .D(n4852), .CLK(CLK), .Q(n9947), .Q_N(n5701) );
	dfxtp_1 DFF_920_Q_reg( .D(n4857), .CLK(CLK), .Q(n7683) );
	dfxbp_1 DFF_919_Q_reg( .D(n4856), .CLK(CLK), .Q(n9940), .Q_N(n5726) );
	dfxbp_1 DFF_918_Q_reg( .D(n4855), .CLK(CLK), .Q(n9941), .Q_N(n5684) );
	dfxtp_1 DFF_926_Q_reg( .D(n4863), .CLK(CLK), .Q(n7680) );
	dfxbp_1 DFF_925_Q_reg( .D(n4862), .CLK(CLK), .Q_N(n5534) );
	dfxbp_1 DFF_924_Q_reg( .D(n4861), .CLK(CLK), .Q(n9942), .Q_N(n5700) );
	dfxtp_1 DFF_929_Q_reg( .D(n4866), .CLK(CLK), .Q(n7685) );
	dfxbp_1 DFF_928_Q_reg( .D(n4865), .CLK(CLK), .Q(n9945), .Q_N(n5724) );
	dfxbp_1 DFF_927_Q_reg( .D(n4864), .CLK(CLK), .Q(n9946), .Q_N(n5682) );
	dfxtp_1 DFF_932_Q_reg( .D(n4869), .CLK(CLK), .Q(n7687) );
	dfxbp_1 DFF_931_Q_reg( .D(n4868), .CLK(CLK), .Q_N(n5533) );
	dfxbp_1 DFF_930_Q_reg( .D(n4867), .CLK(CLK), .Q(n9948), .Q_N(n5699) );
	dfxtp_1 DFF_935_Q_reg( .D(n4872), .CLK(CLK), .Q(n7684) );
	dfxbp_1 DFF_934_Q_reg( .D(n4871), .CLK(CLK), .Q(n9937), .Q_N(n5723) );
	dfxbp_1 DFF_933_Q_reg( .D(n4870), .CLK(CLK), .Q(n9938), .Q_N(n5681) );
	dfxtp_1 DFF_991_Q_reg( .D(n4910), .CLK(CLK), .Q(n7580) );
	dfxtp_1 DFF_990_Q_reg( .D(n4909), .CLK(CLK), .Q(n7579) );
	dfxbp_1 DFF_989_Q_reg( .D(n4908), .CLK(CLK), .Q(n9934), .Q_N(n5617) );
	dfxtp_1 DFF_994_Q_reg( .D(n4913), .CLK(CLK), .Q(n7329) );
	dfxtp_1 DFF_993_Q_reg( .D(n4912), .CLK(CLK), .Q(n7330) );
	dfxtp_1 DFF_911_Q_reg( .D(n4848), .CLK(CLK), .Q(n7682) );
	dfxbp_1 DFF_910_Q_reg( .D(n4847), .CLK(CLK), .Q_N(n5530) );
	dfxbp_1 DFF_909_Q_reg( .D(n4846), .CLK(CLK), .Q(n9936), .Q_N(n5703) );
	dfxtp_1 DFF_1094_Q_reg( .D(n4089), .CLK(CLK), .Q(g1852) );
	dfxtp_1 DFF_1075_Q_reg( .D(n27), .CLK(CLK), .Q(g1948) );
	dfxbp_1 DFF_1076_Q_reg( .D(n4935), .CLK(CLK), .Q_N(n15642) );
	dfxtp_1 DFF_1093_Q_reg( .D(n4088), .CLK(CLK), .Q(g1849) );
	dfxtp_1 DFF_1073_Q_reg( .D(n26), .CLK(CLK), .Q(g1946) );
	dfxtp_1 DFF_1074_Q_reg( .D(n4164), .CLK(CLK), .Q(g1947) );
	dfxtp_1 DFF_1092_Q_reg( .D(n4087), .CLK(CLK), .Q(g1846) );
	dfxtp_1 DFF_1071_Q_reg( .D(n25), .CLK(CLK), .Q(g1954) );
	dfxbp_1 DFF_1072_Q_reg( .D(n4934), .CLK(CLK), .Q(n9925) );
	dfxtp_1 DFF_1095_Q_reg( .D(n4038), .CLK(CLK), .Q(g1908) );
	dfxtp_1 DFF_1096_Q_reg( .D(n3985), .CLK(CLK), .Q(g1915) );
	dfxtp_1 DFF_1097_Q_reg( .D(n4143), .CLK(CLK), .Q(g1922) );
	dfxtp_1 DFF_961_Q_reg( .D(n4253), .CLK(CLK), .Q(g1757) );
	dfxtp_1 DFF_1045_Q_reg( .D(n17), .CLK(CLK), .Q(g1763) );
	dfxbp_1 DFF_1046_Q_reg( .D(n4925), .CLK(CLK), .Q_N(n15048) );
	dfxtp_1 DFF_960_Q_reg( .D(n4252), .CLK(CLK), .Q(g1754) );
	dfxtp_1 DFF_1043_Q_reg( .D(n16), .CLK(CLK), .Q(g1761) );
	dfxbp_1 DFF_1044_Q_reg( .D(n4924), .CLK(CLK), .Q_N(n15049) );
	dfxtp_1 DFF_958_Q_reg( .D(n4251), .CLK(CLK), .Q(g1742) );
	dfxtp_1 DFF_1039_Q_reg( .D(n15), .CLK(CLK), .Q(g1748) );
	dfxbp_1 DFF_1040_Q_reg( .D(n4923), .CLK(CLK), .Q_N(n15051) );
	dfxtp_1 DFF_957_Q_reg( .D(n4250), .CLK(CLK), .Q(g1739) );
	dfxtp_1 DFF_1037_Q_reg( .D(n14), .CLK(CLK), .Q(g1746) );
	dfxbp_1 DFF_1038_Q_reg( .D(n4922), .CLK(CLK), .Q_N(n15053) );
	dfxtp_1 DFF_964_Q_reg( .D(n4255), .CLK(CLK), .Q(g1772) );
	dfxtp_1 DFF_1051_Q_reg( .D(n19), .CLK(CLK), .Q(g1778) );
	dfxbp_1 DFF_1052_Q_reg( .D(n4927), .CLK(CLK), .Q_N(n15044) );
	dfxtp_1 DFF_963_Q_reg( .D(n4254), .CLK(CLK), .Q(g1769) );
	dfxtp_1 DFF_1049_Q_reg( .D(n18), .CLK(CLK), .Q(g1776) );
	dfxbp_1 DFF_1050_Q_reg( .D(n4926), .CLK(CLK), .Q_N(n15045) );
	dfxtp_1 DFF_1047_Q_reg( .D(n3983), .CLK(CLK), .Q(g1768) );
	dfxtp_1 DFF_1048_Q_reg( .D(n4163), .CLK(CLK), .Q(g1775) );
	dfxtp_1 DFF_1035_Q_reg( .D(n3981), .CLK(CLK), .Q(g1738) );
	dfxtp_1 DFF_1036_Q_reg( .D(n4140), .CLK(CLK), .Q(g1745) );
	dfxtp_1 DFF_1041_Q_reg( .D(n3982), .CLK(CLK), .Q(g1753) );
	dfxtp_1 DFF_1042_Q_reg( .D(n4162), .CLK(CLK), .Q(g1760) );
	dfxtp_1 DFF_955_Q_reg( .D(n4249), .CLK(CLK), .Q(g1727) );
	dfxtp_1 DFF_1033_Q_reg( .D(n13), .CLK(CLK), .Q(g1733) );
	dfxbp_1 DFF_1034_Q_reg( .D(n4921), .CLK(CLK), .Q_N(n15046) );
	dfxtp_1 DFF_954_Q_reg( .D(n4248), .CLK(CLK), .Q(g1724) );
	dfxtp_1 DFF_1031_Q_reg( .D(n12), .CLK(CLK), .Q(g1731) );
	dfxbp_1 DFF_1032_Q_reg( .D(n4920), .CLK(CLK), .Q_N(n15047) );
	dfxtp_1 DFF_1029_Q_reg( .D(n3980), .CLK(CLK), .Q(g1723) );
	dfxtp_1 DFF_1030_Q_reg( .D(n4161), .CLK(CLK), .Q(g1730) );
	dfxtp_1 DFF_1085_Q_reg( .D(n4086), .CLK(CLK), .Q(g1842) );
	dfxtp_1 DFF_1069_Q_reg( .D(n24), .CLK(CLK), .Q(g1952) );
	dfxbp_1 DFF_1070_Q_reg( .D(n4933), .CLK(CLK), .Q_N(n15629) );
	dfxtp_1 DFF_1084_Q_reg( .D(n4085), .CLK(CLK), .Q(g1839) );
	dfxtp_1 DFF_1067_Q_reg( .D(n23), .CLK(CLK), .Q(g1950) );
	dfxtp_1 DFF_1068_Q_reg( .D(n4142), .CLK(CLK), .Q(g1951) );
	dfxtp_1 DFF_1083_Q_reg( .D(n4084), .CLK(CLK), .Q(g1836) );
	dfxtp_1 DFF_1065_Q_reg( .D(n22), .CLK(CLK), .Q(g1944) );
	dfxbp_1 DFF_1066_Q_reg( .D(n4932), .CLK(CLK), .Q(n9930) );
	dfxtp_1 DFF_1062_Q_reg( .D(n4037), .CLK(CLK), .Q(g1893) );
	dfxtp_1 DFF_1063_Q_reg( .D(n3984), .CLK(CLK), .Q(g1903) );
	dfxtp_1 DFF_1064_Q_reg( .D(n4141), .CLK(CLK), .Q(g1904) );
	dfxtp_1 DFF_1028_Q_reg( .D(n4160), .CLK(CLK), .Q(g1679) );
	dfxbp_1 DFF_1017_Q_reg( .D(n4919), .CLK(CLK), .Q(n9966), .Q_N(n5674) );
	dfxtp_1 DFF_1367_Q_reg( .D(n5149), .CLK(CLK), .Q(n7632) );
	dfxbp_1 DFF_1088_Q_reg( .D(n4941), .CLK(CLK), .Q(n9928), .Q_N(n5649) );
	dfxtp_1 DFF_1087_Q_reg( .D(n4940), .CLK(CLK), .Q(n7455) );
	dfxbp_1 DFF_1086_Q_reg( .D(n4939), .CLK(CLK), .Q_N(n5420) );
	dfxtp_1 DFF_1098_Q_reg( .D(n4039), .CLK(CLK), .Q(g1923) );
	dfxbp_1 DFF_1099_Q_reg( .D(n4945), .CLK(CLK), .Q_N(n14880) );
	dfxbp_1 DFF_1100_Q_reg( .D(n4946), .CLK(CLK), .Q(n9922) );
	dfxbp_1 DFF_115_Q_reg( .D(n4316), .CLK(CLK), .Q_N(n5387) );
	dfxbp_1 DFF_114_Q_reg( .D(n4315), .CLK(CLK), .Q(n9915), .Q_N(n5577) );
	dfxbp_1 DFF_113_Q_reg( .D(n4314), .CLK(CLK), .Q_N(n5388) );
	dfxbp_1 DFF_1450_Q_reg( .D(n34), .CLK(CLK), .Q(n9913) );
	dfxbp_1 DFF_118_Q_reg( .D(n4319), .CLK(CLK), .Q(n9982), .Q_N(n5583) );
	dfxbp_1 DFF_117_Q_reg( .D(n4318), .CLK(CLK), .Q(n9912), .Q_N(n5584) );
	dfxbp_1 DFF_116_Q_reg( .D(n4317), .CLK(CLK), .Q_N(n5312) );
	dfxbp_1 DFF_156_Q_reg( .D(n4337), .CLK(CLK), .Q(n9888) );
	dfxbp_1 DFF_142_Q_reg( .D(n4337), .CLK(CLK), .Q(n9887) );
	dfxbp_1 DFF_136_Q_reg( .D(n4340), .CLK(CLK), .Q(n10055), .Q_N(n5483) );
	dfxbp_1 DFF_158_Q_reg( .D(n4339), .CLK(CLK), .Q(n9979) );
	dfxbp_1 DFF_157_Q_reg( .D(n4338), .CLK(CLK), .Q(n9980), .Q_N(n5382) );
	dfxbp_1 DFF_138_Q_reg( .D(n4338), .CLK(CLK), .Q(n10054), .Q_N(n5352) );
	dfxbp_1 DFF_152_Q_reg( .D(n4336), .CLK(CLK), .Q_N(n15211) );
	dfxtp_1 DFF_132_Q_reg( .D(n4336), .CLK(CLK), .Q(g3194) );
	dfxbp_1 DFF_131_Q_reg( .D(n4332), .CLK(CLK), .Q(n10057) );
	dfxbp_1 DFF_146_Q_reg( .D(n4333), .CLK(CLK), .Q(n10053) );
	dfxbp_1 DFF_150_Q_reg( .D(n4334), .CLK(CLK), .Q_N(n15214) );
	dfxtp_1 DFF_134_Q_reg( .D(n4334), .CLK(CLK), .Q(g3198) );
	dfxbp_1 DFF_143_Q_reg( .D(n4334), .CLK(CLK), .Q_N(n15217) );
	dfxbp_1 DFF_151_Q_reg( .D(n4335), .CLK(CLK), .Q_N(n15213) );
	dfxbp_1 DFF_133_Q_reg( .D(n4335), .CLK(CLK), .Q(n10056), .Q_N(n5739) );
	dfxtp_1 DFF_144_Q_reg( .D(n4098), .CLK(CLK), .Q(g3125) );
	dfxbp_1 DFF_145_Q_reg( .D(n4336), .CLK(CLK), .Q_N(n15212) );
	dfxbp_1 DFF_153_Q_reg( .D(n4338), .CLK(CLK), .Q_N(n5567) );
	dfxtp_1 DFF_91_Q_reg( .D(n4071), .CLK(CLK), .Q(g2878) );
	dfxtp_1 DFF_1364_Q_reg( .D(n57), .CLK(CLK), .Q(g2365) );
	dfxbp_1 DFF_1365_Q_reg( .D(n5147), .CLK(CLK), .Q_N(DFF_1503_D) );
	dfxbp_1 DFF_1503_Q_reg( .D(n69), .CLK(CLK), .Q(n9863) );
	dfxbp_1 DFF_1502_Q_reg( .D(n5205), .CLK(CLK), .Q(n9872) );
	dfxtp_1 DFF_63_Q_reg( .D(n4061), .CLK(CLK), .Q(g7519) );
	dfxtp_1 DFF_64_Q_reg( .D(n148), .CLK(CLK), .Q(g2873) );
	dfxtp_1 DFF_664_Q_reg( .D(n3973), .CLK(CLK), .Q(g977) );
	dfxbp_1 DFF_665_Q_reg( .D(n4688), .CLK(CLK), .Q_N(DFF_803_D) );
	dfxbp_1 DFF_803_Q_reg( .D(n167), .CLK(CLK), .Q(n9865) );
	dfxbp_1 DFF_802_Q_reg( .D(n4747), .CLK(CLK), .Q(n9866) );
	dfxtp_1 DFF_81_Q_reg( .D(n4070), .CLK(CLK), .Q(g8096) );
	dfxtp_1 DFF_82_Q_reg( .D(n168), .CLK(CLK), .Q(g2857) );
	dfxtp_1 DFF_314_Q_reg( .D(n3966), .CLK(CLK), .Q(g290) );
	dfxbp_1 DFF_315_Q_reg( .D(n4458), .CLK(CLK), .Q_N(DFF_453_D) );
	dfxbp_1 DFF_453_Q_reg( .D(n119), .CLK(CLK), .Q(n9868) );
	dfxbp_1 DFF_452_Q_reg( .D(n4518), .CLK(CLK), .Q(n9869) );
	dfxtp_1 DFF_46_Q_reg( .D(n4052), .CLK(CLK), .Q(g2877) );
	dfxtp_1 DFF_1014_Q_reg( .D(n11), .CLK(CLK), .Q(g1671) );
	dfxbp_1 DFF_1015_Q_reg( .D(n4917), .CLK(CLK), .Q_N(DFF_1153_D) );
	dfxbp_1 DFF_1153_Q_reg( .D(n33), .CLK(CLK), .Q(n9864) );
	dfxbp_1 DFF_1152_Q_reg( .D(n4977), .CLK(CLK), .Q(n9914) );
	dfxbp_1 DFF_770_Q_reg( .D(n4733), .CLK(CLK), .Q_N(n5406) );
	dfxbp_1 DFF_772_Q_reg( .D(n4735), .CLK(CLK), .Q(n9798), .Q_N(n5623) );
	dfxbp_1 DFF_771_Q_reg( .D(n4734), .CLK(CLK), .Q(n9799), .Q_N(n5597) );
	dfxbp_1 DFF_767_Q_reg( .D(n4730), .CLK(CLK), .Q_N(n5407) );
	dfxbp_1 DFF_769_Q_reg( .D(n4732), .CLK(CLK), .Q(n9800), .Q_N(n5624) );
	dfxbp_1 DFF_768_Q_reg( .D(n4731), .CLK(CLK), .Q(n9801), .Q_N(n5598) );
	dfxbp_1 DFF_778_Q_reg( .D(n4741), .CLK(CLK), .Q_N(n5556) );
	dfxbp_1 DFF_777_Q_reg( .D(n4740), .CLK(CLK), .Q_N(n5346) );
	dfxtp_1 DFF_776_Q_reg( .D(n4739), .CLK(CLK), .Q(n7663) );
	dfxbp_1 DFF_783_Q_reg( .D(n4745), .CLK(CLK), .Q_N(n15150) );
	dfxbp_1 DFF_755_Q_reg( .D(n4718), .CLK(CLK), .Q_N(n5509) );
	dfxtp_1 DFF_763_Q_reg( .D(n4726), .CLK(CLK), .Q(n7359) );
	dfxtp_1 DFF_762_Q_reg( .D(n4725), .CLK(CLK), .Q(n7360) );
	dfxbp_1 DFF_761_Q_reg( .D(n4724), .CLK(CLK), .Q_N(n5511) );
	dfxtp_1 DFF_760_Q_reg( .D(n4723), .CLK(CLK), .Q(n7361) );
	dfxtp_1 DFF_759_Q_reg( .D(n4722), .CLK(CLK), .Q(n7362) );
	dfxbp_1 DFF_758_Q_reg( .D(n4721), .CLK(CLK), .Q_N(n5510) );
	dfxtp_1 DFF_766_Q_reg( .D(n4729), .CLK(CLK), .Q(n7365) );
	dfxtp_1 DFF_765_Q_reg( .D(n4728), .CLK(CLK), .Q(n7366) );
	dfxbp_1 DFF_764_Q_reg( .D(n4727), .CLK(CLK), .Q_N(n5512) );
	dfxbp_1 DFF_775_Q_reg( .D(n4738), .CLK(CLK), .Q_N(n5555) );
	dfxbp_1 DFF_774_Q_reg( .D(n4737), .CLK(CLK), .Q_N(n5345) );
	dfxtp_1 DFF_773_Q_reg( .D(n4736), .CLK(CLK), .Q(n7662) );
	dfxbp_1 DFF_851_Q_reg( .D(n4791), .CLK(CLK), .Q(n9988), .Q_N(n5621) );
	dfxtp_1 DFF_850_Q_reg( .D(n4790), .CLK(CLK), .Q(n7449) );
	dfxbp_1 DFF_849_Q_reg( .D(n4789), .CLK(CLK), .Q_N(n5392) );
	dfxbp_1 DFF_781_Q_reg( .D(n4744), .CLK(CLK), .Q_N(n5564) );
	dfxbp_1 DFF_780_Q_reg( .D(n4743), .CLK(CLK), .Q(n9802), .Q_N(n5727) );
	dfxtp_1 DFF_779_Q_reg( .D(n4742), .CLK(CLK), .Q(n7638) );
	dfxtp_1 DFF_757_Q_reg( .D(n4720), .CLK(CLK), .Q(n7363) );
	dfxtp_1 DFF_756_Q_reg( .D(n4719), .CLK(CLK), .Q(n7364) );
	dfxbp_1 DFF_854_Q_reg( .D(n4794), .CLK(CLK), .Q(n9867), .Q_N(n5572) );
	dfxtp_1 DFF_853_Q_reg( .D(n4793), .CLK(CLK), .Q(n7534) );
	dfxbp_1 DFF_852_Q_reg( .D(n4792), .CLK(CLK), .Q_N(n5458) );
	dfxbp_1 DFF_420_Q_reg( .D(n4504), .CLK(CLK), .Q_N(n5408) );
	dfxbp_1 DFF_422_Q_reg( .D(n4506), .CLK(CLK), .Q(n9829), .Q_N(n5627) );
	dfxbp_1 DFF_421_Q_reg( .D(n4505), .CLK(CLK), .Q(n9830), .Q_N(n5599) );
	dfxbp_1 DFF_417_Q_reg( .D(n4501), .CLK(CLK), .Q_N(n5409) );
	dfxbp_1 DFF_419_Q_reg( .D(n4503), .CLK(CLK), .Q(n9831), .Q_N(n5628) );
	dfxbp_1 DFF_418_Q_reg( .D(n4502), .CLK(CLK), .Q(n9832), .Q_N(n5600) );
	dfxbp_1 DFF_428_Q_reg( .D(n4512), .CLK(CLK), .Q_N(n5558) );
	dfxbp_1 DFF_427_Q_reg( .D(n4511), .CLK(CLK), .Q_N(n5348) );
	dfxtp_1 DFF_426_Q_reg( .D(n4510), .CLK(CLK), .Q(n7665) );
	dfxbp_1 DFF_433_Q_reg( .D(n4516), .CLK(CLK), .Q_N(n15423) );
	dfxtp_1 DFF_442_Q_reg( .D(n4049), .CLK(CLK), .Q(g16297) );
	dfxbp_1 DFF_443_Q_reg( .D(n4517), .CLK(CLK), .Q(n9976), .Q_N(n5518) );
	dfxtp_1 DFF_498_Q_reg( .D(n4559), .CLK(CLK), .Q(n7549) );
	dfxtp_1 DFF_495_Q_reg( .D(n4556), .CLK(CLK), .Q(n7551) );
	dfxtp_1 DFF_492_Q_reg( .D(n4553), .CLK(CLK), .Q(n7560) );
	dfxtp_1 DFF_489_Q_reg( .D(n4550), .CLK(CLK), .Q(n7562) );
	dfxtp_1 DFF_486_Q_reg( .D(n4547), .CLK(CLK), .Q(n7564) );
	dfxtp_1 DFF_483_Q_reg( .D(n4544), .CLK(CLK), .Q(n7566) );
	dfxtp_1 DFF_480_Q_reg( .D(n4541), .CLK(CLK), .Q(n7557) );
	dfxtp_1 DFF_477_Q_reg( .D(n4538), .CLK(CLK), .Q(n7553) );
	dfxtp_1 DFF_474_Q_reg( .D(n4535), .CLK(CLK), .Q(n7555) );
	dfxtp_1 DFF_471_Q_reg( .D(n4532), .CLK(CLK), .Q(n7568) );
	dfxtp_1 DFF_510_Q_reg( .D(n4571), .CLK(CLK), .Q(n7318) );
	dfxtp_1 DFF_497_Q_reg( .D(n4558), .CLK(CLK), .Q(n7548) );
	dfxtp_1 DFF_494_Q_reg( .D(n4555), .CLK(CLK), .Q(n7550) );
	dfxtp_1 DFF_491_Q_reg( .D(n4552), .CLK(CLK), .Q(n7559) );
	dfxtp_1 DFF_488_Q_reg( .D(n4549), .CLK(CLK), .Q(n7561) );
	dfxtp_1 DFF_485_Q_reg( .D(n4546), .CLK(CLK), .Q(n7563) );
	dfxtp_1 DFF_482_Q_reg( .D(n4543), .CLK(CLK), .Q(n7565) );
	dfxtp_1 DFF_479_Q_reg( .D(n4540), .CLK(CLK), .Q(n7556) );
	dfxtp_1 DFF_476_Q_reg( .D(n4537), .CLK(CLK), .Q(n7552) );
	dfxtp_1 DFF_473_Q_reg( .D(n4534), .CLK(CLK), .Q(n7554) );
	dfxtp_1 DFF_470_Q_reg( .D(n4531), .CLK(CLK), .Q(n7567) );
	dfxbp_1 DFF_509_Q_reg( .D(n4570), .CLK(CLK), .Q_N(n5336) );
	dfxbp_1 DFF_496_Q_reg( .D(n4557), .CLK(CLK), .Q_N(n5463) );
	dfxbp_1 DFF_493_Q_reg( .D(n4554), .CLK(CLK), .Q_N(n5466) );
	dfxbp_1 DFF_490_Q_reg( .D(n4551), .CLK(CLK), .Q_N(n5472) );
	dfxbp_1 DFF_487_Q_reg( .D(n4548), .CLK(CLK), .Q_N(n5469) );
	dfxbp_1 DFF_484_Q_reg( .D(n4545), .CLK(CLK), .Q_N(n5470) );
	dfxbp_1 DFF_481_Q_reg( .D(n4542), .CLK(CLK), .Q_N(n5467) );
	dfxbp_1 DFF_478_Q_reg( .D(n4539), .CLK(CLK), .Q_N(n5465) );
	dfxbp_1 DFF_475_Q_reg( .D(n4536), .CLK(CLK), .Q(n10036), .Q_N(n5626) );
	dfxbp_1 DFF_472_Q_reg( .D(n4533), .CLK(CLK), .Q_N(n5464) );
	dfxbp_1 DFF_469_Q_reg( .D(n4530), .CLK(CLK), .Q_N(n5471) );
	dfxbp_1 DFF_508_Q_reg( .D(n4569), .CLK(CLK), .Q_N(n5545) );
	dfxbp_1 DFF_793_Q_reg( .D(n4746), .CLK(CLK), .Q(n9971), .Q_N(n5517) );
	dfxtp_1 DFF_848_Q_reg( .D(n4788), .CLK(CLK), .Q(n7525) );
	dfxtp_1 DFF_845_Q_reg( .D(n4785), .CLK(CLK), .Q(n7527) );
	dfxtp_1 DFF_842_Q_reg( .D(n4782), .CLK(CLK), .Q(n7536) );
	dfxtp_1 DFF_839_Q_reg( .D(n4779), .CLK(CLK), .Q(n7538) );
	dfxtp_1 DFF_836_Q_reg( .D(n4776), .CLK(CLK), .Q(n7540) );
	dfxtp_1 DFF_833_Q_reg( .D(n4773), .CLK(CLK), .Q(n7542) );
	dfxtp_1 DFF_830_Q_reg( .D(n4770), .CLK(CLK), .Q(n7533) );
	dfxtp_1 DFF_827_Q_reg( .D(n4767), .CLK(CLK), .Q(n7529) );
	dfxtp_1 DFF_824_Q_reg( .D(n4764), .CLK(CLK), .Q(n7531) );
	dfxtp_1 DFF_821_Q_reg( .D(n4761), .CLK(CLK), .Q(n7544) );
	dfxtp_1 DFF_860_Q_reg( .D(n4800), .CLK(CLK), .Q(n7317) );
	dfxtp_1 DFF_847_Q_reg( .D(n4787), .CLK(CLK), .Q(n7524) );
	dfxtp_1 DFF_844_Q_reg( .D(n4784), .CLK(CLK), .Q(n7526) );
	dfxtp_1 DFF_841_Q_reg( .D(n4781), .CLK(CLK), .Q(n7535) );
	dfxtp_1 DFF_838_Q_reg( .D(n4778), .CLK(CLK), .Q(n7537) );
	dfxtp_1 DFF_835_Q_reg( .D(n4775), .CLK(CLK), .Q(n7539) );
	dfxtp_1 DFF_832_Q_reg( .D(n4772), .CLK(CLK), .Q(n7541) );
	dfxtp_1 DFF_829_Q_reg( .D(n4769), .CLK(CLK), .Q(n7532) );
	dfxtp_1 DFF_826_Q_reg( .D(n4766), .CLK(CLK), .Q(n7528) );
	dfxtp_1 DFF_823_Q_reg( .D(n4763), .CLK(CLK), .Q(n7530) );
	dfxtp_1 DFF_820_Q_reg( .D(n4760), .CLK(CLK), .Q(n7543) );
	dfxbp_1 DFF_859_Q_reg( .D(n4799), .CLK(CLK), .Q_N(n5335) );
	dfxbp_1 DFF_846_Q_reg( .D(n4786), .CLK(CLK), .Q_N(n5453) );
	dfxbp_1 DFF_843_Q_reg( .D(n4783), .CLK(CLK), .Q_N(n5456) );
	dfxbp_1 DFF_840_Q_reg( .D(n4780), .CLK(CLK), .Q_N(n5462) );
	dfxbp_1 DFF_837_Q_reg( .D(n4777), .CLK(CLK), .Q_N(n5459) );
	dfxbp_1 DFF_834_Q_reg( .D(n4774), .CLK(CLK), .Q_N(n5460) );
	dfxbp_1 DFF_831_Q_reg( .D(n4771), .CLK(CLK), .Q_N(n5457) );
	dfxbp_1 DFF_828_Q_reg( .D(n4768), .CLK(CLK), .Q_N(n5455) );
	dfxbp_1 DFF_825_Q_reg( .D(n4765), .CLK(CLK), .Q(n10035), .Q_N(n5622) );
	dfxbp_1 DFF_822_Q_reg( .D(n4762), .CLK(CLK), .Q_N(n5454) );
	dfxbp_1 DFF_819_Q_reg( .D(n4759), .CLK(CLK), .Q_N(n5461) );
	dfxtp_1 DFF_857_Q_reg( .D(n4797), .CLK(CLK), .Q(n7523) );
	dfxtp_1 DFF_856_Q_reg( .D(n4796), .CLK(CLK), .Q(n7546) );
	dfxtp_1 DFF_855_Q_reg( .D(n4795), .CLK(CLK), .Q(n7545) );
	dfxbp_1 DFF_858_Q_reg( .D(n4798), .CLK(CLK), .Q_N(n5544) );
	dfxtp_1 DFF_1581_Q_reg( .D(n4186), .CLK(CLK), .Q(g3061) );
	dfxtp_1 DFF_1580_Q_reg( .D(n4185), .CLK(CLK), .Q(g3060) );
	dfxtp_1 DFF_1579_Q_reg( .D(n4184), .CLK(CLK), .Q(g3059) );
	dfxtp_1 DFF_1578_Q_reg( .D(n4183), .CLK(CLK), .Q(g3058) );
	dfxtp_1 DFF_1577_Q_reg( .D(n4182), .CLK(CLK), .Q(g3057) );
	dfxtp_1 DFF_1576_Q_reg( .D(n4181), .CLK(CLK), .Q(g3056) );
	dfxtp_1 DFF_1575_Q_reg( .D(n4180), .CLK(CLK), .Q(g3055) );
	dfxtp_1 DFF_1574_Q_reg( .D(n4179), .CLK(CLK), .Q(g3053) );
	dfxtp_1 DFF_1573_Q_reg( .D(n4178), .CLK(CLK), .Q(g3052) );
	dfxbp_1 DFF_405_Q_reg( .D(n4489), .CLK(CLK), .Q_N(n5513) );
	dfxtp_1 DFF_413_Q_reg( .D(n4497), .CLK(CLK), .Q(n7367) );
	dfxtp_1 DFF_412_Q_reg( .D(n4496), .CLK(CLK), .Q(n7368) );
	dfxbp_1 DFF_411_Q_reg( .D(n4495), .CLK(CLK), .Q_N(n5515) );
	dfxtp_1 DFF_410_Q_reg( .D(n4494), .CLK(CLK), .Q(n7369) );
	dfxtp_1 DFF_409_Q_reg( .D(n4493), .CLK(CLK), .Q(n7370) );
	dfxbp_1 DFF_408_Q_reg( .D(n4492), .CLK(CLK), .Q_N(n5514) );
	dfxtp_1 DFF_416_Q_reg( .D(n4500), .CLK(CLK), .Q(n7373) );
	dfxtp_1 DFF_415_Q_reg( .D(n4499), .CLK(CLK), .Q(n7374) );
	dfxbp_1 DFF_414_Q_reg( .D(n4498), .CLK(CLK), .Q_N(n5516) );
	dfxbp_1 DFF_425_Q_reg( .D(n4509), .CLK(CLK), .Q_N(n5557) );
	dfxbp_1 DFF_424_Q_reg( .D(n4508), .CLK(CLK), .Q_N(n5347) );
	dfxtp_1 DFF_423_Q_reg( .D(n4507), .CLK(CLK), .Q(n7664) );
	dfxbp_1 DFF_501_Q_reg( .D(n4562), .CLK(CLK), .Q(n10010), .Q_N(n5625) );
	dfxtp_1 DFF_500_Q_reg( .D(n4561), .CLK(CLK), .Q(n7450) );
	dfxbp_1 DFF_499_Q_reg( .D(n4560), .CLK(CLK), .Q_N(n5393) );
	dfxbp_1 DFF_431_Q_reg( .D(n4515), .CLK(CLK), .Q_N(n5565) );
	dfxbp_1 DFF_430_Q_reg( .D(n4514), .CLK(CLK), .Q(n9833), .Q_N(n5730) );
	dfxtp_1 DFF_429_Q_reg( .D(n4513), .CLK(CLK), .Q(n7639) );
	dfxtp_1 DFF_407_Q_reg( .D(n4491), .CLK(CLK), .Q(n7371) );
	dfxtp_1 DFF_406_Q_reg( .D(n4490), .CLK(CLK), .Q(n7372) );
	dfxbp_1 DFF_504_Q_reg( .D(n4565), .CLK(CLK), .Q(n9870), .Q_N(n5573) );
	dfxtp_1 DFF_503_Q_reg( .D(n4564), .CLK(CLK), .Q(n7558) );
	dfxbp_1 DFF_502_Q_reg( .D(n4563), .CLK(CLK), .Q_N(n5468) );
	dfxtp_1 DFF_507_Q_reg( .D(n4568), .CLK(CLK), .Q(n7547) );
	dfxtp_1 DFF_506_Q_reg( .D(n4567), .CLK(CLK), .Q(n7570) );
	dfxtp_1 DFF_505_Q_reg( .D(n4566), .CLK(CLK), .Q(n7569) );
	dfxtp_1 DFF_1571_Q_reg( .D(n4176), .CLK(CLK), .Q(g3050) );
	dfxtp_1 DFF_1569_Q_reg( .D(n4174), .CLK(CLK), .Q(g3048) );
	dfxtp_1 DFF_1565_Q_reg( .D(n4170), .CLK(CLK), .Q(g3044) );
	dfxtp_1 DFF_1567_Q_reg( .D(n4172), .CLK(CLK), .Q(g3046) );
	dfxtp_1 DFF_1566_Q_reg( .D(n4171), .CLK(CLK), .Q(g3045) );
	dfxtp_1 DFF_1564_Q_reg( .D(n4169), .CLK(CLK), .Q(g3043) );
	dfxtp_1 DFF_1570_Q_reg( .D(n4175), .CLK(CLK), .Q(g3049) );
	dfxtp_1 DFF_1572_Q_reg( .D(n4177), .CLK(CLK), .Q(g3051) );
	dfxtp_1 DFF_1568_Q_reg( .D(n4173), .CLK(CLK), .Q(g3047) );
	dfxbp_1 DFF_1470_Q_reg( .D(n5193), .CLK(CLK), .Q_N(n5402) );
	dfxbp_1 DFF_1472_Q_reg( .D(n5195), .CLK(CLK), .Q(n9873), .Q_N(n5607) );
	dfxbp_1 DFF_1471_Q_reg( .D(n5194), .CLK(CLK), .Q(n9874), .Q_N(n5593) );
	dfxbp_1 DFF_1467_Q_reg( .D(n5190), .CLK(CLK), .Q_N(n5403) );
	dfxbp_1 DFF_1469_Q_reg( .D(n5192), .CLK(CLK), .Q(n9875), .Q_N(n5608) );
	dfxbp_1 DFF_1468_Q_reg( .D(n5191), .CLK(CLK), .Q(n9876), .Q_N(n5594) );
	dfxbp_1 DFF_1478_Q_reg( .D(n5201), .CLK(CLK), .Q_N(n5561) );
	dfxbp_1 DFF_1477_Q_reg( .D(n5200), .CLK(CLK), .Q_N(n5351) );
	dfxtp_1 DFF_1476_Q_reg( .D(n5199), .CLK(CLK), .Q(n7659) );
	dfxtp_1 DFF_1483_Q_reg( .D(n4148), .CLK(CLK), .Q(g2581) );
	dfxbp_1 DFF_1455_Q_reg( .D(n5178), .CLK(CLK), .Q_N(n5501) );
	dfxtp_1 DFF_1463_Q_reg( .D(n5186), .CLK(CLK), .Q(n7343) );
	dfxtp_1 DFF_1462_Q_reg( .D(n5185), .CLK(CLK), .Q(n7344) );
	dfxbp_1 DFF_1461_Q_reg( .D(n5184), .CLK(CLK), .Q_N(n5503) );
	dfxtp_1 DFF_1460_Q_reg( .D(n5183), .CLK(CLK), .Q(n7345) );
	dfxtp_1 DFF_1459_Q_reg( .D(n5182), .CLK(CLK), .Q(n7346) );
	dfxbp_1 DFF_1458_Q_reg( .D(n5181), .CLK(CLK), .Q_N(n5502) );
	dfxtp_1 DFF_1466_Q_reg( .D(n5189), .CLK(CLK), .Q(n7349) );
	dfxtp_1 DFF_1465_Q_reg( .D(n5188), .CLK(CLK), .Q(n7350) );
	dfxbp_1 DFF_1464_Q_reg( .D(n5187), .CLK(CLK), .Q_N(n5504) );
	dfxbp_1 DFF_1475_Q_reg( .D(n5198), .CLK(CLK), .Q_N(n5560) );
	dfxbp_1 DFF_1474_Q_reg( .D(n5197), .CLK(CLK), .Q_N(n5350) );
	dfxtp_1 DFF_1473_Q_reg( .D(n5196), .CLK(CLK), .Q(n7658) );
	dfxbp_1 DFF_1551_Q_reg( .D(n5249), .CLK(CLK), .Q(n10037), .Q_N(n5605) );
	dfxtp_1 DFF_1550_Q_reg( .D(n5248), .CLK(CLK), .Q(n7447) );
	dfxbp_1 DFF_1549_Q_reg( .D(n5247), .CLK(CLK), .Q_N(n5390) );
	dfxbp_1 DFF_1481_Q_reg( .D(n5204), .CLK(CLK), .Q_N(n5566) );
	dfxbp_1 DFF_1480_Q_reg( .D(n5203), .CLK(CLK), .Q(n9877), .Q_N(n5719) );
	dfxtp_1 DFF_1479_Q_reg( .D(n5202), .CLK(CLK), .Q(n7636) );
	dfxtp_1 DFF_1457_Q_reg( .D(n5180), .CLK(CLK), .Q(n7347) );
	dfxtp_1 DFF_1456_Q_reg( .D(n5179), .CLK(CLK), .Q(n7348) );
	dfxbp_1 DFF_1554_Q_reg( .D(n5252), .CLK(CLK), .Q(n9871), .Q_N(n5570) );
	dfxtp_1 DFF_1553_Q_reg( .D(n5251), .CLK(CLK), .Q(n7486) );
	dfxbp_1 DFF_1552_Q_reg( .D(n5250), .CLK(CLK), .Q_N(n5448) );
	dfxbp_1 DFF_1120_Q_reg( .D(n4963), .CLK(CLK), .Q_N(n5404) );
	dfxbp_1 DFF_1122_Q_reg( .D(n4965), .CLK(CLK), .Q(n9917), .Q_N(n5615) );
	dfxbp_1 DFF_1121_Q_reg( .D(n4964), .CLK(CLK), .Q(n9918), .Q_N(n5595) );
	dfxbp_1 DFF_1117_Q_reg( .D(n4960), .CLK(CLK), .Q_N(n5405) );
	dfxbp_1 DFF_1119_Q_reg( .D(n4962), .CLK(CLK), .Q(n9919), .Q_N(n5616) );
	dfxbp_1 DFF_1118_Q_reg( .D(n4961), .CLK(CLK), .Q(n9920), .Q_N(n5596) );
	dfxbp_1 DFF_1128_Q_reg( .D(n4971), .CLK(CLK), .Q_N(n5559) );
	dfxbp_1 DFF_1127_Q_reg( .D(n4970), .CLK(CLK), .Q_N(n5349) );
	dfxtp_1 DFF_1126_Q_reg( .D(n4969), .CLK(CLK), .Q(n7661) );
	dfxbp_1 DFF_1204_Q_reg( .D(n5024), .CLK(CLK), .Q(n9911), .Q_N(n5571) );
	dfxtp_1 DFF_1203_Q_reg( .D(n5023), .CLK(CLK), .Q(n7510) );
	dfxbp_1 DFF_1202_Q_reg( .D(n5022), .CLK(CLK), .Q_N(n5478) );
	dfxbp_1 DFF_1133_Q_reg( .D(n4975), .CLK(CLK), .Q_N(n15018) );
	dfxbp_1 DFF_1143_Q_reg( .D(n4976), .CLK(CLK), .Q(n9964) );
	dfxtp_1 DFF_1198_Q_reg( .D(n5018), .CLK(CLK), .Q(n7501) );
	dfxtp_1 DFF_1195_Q_reg( .D(n5015), .CLK(CLK), .Q(n7503) );
	dfxtp_1 DFF_1192_Q_reg( .D(n5012), .CLK(CLK), .Q(n7512) );
	dfxtp_1 DFF_1189_Q_reg( .D(n5009), .CLK(CLK), .Q(n7514) );
	dfxtp_1 DFF_1186_Q_reg( .D(n5006), .CLK(CLK), .Q(n7516) );
	dfxtp_1 DFF_1183_Q_reg( .D(n5003), .CLK(CLK), .Q(n7518) );
	dfxtp_1 DFF_1180_Q_reg( .D(n5000), .CLK(CLK), .Q(n7509) );
	dfxtp_1 DFF_1177_Q_reg( .D(n4997), .CLK(CLK), .Q(n7505) );
	dfxtp_1 DFF_1174_Q_reg( .D(n4994), .CLK(CLK), .Q(n7507) );
	dfxtp_1 DFF_1171_Q_reg( .D(n4991), .CLK(CLK), .Q(n7520) );
	dfxtp_1 DFF_1210_Q_reg( .D(n5030), .CLK(CLK), .Q(n7316) );
	dfxtp_1 DFF_1197_Q_reg( .D(n5017), .CLK(CLK), .Q(n7500) );
	dfxtp_1 DFF_1194_Q_reg( .D(n5014), .CLK(CLK), .Q(n7502) );
	dfxtp_1 DFF_1191_Q_reg( .D(n5011), .CLK(CLK), .Q(n7511) );
	dfxtp_1 DFF_1188_Q_reg( .D(n5008), .CLK(CLK), .Q(n7513) );
	dfxtp_1 DFF_1185_Q_reg( .D(n5005), .CLK(CLK), .Q(n7515) );
	dfxtp_1 DFF_1182_Q_reg( .D(n5002), .CLK(CLK), .Q(n7517) );
	dfxtp_1 DFF_1179_Q_reg( .D(n4999), .CLK(CLK), .Q(n7508) );
	dfxtp_1 DFF_1176_Q_reg( .D(n4996), .CLK(CLK), .Q(n7504) );
	dfxtp_1 DFF_1173_Q_reg( .D(n4993), .CLK(CLK), .Q(n7506) );
	dfxtp_1 DFF_1170_Q_reg( .D(n4990), .CLK(CLK), .Q(n7519) );
	dfxbp_1 DFF_1209_Q_reg( .D(n5029), .CLK(CLK), .Q_N(n5337) );
	dfxbp_1 DFF_1196_Q_reg( .D(n5016), .CLK(CLK), .Q_N(n5473) );
	dfxbp_1 DFF_1193_Q_reg( .D(n5013), .CLK(CLK), .Q_N(n5476) );
	dfxbp_1 DFF_1190_Q_reg( .D(n5010), .CLK(CLK), .Q_N(n5482) );
	dfxbp_1 DFF_1187_Q_reg( .D(n5007), .CLK(CLK), .Q_N(n5479) );
	dfxbp_1 DFF_1184_Q_reg( .D(n5004), .CLK(CLK), .Q_N(n5480) );
	dfxbp_1 DFF_1181_Q_reg( .D(n5001), .CLK(CLK), .Q_N(n5477) );
	dfxbp_1 DFF_1178_Q_reg( .D(n4998), .CLK(CLK), .Q_N(n5475) );
	dfxbp_1 DFF_1175_Q_reg( .D(n4995), .CLK(CLK), .Q(n10069), .Q_N(n5614) );
	dfxbp_1 DFF_1172_Q_reg( .D(n4992), .CLK(CLK), .Q_N(n5474) );
	dfxbp_1 DFF_1169_Q_reg( .D(n4989), .CLK(CLK), .Q_N(n5481) );
	dfxbp_1 DFF_1208_Q_reg( .D(n5028), .CLK(CLK), .Q_N(n5546) );
	dfxtp_1 DFF_1588_Q_reg( .D(n4192), .CLK(CLK), .Q(g3068) );
	dfxtp_1 DFF_1586_Q_reg( .D(n4149), .CLK(CLK), .Q(g3066) );
	dfxtp_1 DFF_1492_Q_reg( .D(n4096), .CLK(CLK), .Q(g16437) );
	dfxbp_1 DFF_1493_Q_reg( .D(n68), .CLK(CLK), .Q(n9959), .Q_N(n5574) );
	dfxtp_1 DFF_1548_Q_reg( .D(n5246), .CLK(CLK), .Q(n7477) );
	dfxtp_1 DFF_1545_Q_reg( .D(n5243), .CLK(CLK), .Q(n7479) );
	dfxtp_1 DFF_1542_Q_reg( .D(n5240), .CLK(CLK), .Q(n7488) );
	dfxtp_1 DFF_1539_Q_reg( .D(n5237), .CLK(CLK), .Q(n7490) );
	dfxtp_1 DFF_1536_Q_reg( .D(n5234), .CLK(CLK), .Q(n7492) );
	dfxtp_1 DFF_1533_Q_reg( .D(n5231), .CLK(CLK), .Q(n7494) );
	dfxtp_1 DFF_1530_Q_reg( .D(n5228), .CLK(CLK), .Q(n7485) );
	dfxtp_1 DFF_1527_Q_reg( .D(n5225), .CLK(CLK), .Q(n7481) );
	dfxtp_1 DFF_1524_Q_reg( .D(n5222), .CLK(CLK), .Q(n7483) );
	dfxtp_1 DFF_1521_Q_reg( .D(n5219), .CLK(CLK), .Q(n7496) );
	dfxtp_1 DFF_1560_Q_reg( .D(n5258), .CLK(CLK), .Q(n7315) );
	dfxtp_1 DFF_1547_Q_reg( .D(n5245), .CLK(CLK), .Q(n7476) );
	dfxtp_1 DFF_1544_Q_reg( .D(n5242), .CLK(CLK), .Q(n7478) );
	dfxtp_1 DFF_1541_Q_reg( .D(n5239), .CLK(CLK), .Q(n7487) );
	dfxtp_1 DFF_1538_Q_reg( .D(n5236), .CLK(CLK), .Q(n7489) );
	dfxtp_1 DFF_1535_Q_reg( .D(n5233), .CLK(CLK), .Q(n7491) );
	dfxtp_1 DFF_1532_Q_reg( .D(n5230), .CLK(CLK), .Q(n7493) );
	dfxtp_1 DFF_1529_Q_reg( .D(n5227), .CLK(CLK), .Q(n7484) );
	dfxtp_1 DFF_1526_Q_reg( .D(n5224), .CLK(CLK), .Q(n7480) );
	dfxtp_1 DFF_1523_Q_reg( .D(n5221), .CLK(CLK), .Q(n7482) );
	dfxtp_1 DFF_1520_Q_reg( .D(n5218), .CLK(CLK), .Q(n7495) );
	dfxbp_1 DFF_1559_Q_reg( .D(n5257), .CLK(CLK), .Q_N(n5334) );
	dfxbp_1 DFF_1546_Q_reg( .D(n5244), .CLK(CLK), .Q_N(n5443) );
	dfxbp_1 DFF_1543_Q_reg( .D(n5241), .CLK(CLK), .Q_N(n5446) );
	dfxbp_1 DFF_1540_Q_reg( .D(n5238), .CLK(CLK), .Q_N(n5452) );
	dfxbp_1 DFF_1537_Q_reg( .D(n5235), .CLK(CLK), .Q_N(n5450) );
	dfxbp_1 DFF_1534_Q_reg( .D(n5232), .CLK(CLK), .Q_N(n5449) );
	dfxbp_1 DFF_1531_Q_reg( .D(n5229), .CLK(CLK), .Q_N(n5447) );
	dfxbp_1 DFF_1528_Q_reg( .D(n5226), .CLK(CLK), .Q_N(n5445) );
	dfxbp_1 DFF_1525_Q_reg( .D(n5223), .CLK(CLK), .Q(n10039), .Q_N(n5606) );
	dfxbp_1 DFF_1522_Q_reg( .D(n5220), .CLK(CLK), .Q_N(n5444) );
	dfxbp_1 DFF_1519_Q_reg( .D(n5217), .CLK(CLK), .Q_N(n5451) );
	dfxtp_1 DFF_1557_Q_reg( .D(n5255), .CLK(CLK), .Q(n7475) );
	dfxtp_1 DFF_1556_Q_reg( .D(n5254), .CLK(CLK), .Q(n7498) );
	dfxtp_1 DFF_1555_Q_reg( .D(n5253), .CLK(CLK), .Q(n7497) );
	dfxbp_1 DFF_1558_Q_reg( .D(n5256), .CLK(CLK), .Q_N(n5543) );
	dfxtp_1 DFF_1598_Q_reg( .D(n4202), .CLK(CLK), .Q(g3078) );
	dfxtp_1 DFF_1596_Q_reg( .D(n4200), .CLK(CLK), .Q(g3076) );
	dfxtp_1 DFF_1597_Q_reg( .D(n4201), .CLK(CLK), .Q(g3077) );
	dfxtp_1 DFF_1599_Q_reg( .D(n4203), .CLK(CLK), .Q(g2997) );
	dfxtp_1 DFF_1633_Q_reg( .D(n89), .CLK(CLK), .Q(g2990) );
	dfxtp_1 DFF_1595_Q_reg( .D(n4199), .CLK(CLK), .Q(g3075) );
	dfxtp_1 DFF_1629_Q_reg( .D(n85), .CLK(CLK), .Q(g8263) );
	dfxtp_1 DFF_1594_Q_reg( .D(n4198), .CLK(CLK), .Q(g3074) );
	dfxtp_1 DFF_1591_Q_reg( .D(n4195), .CLK(CLK), .Q(g3071) );
	dfxtp_1 DFF_1593_Q_reg( .D(n4197), .CLK(CLK), .Q(g3073) );
	dfxtp_1 DFF_1592_Q_reg( .D(n4196), .CLK(CLK), .Q(g3072) );
	dfxbp_1 DFF_1634_Q_reg( .D(n5274), .CLK(CLK), .Q_N(n15173) );
	dfxbp_1 DFF_1105_Q_reg( .D(n4948), .CLK(CLK), .Q_N(n5505) );
	dfxtp_1 DFF_1113_Q_reg( .D(n4956), .CLK(CLK), .Q(n7351) );
	dfxtp_1 DFF_1112_Q_reg( .D(n4955), .CLK(CLK), .Q(n7352) );
	dfxbp_1 DFF_1111_Q_reg( .D(n4954), .CLK(CLK), .Q_N(n5507) );
	dfxtp_1 DFF_1110_Q_reg( .D(n4953), .CLK(CLK), .Q(n7353) );
	dfxtp_1 DFF_1109_Q_reg( .D(n4952), .CLK(CLK), .Q(n7354) );
	dfxbp_1 DFF_1108_Q_reg( .D(n4951), .CLK(CLK), .Q_N(n5506) );
	dfxtp_1 DFF_1116_Q_reg( .D(n4959), .CLK(CLK), .Q(n7357) );
	dfxtp_1 DFF_1115_Q_reg( .D(n4958), .CLK(CLK), .Q(n7358) );
	dfxbp_1 DFF_1114_Q_reg( .D(n4957), .CLK(CLK), .Q_N(n5508) );
	dfxbp_1 DFF_1125_Q_reg( .D(n4968), .CLK(CLK), .Q_N(n5554) );
	dfxbp_1 DFF_1124_Q_reg( .D(n4967), .CLK(CLK), .Q_N(n5344) );
	dfxtp_1 DFF_1123_Q_reg( .D(n4966), .CLK(CLK), .Q(n7660) );
	dfxbp_1 DFF_1131_Q_reg( .D(n4974), .CLK(CLK), .Q_N(n5563) );
	dfxbp_1 DFF_1130_Q_reg( .D(n4973), .CLK(CLK), .Q(n9921), .Q_N(n5722) );
	dfxtp_1 DFF_1129_Q_reg( .D(n4972), .CLK(CLK), .Q(n7637) );
	dfxbp_1 DFF_1201_Q_reg( .D(n5021), .CLK(CLK), .Q(n10067), .Q_N(n5613) );
	dfxtp_1 DFF_1200_Q_reg( .D(n5020), .CLK(CLK), .Q(n7448) );
	dfxbp_1 DFF_1199_Q_reg( .D(n5019), .CLK(CLK), .Q_N(n5391) );
	dfxtp_1 DFF_1207_Q_reg( .D(n5027), .CLK(CLK), .Q(n7499) );
	dfxtp_1 DFF_1206_Q_reg( .D(n5026), .CLK(CLK), .Q(n7522) );
	dfxtp_1 DFF_1205_Q_reg( .D(n5025), .CLK(CLK), .Q(n7521) );
	dfxtp_1 DFF_1584_Q_reg( .D(n4189), .CLK(CLK), .Q(g3064) );
	dfxtp_1 DFF_1582_Q_reg( .D(n4187), .CLK(CLK), .Q(g3062) );
	dfxtp_1 DFF_1585_Q_reg( .D(n4190), .CLK(CLK), .Q(g3065) );
	dfxtp_1 DFF_1583_Q_reg( .D(n4188), .CLK(CLK), .Q(g3063) );
	dfxtp_1 DFF_1589_Q_reg( .D(n4193), .CLK(CLK), .Q(g3069) );
	dfxtp_1 DFF_1590_Q_reg( .D(n4194), .CLK(CLK), .Q(g3070) );
	dfxtp_1 DFF_1622_Q_reg( .D(n80), .CLK(CLK), .Q(g3083) );
	dfxtp_1 DFF_1587_Q_reg( .D(n4191), .CLK(CLK), .Q(g3067) );
	dfxtp_1 DFF_1619_Q_reg( .D(n77), .CLK(CLK), .Q(g8269) );
	dfxbp_1 DFF_1624_Q_reg( .D(n5273), .CLK(CLK), .Q_N(n15172) );
	dfxtp_1 DFF_1107_Q_reg( .D(n4950), .CLK(CLK), .Q(n7355) );
	dfxtp_1 DFF_1106_Q_reg( .D(n4949), .CLK(CLK), .Q(n7356) );
	dfxbp_1 DFF_139_Q_reg( .D(n4341), .CLK(CLK), .Q(n9883) );
	dfxbp_1 DFF_140_Q_reg( .D(n4339), .CLK(CLK), .Q_N(n15165) );
	dfxbp_1 DFF_154_Q_reg( .D(n4339), .CLK(CLK), .Q_N(n5414) );
	dfxtp_1 DFF_1635_Q_reg( .D(n4025), .CLK(CLK), .Q(g8258) );
	dfxtp_1 DFF_1623_Q_reg( .D(n4024), .CLK(CLK), .Q(g8267) );
	dfxbp_1 DFF_155_Q_reg( .D(n4340), .CLK(CLK), .Q_N(n15162) );
	dfxtp_1 DFF_141_Q_reg( .D(n4097), .CLK(CLK), .Q(g3128) );
	dfxbp_1 DFF_149_Q_reg( .D(n4337), .CLK(CLK), .Q(n9886) );
	dfxtp_1 DFF_34_Q_reg( .D(n4291), .CLK(CLK), .Q(n7602) );
	dfxtp_1 DFF_33_Q_reg( .D(n4290), .CLK(CLK), .Q(n7597) );
	dfxtp_1 DFF_32_Q_reg( .D(n4289), .CLK(CLK), .Q(n7604) );
	dfxtp_1 DFF_27_Q_reg( .D(n4285), .CLK(CLK), .Q(n7608) );
	dfxtp_1 DFF_25_Q_reg( .D(n4283), .CLK(CLK), .Q(n7600) );
	dfxtp_1 DFF_24_Q_reg( .D(n4282), .CLK(CLK), .Q(n7606) );
	dfxtp_1 DFF_92_Q_reg( .D(n4231), .CLK(CLK), .Q(g8106) );
	dfxtp_1 DFF_93_Q_reg( .D(n4209), .CLK(CLK), .Q(g8030) );
	dfxtp_1 DFF_354_Q_reg( .D(n4204), .CLK(CLK), .Q(g5648) );
	dfxtp_1 DFF_1054_Q_reg( .D(n4206), .CLK(CLK), .Q(g5738) );
	dfxtp_1 DFF_1404_Q_reg( .D(n4207), .CLK(CLK), .Q(g5796) );
	dfxtp_1 DFF_704_Q_reg( .D(n4205), .CLK(CLK), .Q(g5686) );
	dfxtp_1 DFF_178_Q_reg( .D(n4356), .CLK(CLK), .Q(n7325) );
	dfxtp_1 DFF_280_Q_reg( .D(n4440), .CLK(CLK), .Q(n7715) );
	dfxtp_1 DFF_271_Q_reg( .D(n4431), .CLK(CLK), .Q(n7735) );
	dfxtp_1 DFF_295_Q_reg( .D(n4455), .CLK(CLK), .Q(n7740) );
	dfxtp_1 DFF_528_Q_reg( .D(n4586), .CLK(CLK), .Q(n7323) );
	dfxtp_1 DFF_630_Q_reg( .D(n4670), .CLK(CLK), .Q(n7736) );
	dfxtp_1 DFF_622_Q_reg( .D(n4662), .CLK(CLK), .Q(n7734) );
	dfxtp_1 DFF_646_Q_reg( .D(n4686), .CLK(CLK), .Q(n7739) );
	dfxtp_1 DFF_1345_Q_reg( .D(n5144), .CLK(CLK), .Q(n7737) );
	dfxtp_1 DFF_1330_Q_reg( .D(n5129), .CLK(CLK), .Q(n7713) );
	dfxtp_1 DFF_1321_Q_reg( .D(n5120), .CLK(CLK), .Q(n7732) );
	dfxtp_1 DFF_872_Q_reg( .D(n4809), .CLK(CLK), .Q(n7324) );
	dfxtp_1 DFF_980_Q_reg( .D(n4899), .CLK(CLK), .Q(n7714) );
	dfxtp_1 DFF_971_Q_reg( .D(n4890), .CLK(CLK), .Q(n7733) );
	dfxtp_1 DFF_995_Q_reg( .D(n4914), .CLK(CLK), .Q(n7738) );
	dfxtp_1 DFF_792_Q_reg( .D(n4229), .CLK(CLK), .Q(g16355) );
	dfxtp_1 DFF_1142_Q_reg( .D(n4230), .CLK(CLK), .Q(g16399) );
	dfxtp_1 DFF_1620_Q_reg( .D(n78), .CLK(CLK), .Q(g8270) );
	dfxtp_1 DFF_1631_Q_reg( .D(n87), .CLK(CLK), .Q(g8261) );
	dfxtp_1 DFF_1628_Q_reg( .D(n84), .CLK(CLK), .Q(g8262) );
	dfxtp_1 DFF_1621_Q_reg( .D(n79), .CLK(CLK), .Q(g8271) );
	dfxtp_1 DFF_1618_Q_reg( .D(n76), .CLK(CLK), .Q(g8268) );
	dfxtp_1 DFF_1632_Q_reg( .D(n88), .CLK(CLK), .Q(g8259) );
	dfxtp_1 DFF_1626_Q_reg( .D(n82), .CLK(CLK), .Q(g8265) );
	dfxtp_1 DFF_1617_Q_reg( .D(n75), .CLK(CLK), .Q(g8272) );
	dfxtp_1 DFF_1615_Q_reg( .D(n73), .CLK(CLK), .Q(g8274) );
	dfxtp_1 DFF_1630_Q_reg( .D(n86), .CLK(CLK), .Q(g8260) );
	dfxtp_1 DFF_1625_Q_reg( .D(n81), .CLK(CLK), .Q(g8266) );
	dfxtp_1 DFF_1627_Q_reg( .D(n83), .CLK(CLK), .Q(g8264) );
	dfxtp_1 DFF_1616_Q_reg( .D(n74), .CLK(CLK), .Q(g8273) );
	dfxtp_1 DFF_1614_Q_reg( .D(n72), .CLK(CLK), .Q(g8275) );
	dfxtp_1 DFF_3_Q_reg( .D(n4048), .CLK(CLK), .Q(g2950) );
	dfxtp_1 DFF_184_Q_reg( .D(n4362), .CLK(CLK), .Q(n7613) );
	dfxtp_1 DFF_534_Q_reg( .D(n4592), .CLK(CLK), .Q(n7612) );
	dfxtp_1 DFF_175_Q_reg( .D(n4353), .CLK(CLK), .Q(n7616) );
	dfxtp_1 DFF_525_Q_reg( .D(n4583), .CLK(CLK), .Q(n7615) );
	dfxtp_1 DFF_887_Q_reg( .D(n4824), .CLK(CLK), .Q(n7610) );
	dfxtp_1 DFF_1237_Q_reg( .D(n5054), .CLK(CLK), .Q(n7609) );
	dfxtp_1 DFF_875_Q_reg( .D(n4812), .CLK(CLK), .Q(n7614) );
	dfxtp_1 DFF_881_Q_reg( .D(n4818), .CLK(CLK), .Q(n7322) );
	dfxtp_1 DFF_884_Q_reg( .D(n4821), .CLK(CLK), .Q(n7611) );
	dfxtp_1 DFF_253_Q_reg( .D(n4213), .CLK(CLK), .Q(g354) );
	dfxtp_1 DFF_259_Q_reg( .D(n4215), .CLK(CLK), .Q(g384) );
	dfxtp_1 DFF_256_Q_reg( .D(n4214), .CLK(CLK), .Q(g369) );
	dfxtp_1 DFF_262_Q_reg( .D(n4216), .CLK(CLK), .Q(g398) );
	dfxtp_1 DFF_1303_Q_reg( .D(n4225), .CLK(CLK), .Q(g2429) );
	dfxtp_1 DFF_1309_Q_reg( .D(n4227), .CLK(CLK), .Q(g2459) );
	dfxtp_1 DFF_1306_Q_reg( .D(n4226), .CLK(CLK), .Q(g2444) );
	dfxtp_1 DFF_1312_Q_reg( .D(n4228), .CLK(CLK), .Q(g2473) );
	dfxtp_1 DFF_953_Q_reg( .D(n4221), .CLK(CLK), .Q(g1735) );
	dfxtp_1 DFF_959_Q_reg( .D(n4223), .CLK(CLK), .Q(g1765) );
	dfxtp_1 DFF_956_Q_reg( .D(n4222), .CLK(CLK), .Q(g1750) );
	dfxtp_1 DFF_962_Q_reg( .D(n4224), .CLK(CLK), .Q(g1779) );
	dfxtp_1 DFF_316_Q_reg( .D(n4459), .CLK(CLK), .Q(n7745) );
	dfxtp_1 DFF_432_Q_reg( .D(n35), .CLK(CLK), .Q(n7744) );
	dfxtp_1 DFF_666_Q_reg( .D(n4689), .CLK(CLK), .Q(n7742) );
	dfxtp_1 DFF_782_Q_reg( .D(n44), .CLK(CLK), .Q(n7741) );
	dfxtp_1 DFF_1366_Q_reg( .D(n5148), .CLK(CLK), .Q(n7743) );
	dfxtp_1 DFF_1482_Q_reg( .D(n47), .CLK(CLK), .Q(n7725) );
	dfxtp_1 DFF_1016_Q_reg( .D(n4918), .CLK(CLK), .Q(n7731) );
	dfxtp_1 DFF_1132_Q_reg( .D(n32), .CLK(CLK), .Q(n7730) );
	dfxtp_1 DFF_80_Q_reg( .D(n166), .CLK(CLK), .Q(n7594) );
	dfxtp_1 DFF_90_Q_reg( .D(n5290), .CLK(CLK), .Q(n7242) );
	dfxtp_1 DFF_610_Q_reg( .D(n4219), .CLK(CLK), .Q(g1060) );
	dfxtp_1 DFF_607_Q_reg( .D(n4218), .CLK(CLK), .Q(g1045) );
	dfxtp_1 DFF_613_Q_reg( .D(n4220), .CLK(CLK), .Q(g1075) );
	dfxtp_1 DFF_604_Q_reg( .D(n4217), .CLK(CLK), .Q(g1030) );
	dfxtp_1 DFF_458_Q_reg( .D(n4520), .CLK(CLK), .Q(n7278) );
	dfxtp_1 DFF_1158_Q_reg( .D(n4979), .CLK(CLK), .Q(n7276) );
	dfxtp_1 DFF_1508_Q_reg( .D(n5207), .CLK(CLK), .Q(n7275) );
	dfxtp_1 DFF_808_Q_reg( .D(n4749), .CLK(CLK), .Q(n7277) );
	dfxtp_1 DFF_292_Q_reg( .D(n4452), .CLK(CLK), .Q(n7729) );
	dfxtp_1 DFF_643_Q_reg( .D(n4683), .CLK(CLK), .Q(n7728) );
	dfxtp_1 DFF_1342_Q_reg( .D(n5141), .CLK(CLK), .Q(n7726) );
	dfxtp_1 DFF_992_Q_reg( .D(n4911), .CLK(CLK), .Q(n7727) );
	dfxtp_1 DFF_754_Q_reg( .D(n4717), .CLK(CLK), .Q(n7288) );
	dfxtp_1 DFF_1454_Q_reg( .D(n5177), .CLK(CLK), .Q(n7294) );
	dfxtp_1 DFF_1104_Q_reg( .D(n4947), .CLK(CLK), .Q(n7289) );
	dfxtp_1 DFF_148_Q_reg( .D(n4340), .CLK(CLK), .Q(n7723) );
	dfxtp_1 DFF_147_Q_reg( .D(n4339), .CLK(CLK), .Q(n7724) );
	dfxtp_1 DFF_1613_Q_reg( .D(n5303), .CLK(CLK), .Q(n7255) );
	dfxtp_1 DFF_19_Q_reg( .D(n3957), .CLK(CLK), .Q(n7587) );
	dfxtp_1 DFF_1060_Q_reg( .D(n4930), .CLK(CLK), .Q(n7291) );
	dfxtp_1 DFF_37_Q_reg( .D(n4294), .CLK(CLK), .Q(n7603) );
	dfxtp_1 DFF_36_Q_reg( .D(n4293), .CLK(CLK), .Q(n7595) );
	dfxtp_1 DFF_35_Q_reg( .D(n4292), .CLK(CLK), .Q(n7601) );
	dfxtp_1 DFF_30_Q_reg( .D(n4287), .CLK(CLK), .Q(n7596) );
	dfxtp_1 DFF_26_Q_reg( .D(n4284), .CLK(CLK), .Q(n7607) );
	dfxtp_1 DFF_23_Q_reg( .D(n4281), .CLK(CLK), .Q(n7599) );
	dfxtp_1 DFF_22_Q_reg( .D(n4280), .CLK(CLK), .Q(n7605) );
	dfxtp_1 DFF_21_Q_reg( .D(n4279), .CLK(CLK), .Q(n7598) );
	dfxtp_1 DFF_1289_Q_reg( .D(n5106), .CLK(CLK), .Q(n7709) );
	dfxtp_1 DFF_1294_Q_reg( .D(n5111), .CLK(CLK), .Q(n7307) );
	dfxtp_1 DFF_939_Q_reg( .D(n4876), .CLK(CLK), .Q(n7710) );
	dfxtp_1 DFF_944_Q_reg( .D(n4881), .CLK(CLK), .Q(n7308) );
	dfxtp_1 DFF_239_Q_reg( .D(n4417), .CLK(CLK), .Q(n7712) );
	dfxtp_1 DFF_244_Q_reg( .D(n4422), .CLK(CLK), .Q(n7306) );
	dfxtp_1 DFF_589_Q_reg( .D(n4647), .CLK(CLK), .Q(n7711) );
	dfxtp_1 DFF_594_Q_reg( .D(n4652), .CLK(CLK), .Q(n7305) );
	dfxtp_1 DFF_8_Q_reg( .D(n4269), .CLK(CLK), .Q(n7321) );
	dfxtp_1 DFF_1411_Q_reg( .D(n5162), .CLK(CLK), .Q(n7588) );
	dfxtp_1 DFF_159_Q_reg( .D(n4340), .CLK(CLK), .Q(n7722) );
	dfxtp_1 DFF_70_Q_reg( .D(n151), .CLK(CLK), .Q(n7269) );
	dfxtp_1 DFF_68_Q_reg( .D(n150), .CLK(CLK), .Q(n7241) );
	dfxtp_1 DFF_52_Q_reg( .D(n127), .CLK(CLK), .Q(n7270) );
	dfxtp_1 DFF_710_Q_reg( .D(n4701), .CLK(CLK), .Q(n7292) );
	dfxtp_1 DFF_360_Q_reg( .D(n4472), .CLK(CLK), .Q(n7293) );
	dfxtp_1 DFF_85_Q_reg( .D(n5285), .CLK(CLK), .Q(n7261) );
	dfxtp_1 DFF_40_Q_reg( .D(n5277), .CLK(CLK), .Q(n7221) );
	dfxtp_1 DFF_1609_Q_reg( .D(n5270), .CLK(CLK), .Q(n7704) );
	dfxtp_1 DFF_937_Q_reg( .D(n4874), .CLK(CLK), .Q(n7700) );
	dfxtp_1 DFF_587_Q_reg( .D(n4645), .CLK(CLK), .Q(n7701) );
	dfxtp_1 DFF_13_Q_reg( .D(n4274), .CLK(CLK), .Q(n7703) );
	dfxtp_1 DFF_727_Q_reg( .D(n4131), .CLK(CLK), .Q(g7961) );
	dfxtp_1 DFF_728_Q_reg( .D(n161), .CLK(CLK), .Q(g8007) );
	dfxtp_1 DFF_729_Q_reg( .D(n162), .CLK(CLK), .Q(n7258) );
	dfxtp_1 DFF_1427_Q_reg( .D(n4131), .CLK(CLK), .Q(g8087) );
	dfxtp_1 DFF_1428_Q_reg( .D(n66), .CLK(CLK), .Q(g8167) );
	dfxtp_1 DFF_1429_Q_reg( .D(n67), .CLK(CLK), .Q(n7260) );
	dfxtp_1 DFF_1077_Q_reg( .D(n4131), .CLK(CLK), .Q(g8012) );
	dfxtp_1 DFF_1078_Q_reg( .D(n28), .CLK(CLK), .Q(g8082) );
	dfxtp_1 DFF_1079_Q_reg( .D(n29), .CLK(CLK), .Q(n7257) );
	dfxtp_1 DFF_377_Q_reg( .D(n4131), .CLK(CLK), .Q(g7909) );
	dfxtp_1 DFF_378_Q_reg( .D(n117), .CLK(CLK), .Q(g7956) );
	dfxtp_1 DFF_379_Q_reg( .D(n118), .CLK(CLK), .Q(n7259) );
	dfxtp_1 DFF_1600_Q_reg( .D(n5261), .CLK(CLK), .Q(n7716) );
	dfxtp_1 DFF_1061_Q_reg( .D(n4931), .CLK(CLK), .Q(n7589) );
	dfxtp_1 DFF_1604_Q_reg( .D(n5265), .CLK(CLK), .Q(n7326) );
	dfxtp_1 DFF_1410_Q_reg( .D(n5161), .CLK(CLK), .Q(n7290) );
	dfxtp_1 DFF_1291_Q_reg( .D(n5108), .CLK(CLK), .Q(n7696) );
	dfxtp_1 DFF_1287_Q_reg( .D(n5104), .CLK(CLK), .Q(n7699) );
	dfxtp_1 DFF_941_Q_reg( .D(n4878), .CLK(CLK), .Q(n7697) );
	dfxtp_1 DFF_237_Q_reg( .D(n4415), .CLK(CLK), .Q(n7702) );
	dfxtp_1 DFF_241_Q_reg( .D(n4419), .CLK(CLK), .Q(n7304) );
	dfxtp_1 DFF_591_Q_reg( .D(n4649), .CLK(CLK), .Q(n7698) );
	dfxtp_1 DFF_62_Q_reg( .D(n147), .CLK(CLK), .Q(n7593) );
	dfxtp_1 DFF_45_Q_reg( .D(n5282), .CLK(CLK), .Q(n7243) );
	dfxtp_1 DFF_76_Q_reg( .D(n164), .CLK(CLK), .Q(n7233) );
	dfxtp_1 DFF_66_Q_reg( .D(n149), .CLK(CLK), .Q(n7223) );
	dfxtp_1 DFF_48_Q_reg( .D(n120), .CLK(CLK), .Q(n7222) );
	dfxtp_1 DFF_711_Q_reg( .D(n4702), .CLK(CLK), .Q(n7590) );
	dfxtp_1 DFF_361_Q_reg( .D(n4473), .CLK(CLK), .Q(n7591) );
	dfxtp_1 DFF_1606_Q_reg( .D(n5267), .CLK(CLK), .Q(n7254) );
	dfxtp_1 DFF_752_Q_reg( .D(n4211), .CLK(CLK), .Q(g1186) );
	dfxtp_1 DFF_1102_Q_reg( .D(n4208), .CLK(CLK), .Q(g1880) );
	dfxtp_1 DFF_11_Q_reg( .D(n4272), .CLK(CLK), .Q(n7303) );
	dfxtp_1 DFF_1300_Q_reg( .D(n3960), .CLK(CLK), .Q(g7264) );
	dfxtp_1 DFF_38_Q_reg( .D(n5275), .CLK(CLK), .Q(n7268) );
	dfxtp_1 DFF_72_Q_reg( .D(n157), .CLK(CLK), .Q(n7244) );
	dfxtp_1 DFF_86_Q_reg( .D(n5286), .CLK(CLK), .Q(n7273) );
	dfxtp_1 DFF_41_Q_reg( .D(n5278), .CLK(CLK), .Q(n7274) );
	dfxtp_1 DFF_1512_Q_reg( .D(n5210), .CLK(CLK), .Q(n7299) );
	dfxtp_1 DFF_462_Q_reg( .D(n4523), .CLK(CLK), .Q(n7302) );
	dfxtp_1 DFF_812_Q_reg( .D(n4752), .CLK(CLK), .Q(n7301) );
	dfxtp_1 DFF_1563_Q_reg( .D(n4047), .CLK(CLK), .Q(g3080) );
	dfxtp_1 DFF_9_Q_reg( .D(n4270), .CLK(CLK), .Q(n7320) );
	dfxtp_1 DFF_593_Q_reg( .D(n4651), .CLK(CLK), .Q(n7707) );
	dfxtp_1 DFF_243_Q_reg( .D(n4421), .CLK(CLK), .Q(n7708) );
	dfxtp_1 DFF_943_Q_reg( .D(n4880), .CLK(CLK), .Q(n7706) );
	dfxtp_1 DFF_1293_Q_reg( .D(n5110), .CLK(CLK), .Q(n7705) );
	dfxtp_1 DFF_44_Q_reg( .D(n5281), .CLK(CLK), .Q(n7585) );
	dfxtp_1 DFF_58_Q_reg( .D(n136), .CLK(CLK), .Q(n7592) );
	dfxtp_1 DFF_1298_Q_reg( .D(n5113), .CLK(CLK), .Q(n7720) );
	dfxtp_1 DFF_948_Q_reg( .D(n4883), .CLK(CLK), .Q(n7717) );
	dfxtp_1 DFF_598_Q_reg( .D(n4654), .CLK(CLK), .Q(n7718) );
	dfxtp_1 DFF_248_Q_reg( .D(n4424), .CLK(CLK), .Q(n7719) );
	dfxtp_1 DFF_84_Q_reg( .D(n5284), .CLK(CLK), .Q(n7232) );
	dfxtp_1 DFF_50_Q_reg( .D(n121), .CLK(CLK), .Q(n7240) );
	dfxtp_1 DFF_78_Q_reg( .D(n165), .CLK(CLK), .Q(n7252) );
	dfxtp_1 DFF_60_Q_reg( .D(n137), .CLK(CLK), .Q(n7251) );
	dfxtp_1 DFF_89_Q_reg( .D(n5289), .CLK(CLK), .Q(n7586) );
	dfxtp_1 DFF_39_Q_reg( .D(n5276), .CLK(CLK), .Q(n7234) );
	dfxtp_1 DFF_402_Q_reg( .D(n4210), .CLK(CLK), .Q(g499) );
	dfxtp_1 DFF_1452_Q_reg( .D(n4212), .CLK(CLK), .Q(g2574) );
	dfxtp_1 DFF_708_Q_reg( .D(n153), .CLK(CLK), .Q(n7226) );
	dfxtp_1 DFF_1408_Q_reg( .D(n59), .CLK(CLK), .Q(n7224) );
	dfxtp_1 DFF_1058_Q_reg( .D(n21), .CLK(CLK), .Q(n7225) );
	dfxtp_1 DFF_358_Q_reg( .D(n110), .CLK(CLK), .Q(n7227) );
	dfxtp_1 DFF_250_Q_reg( .D(n3958), .CLK(CLK), .Q(g6447) );
	dfxtp_1 DFF_7_Q_reg( .D(n4268), .CLK(CLK), .Q(n7279) );
	dfxtp_1 DFF_5_Q_reg( .D(n4266), .CLK(CLK), .Q(n7721) );
	dfxtp_1 DFF_1603_Q_reg( .D(n5264), .CLK(CLK), .Q(n7249) );
	dfxtp_1 DFF_950_Q_reg( .D(n3959), .CLK(CLK), .Q(g7014) );
	dfxtp_1 DFF_135_Q_reg( .D(n4337), .CLK(CLK), .Q(n7319) );
	dfxtp_1 DFF_87_Q_reg( .D(n5287), .CLK(CLK), .Q(n7235) );
	dfxtp_1 DFF_88_Q_reg( .D(n5288), .CLK(CLK), .Q(n7250) );
	dfxtp_1 DFF_43_Q_reg( .D(n5280), .CLK(CLK), .Q(n7246) );
	dfxtp_1 DFF_74_Q_reg( .D(n163), .CLK(CLK), .Q(n7282) );
	dfxtp_1 DFF_56_Q_reg( .D(n135), .CLK(CLK), .Q(n7248) );
	dfxtp_1 DFF_83_Q_reg( .D(n5283), .CLK(CLK), .Q(n7267) );
	dfxtp_1 DFF_54_Q_reg( .D(n134), .CLK(CLK), .Q(n7245) );
	dfxtp_1 DFF_42_Q_reg( .D(n5279), .CLK(CLK), .Q(n7271) );
	dfxtp_1 DFF_1162_Q_reg( .D(n4982), .CLK(CLK), .Q(n7300) );
	dfxtp_1 DFF_1160_Q_reg( .D(n4981), .CLK(CLK), .Q(n7690) );
	dfxtp_1 DFF_1164_Q_reg( .D(n4984), .CLK(CLK), .Q(n7296) );
	dfxtp_1 DFF_1510_Q_reg( .D(n5209), .CLK(CLK), .Q(n7689) );
	dfxtp_1 DFF_1514_Q_reg( .D(n5212), .CLK(CLK), .Q(n7295) );
	dfxtp_1 DFF_460_Q_reg( .D(n4522), .CLK(CLK), .Q(n7688) );
	dfxtp_1 DFF_810_Q_reg( .D(n4751), .CLK(CLK), .Q(n7691) );
	dfxtp_1 DFF_952_Q_reg( .D(n4883), .CLK(CLK), .Q(n7265) );
	dfxtp_1 DFF_464_Q_reg( .D(n4525), .CLK(CLK), .Q(n7298) );
	dfxtp_1 DFF_814_Q_reg( .D(n4754), .CLK(CLK), .Q(n7297) );
	dfxtp_1 DFF_455_Q_reg( .D(n5291), .CLK(CLK), .Q(g6911) );
	dfxtp_1 DFF_1155_Q_reg( .D(n5297), .CLK(CLK), .Q(g7357) );
	dfxtp_1 DFF_1505_Q_reg( .D(n5300), .CLK(CLK), .Q(g7487) );
	dfxtp_1 DFF_805_Q_reg( .D(n5294), .CLK(CLK), .Q(g7161) );
	dfxtp_1 DFF_249_Q_reg( .D(n4131), .CLK(CLK), .Q(g5437) );
	dfxtp_1 DFF_1299_Q_reg( .D(n4131), .CLK(CLK), .Q(g5555) );
	dfxtp_1 DFF_456_Q_reg( .D(n5292), .CLK(CLK), .Q(n7239) );
	dfxtp_1 DFF_1156_Q_reg( .D(n5298), .CLK(CLK), .Q(n7237) );
	dfxtp_1 DFF_1506_Q_reg( .D(n5301), .CLK(CLK), .Q(n7236) );
	dfxtp_1 DFF_806_Q_reg( .D(n5295), .CLK(CLK), .Q(n7238) );
	dfxtp_1 DFF_1166_Q_reg( .D(n4986), .CLK(CLK), .Q(n7692) );
	dfxtp_1 DFF_1516_Q_reg( .D(n5214), .CLK(CLK), .Q(n7695) );
	dfxtp_1 DFF_466_Q_reg( .D(n4527), .CLK(CLK), .Q(n7694) );
	dfxtp_1 DFF_816_Q_reg( .D(n4756), .CLK(CLK), .Q(n7693) );
	dfxtp_1 DFF_137_Q_reg( .D(n4339), .CLK(CLK), .Q(n7262) );
	dfxtp_1 DFF_600_Q_reg( .D(n138), .CLK(CLK), .Q(g6712) );
	dfxtp_1 DFF_863_Q_reg( .D(n170), .CLK(CLK), .Q(n7229) );
	dfxtp_1 DFF_163_Q_reg( .D(n91), .CLK(CLK), .Q(n7230) );
	dfxtp_1 DFF_513_Q_reg( .D(n124), .CLK(CLK), .Q(n7231) );
	dfxtp_1 DFF_1302_Q_reg( .D(n5113), .CLK(CLK), .Q(n7264) );
	dfxtp_1 DFF_252_Q_reg( .D(n4424), .CLK(CLK), .Q(n7266) );
	dfxtp_1 DFF_602_Q_reg( .D(n4654), .CLK(CLK), .Q(n7263) );
	dfxtp_1 DFF_951_Q_reg( .D(n172), .CLK(CLK), .Q(n7782) );
	dfxtp_1 DFF_949_Q_reg( .D(n4131), .CLK(CLK), .Q(g5511) );
	dfxtp_1 DFF_160_Q_reg( .D(n4341), .CLK(CLK), .Q(n7256) );
	dfxtp_1 DFF_1301_Q_reg( .D(n48), .CLK(CLK), .Q(n7780) );
	dfxtp_1 DFF_251_Q_reg( .D(n100), .CLK(CLK), .Q(n7784) );
	dfxtp_1 DFF_1213_Q_reg( .D(n37), .CLK(CLK), .Q(n7228) );
	dfxtp_1 DFF_599_Q_reg( .D(n4131), .CLK(CLK), .Q(g5472) );
	dfxtp_1 DFF_601_Q_reg( .D(n3961), .CLK(CLK), .Q(n7775) );
	dfxtp_1 DFF_707_Q_reg( .D(n152), .CLK(CLK), .Q(g6944) );
	dfxtp_1 DFF_1407_Q_reg( .D(n58), .CLK(CLK), .Q(g7390) );
	dfxtp_1 DFF_1057_Q_reg( .D(n20), .CLK(CLK), .Q(g7194) );
	dfxtp_1 DFF_706_Q_reg( .D(n4231), .CLK(CLK), .Q(g6750) );
	dfxtp_1 DFF_1406_Q_reg( .D(n4231), .CLK(CLK), .Q(g7302) );
	dfxtp_1 DFF_1056_Q_reg( .D(n4231), .CLK(CLK), .Q(g7052) );
	dfxtp_1 DFF_357_Q_reg( .D(n109), .CLK(CLK), .Q(g6642) );
	dfxtp_1 DFF_356_Q_reg( .D(n4231), .CLK(CLK), .Q(g6485) );
	dfxtp_1 DFF_454_Q_reg( .D(n4231), .CLK(CLK), .Q(g6677) );
	dfxtp_1 DFF_1154_Q_reg( .D(n4231), .CLK(CLK), .Q(g7229) );
	dfxtp_1 DFF_1504_Q_reg( .D(n4231), .CLK(CLK), .Q(g7425) );
	dfxtp_1 DFF_804_Q_reg( .D(n4231), .CLK(CLK), .Q(g6979) );
	dfxtp_1 DFF_512_Q_reg( .D(n123), .CLK(CLK), .Q(g6518) );
	dfxtp_1 DFF_1212_Q_reg( .D(n36), .CLK(CLK), .Q(g7084) );
	dfxtp_1 DFF_862_Q_reg( .D(n169), .CLK(CLK), .Q(g6782) );
	dfxtp_1 DFF_162_Q_reg( .D(n90), .CLK(CLK), .Q(g6313) );
	dfxtp_1 DFF_1211_Q_reg( .D(n4131), .CLK(CLK), .Q(g6837) );
	dfxtp_1 DFF_511_Q_reg( .D(n4131), .CLK(CLK), .Q(g6368) );
	dfxtp_1 DFF_861_Q_reg( .D(n4131), .CLK(CLK), .Q(g6573) );
	dfxtp_1 DFF_161_Q_reg( .D(n4131), .CLK(CLK), .Q(g6231) );
	inv_2 U5578( .A(RST), .Y(n5740) );
	inv_2 U5579( .A(RST), .Y(n5742) );
	inv_2 U5580( .A(RST), .Y(n5746) );
	inv_2 U5581( .A(RST), .Y(n5750) );
	inv_2 U5582( .A(RST), .Y(n5743) );
	inv_2 U5583( .A(RST), .Y(n5744) );
	inv_2 U5584( .A(RST), .Y(n5749) );
	inv_2 U5585( .A(RST), .Y(n5747) );
	inv_2 U5586( .A(RST), .Y(n5748) );
	inv_2 U5587( .A(RST), .Y(n5753) );
	inv_2 U5588( .A(RST), .Y(n5754) );
	inv_2 U5589( .A(RST), .Y(n5745) );
	inv_2 U5590( .A(RST), .Y(n5752) );
	inv_2 U5591( .A(RST), .Y(n5751) );
	inv_2 U5592( .A(RST), .Y(n5741) );
	inv_2 U5593( .A(RST), .Y(n5755) );
	inv_2 U5594( .A(RST), .Y(n5757) );
	inv_2 U5595( .A(RST), .Y(n5756) );
	inv_2 U5596( .A(RST), .Y(n5758) );
	inv_2 U5597( .A(RST), .Y(n5762) );
	inv_2 U5598( .A(RST), .Y(n5760) );
	inv_2 U5599( .A(RST), .Y(n5759) );
	inv_2 U5600( .A(RST), .Y(n5761) );
	inv_2 U5601( .A(RST), .Y(n5763) );
	inv_2 U5602( .A(RST), .Y(n5764) );
	inv_2 U5603( .A(RST), .Y(n5765) );
	inv_1 U5604( .A(n5766), .Y(n89) );
	a22oi_1 U5605( .A1(g2997), .A2(n5767), .B1(g3061), .B2(n5768), .Y(n5766) );
	inv_1 U5606( .A(n5769), .Y(n88) );
	a22oi_1 U5607( .A1(g3078), .A2(n5767), .B1(g3060), .B2(n5768), .Y(n5769) );
	inv_1 U5608( .A(n5770), .Y(n87) );
	a22oi_1 U5609( .A1(g3077), .A2(n5767), .B1(g3059), .B2(n5768), .Y(n5770) );
	inv_1 U5610( .A(n5771), .Y(n86) );
	a22oi_1 U5611( .A1(g3076), .A2(n5767), .B1(g3058), .B2(n5768), .Y(n5771) );
	inv_1 U5612( .A(n5772), .Y(n85) );
	a22oi_1 U5613( .A1(g3075), .A2(n5767), .B1(g3057), .B2(n5768), .Y(n5772) );
	inv_1 U5614( .A(n5773), .Y(n84) );
	a22oi_1 U5615( .A1(g3074), .A2(n5767), .B1(g3056), .B2(n5768), .Y(n5773) );
	inv_1 U5616( .A(n5774), .Y(n83) );
	a22oi_1 U5617( .A1(g3073), .A2(n5767), .B1(g3055), .B2(n5768), .Y(n5774) );
	inv_1 U5618( .A(n5775), .Y(n82) );
	a22oi_1 U5619( .A1(g3072), .A2(n5767), .B1(g3053), .B2(n5768), .Y(n5775) );
	inv_1 U5620( .A(n5776), .Y(n81) );
	a22oi_1 U5621( .A1(g3071), .A2(n5767), .B1(g3052), .B2(n5768), .Y(n5776) );
	inv_1 U5622( .A(n5777), .Y(n80) );
	a22oi_1 U5623( .A1(g3070), .A2(n5767), .B1(g3051), .B2(n5768), .Y(n5777) );
	inv_1 U5624( .A(n5778), .Y(n79) );
	a22oi_1 U5625( .A1(g3069), .A2(n5767), .B1(g3050), .B2(n5768), .Y(n5778) );
	inv_1 U5626( .A(n5779), .Y(n78) );
	a22oi_1 U5627( .A1(g3068), .A2(n5767), .B1(g3049), .B2(n5768), .Y(n5779) );
	inv_1 U5628( .A(n5780), .Y(n77) );
	a22oi_1 U5629( .A1(g3067), .A2(n5767), .B1(g3048), .B2(n5768), .Y(n5780) );
	inv_1 U5630( .A(n5781), .Y(n76) );
	a22oi_1 U5631( .A1(g3066), .A2(n5767), .B1(g3047), .B2(n5768), .Y(n5781) );
	inv_1 U5632( .A(n5782), .Y(n75) );
	a22oi_1 U5633( .A1(g3065), .A2(n5767), .B1(g3046), .B2(n5768), .Y(n5782) );
	inv_1 U5634( .A(n5783), .Y(n74) );
	a22oi_1 U5635( .A1(g3064), .A2(n5767), .B1(g3045), .B2(n5768), .Y(n5783) );
	inv_1 U5636( .A(n5784), .Y(n73) );
	a22oi_1 U5637( .A1(g3063), .A2(n5767), .B1(g3044), .B2(n5768), .Y(n5784) );
	inv_1 U5638( .A(n5785), .Y(n72) );
	a22oi_1 U5639( .A1(g3062), .A2(n5767), .B1(g3043), .B2(n5768), .Y(n5785) );
	nor2_1 U5640( .A(RST), .B(n7255), .Y(n5768) );
	and2_0 U5641( .A(n7255), .B(n5761), .X(n5767) );
	inv_1 U5642( .A(n5786), .Y(n69) );
	inv_1 U5643( .A(n5787), .Y(n67) );
	inv_1 U5644( .A(n5788), .Y(n66) );
	inv_1 U5645( .A(n5789), .Y(n65) );
	inv_1 U5646( .A(n5790), .Y(n64) );
	inv_1 U5647( .A(n5791), .Y(n63) );
	inv_1 U5648( .A(n5792), .Y(n62) );
	inv_1 U5649( .A(n5793), .Y(n61) );
	inv_1 U5650( .A(n5794), .Y(n60) );
	inv_1 U5651( .A(n5795), .Y(n57) );
	inv_1 U5652( .A(n5796), .Y(n56) );
	inv_1 U5653( .A(n5797), .Y(n55) );
	inv_1 U5654( .A(n5798), .Y(n54) );
	and2_0 U5655( .A(n5758), .B(g16496), .X(n5303) );
	inv_1 U5656( .A(n5799), .Y(n5302) );
	o211ai_1 U5657( .A1(n9951), .A2(n5800), .B1(n5801), .C1(n5802), .Y(n5799) );
	inv_1 U5658( .A(n5803), .Y(n5300) );
	inv_1 U5659( .A(n5804), .Y(n53) );
	inv_1 U5660( .A(n5805), .Y(n5299) );
	o211ai_1 U5661( .A1(n9952), .A2(n5806), .B1(n5807), .C1(n5808), .Y(n5805) );
	inv_1 U5662( .A(n5809), .Y(n5297) );
	inv_1 U5663( .A(n5810), .Y(n5296) );
	o211ai_1 U5664( .A1(n9953), .A2(n5811), .B1(n5812), .C1(n5813), .Y(n5810) );
	inv_1 U5665( .A(n5814), .Y(n5294) );
	inv_1 U5666( .A(n5815), .Y(n5293) );
	o211ai_1 U5667( .A1(n9954), .A2(n5816), .B1(n5817), .C1(n5818), .Y(n5815) );
	inv_1 U5668( .A(n5819), .Y(n5291) );
	o22ai_1 U5669( .A1(n5820), .A2(n5821), .B1(n5822), .B2(n5823), .Y(n5290) );
	o22ai_1 U5670( .A1(n5820), .A2(n5824), .B1(n5822), .B2(n5825), .Y(n5289) );
	o22ai_1 U5671( .A1(n5820), .A2(n5826), .B1(n5822), .B2(n5827), .Y(n5288) );
	o22ai_1 U5672( .A1(n5820), .A2(n5828), .B1(n5822), .B2(n5829), .Y(n5287) );
	o22ai_1 U5673( .A1(n5820), .A2(n5830), .B1(n5822), .B2(n5831), .Y(n5286) );
	o22ai_1 U5674( .A1(n5820), .A2(n5832), .B1(n5822), .B2(n5833), .Y(n5285) );
	o22ai_1 U5675( .A1(n5820), .A2(n5834), .B1(n5822), .B2(n5835), .Y(n5284) );
	o22ai_1 U5676( .A1(n5820), .A2(n5836), .B1(n5822), .B2(n5837), .Y(n5283) );
	o22ai_1 U5677( .A1(n5820), .A2(n5838), .B1(n5822), .B2(n5839), .Y(n5282) );
	o22ai_1 U5678( .A1(n5820), .A2(n5840), .B1(n5822), .B2(n5841), .Y(n5281) );
	o22ai_1 U5679( .A1(n5820), .A2(n5842), .B1(n5822), .B2(n5843), .Y(n5280) );
	o22ai_1 U5680( .A1(n5820), .A2(n5844), .B1(n5822), .B2(n5845), .Y(n5279) );
	o22ai_1 U5681( .A1(n5820), .A2(n5846), .B1(n5822), .B2(n5847), .Y(n5278) );
	o22ai_1 U5682( .A1(n5820), .A2(n5848), .B1(n5822), .B2(n5849), .Y(n5277) );
	o22ai_1 U5683( .A1(n5820), .A2(n5850), .B1(n5822), .B2(n5851), .Y(n5276) );
	o22ai_1 U5684( .A1(n5820), .A2(n5852), .B1(n5822), .B2(n5853), .Y(n5275) );
	nor2_1 U5685( .A(RST), .B(n5854), .Y(n5274) );
	xor2_1 U5686( .A(n5855), .B(g2990), .X(n5854) );
	nor2_1 U5687( .A(RST), .B(n5856), .Y(n5273) );
	xor2_1 U5688( .A(n5857), .B(g3083), .X(n5856) );
	nor2_1 U5689( .A(RST), .B(n5858), .Y(n5272) );
	nor2_1 U5690( .A(n5859), .B(n5860), .Y(n5271) );
	xnor2_1 U5691( .A(n5861), .B(n10034), .Y(n5859) );
	nor3_1 U5692( .A(n5860), .B(n5861), .C(n5862), .Y(n5270) );
	a21oi_1 U5693( .A1(n9955), .A2(n5863), .B1(n7704), .Y(n5862) );
	nor3_1 U5694( .A(n5864), .B(n5865), .C(n5370), .Y(n5861) );
	nor2_1 U5695( .A(n5866), .B(n5860), .Y(n5269) );
	nand3_1 U5696( .A(n5750), .B(n5867), .C(n5868), .Y(n5860) );
	xnor2_1 U5697( .A(n9955), .B(n5863), .Y(n5866) );
	o211ai_1 U5698( .A1(RST), .A2(n5869), .B1(n5870), .C1(n5871), .Y(n5268) );
	nand3_1 U5699( .A(n5872), .B(n5865), .C(n4231), .Y(n5870) );
	a21oi_1 U5700( .A1(n9956), .A2(n5865), .B1(n5873), .Y(n5869) );
	inv_1 U5701( .A(n5868), .Y(n5873) );
	nand4_1 U5702( .A(n10034), .B(n5863), .C(n5864), .D(n5370), .Y(n5868) );
	inv_1 U5703( .A(n7704), .Y(n5864) );
	inv_1 U5704( .A(n5865), .Y(n5863) );
	nand3_1 U5705( .A(g3080), .B(n5872), .C(n9956), .Y(n5865) );
	inv_1 U5706( .A(n5874), .Y(n5872) );
	nor2_1 U5707( .A(n5875), .B(n5876), .Y(n5267) );
	xnor2_1 U5708( .A(n7254), .B(n5877), .Y(n5875) );
	and2_0 U5709( .A(n5878), .B(n10083), .X(n5877) );
	nor2_1 U5710( .A(n5879), .B(n5876), .Y(n5266) );
	xnor2_1 U5711( .A(n5878), .B(n10083), .Y(n5879) );
	nor3_1 U5712( .A(n5876), .B(n5878), .C(n5880), .Y(n5265) );
	a21oi_1 U5713( .A1(n5881), .A2(n7249), .B1(n7326), .Y(n5880) );
	and3_1 U5714( .A(n7326), .B(n7249), .C(n5881), .X(n5878) );
	nor2_1 U5715( .A(n5882), .B(n5876), .Y(n5264) );
	xnor2_1 U5716( .A(n5881), .B(n7249), .Y(n5882) );
	nor3_1 U5717( .A(n5876), .B(n5881), .C(n5883), .Y(n5263) );
	a21oi_1 U5718( .A1(n5884), .A2(n7283), .B1(n10082), .Y(n5883) );
	and3_1 U5719( .A(n5884), .B(n7283), .C(n10082), .X(n5881) );
	o21ai_0 U5720( .A1(n5885), .A2(n5876), .B1(n5871), .Y(n5262) );
	xnor2_1 U5721( .A(n5884), .B(n7283), .Y(n5885) );
	and2_0 U5722( .A(n7716), .B(g3080), .X(n5884) );
	o22ai_1 U5723( .A1(n5874), .A2(n5886), .B1(n5887), .B2(n5876), .Y(n5261) );
	o211ai_1 U5724( .A1(n5874), .A2(n5888), .B1(n5741), .C1(n5867), .Y(n5876) );
	xnor2_1 U5725( .A(n7716), .B(g3080), .Y(n5887) );
	nor3_1 U5726( .A(n15502), .B(g3234), .C(RST), .Y(n5260) );
	inv_1 U5727( .A(n5886), .Y(n5259) );
	nand2_1 U5728( .A(n4231), .B(n5867), .Y(n5886) );
	a21oi_1 U5729( .A1(n5889), .A2(n5890), .B1(n5891), .Y(n5258) );
	a21oi_1 U5730( .A1(n5334), .A2(n5892), .B1(n5893), .Y(n5257) );
	a21oi_1 U5731( .A1(n5543), .A2(n5894), .B1(n5895), .Y(n5256) );
	o22ai_1 U5732( .A1(n5896), .A2(n5897), .B1(n5898), .B2(n5899), .Y(n5255) );
	inv_1 U5733( .A(n7475), .Y(n5897) );
	o22ai_1 U5734( .A1(n5900), .A2(n5901), .B1(n5898), .B2(n5902), .Y(n5254) );
	inv_1 U5735( .A(n7498), .Y(n5901) );
	o22ai_1 U5736( .A1(n5903), .A2(n5904), .B1(n5898), .B2(n5905), .Y(n5253) );
	nand4_1 U5737( .A(n5906), .B(n5907), .C(n5908), .D(n5909), .Y(n5898) );
	a222oi_1 U5738( .A1(g7487), .A2(n5910), .B1(n7236), .B2(n5911), .C1(g7425), .C2(n5390), .Y(n5909) );
	nand2_1 U5739( .A(n9871), .B(n10037), .Y(n5911) );
	nand4_1 U5740( .A(n5912), .B(n5913), .C(n5914), .D(n5915), .Y(n5908) );
	nor3_1 U5741( .A(n5916), .B(n5917), .C(n5918), .Y(n5915) );
	xor2_1 U5742( .A(n5919), .B(n10040), .X(n5918) );
	xor2_1 U5743( .A(n5920), .B(n7689), .X(n5917) );
	nand3_1 U5744( .A(n5921), .B(n5922), .C(n5923), .Y(n5916) );
	xor2_1 U5745( .A(n9951), .B(n5924), .X(n5923) );
	xnor2_1 U5746( .A(n10041), .B(n5925), .Y(n5922) );
	xnor2_1 U5747( .A(n10042), .B(n5926), .Y(n5921) );
	nor3_1 U5748( .A(n5927), .B(n5928), .C(n5929), .Y(n5914) );
	xor2_1 U5749( .A(n5930), .B(n9957), .X(n5929) );
	xor2_1 U5750( .A(n5931), .B(n7295), .X(n5928) );
	xnor2_1 U5751( .A(n5932), .B(n5933), .Y(n5927) );
	xnor2_1 U5752( .A(n10038), .B(n5934), .Y(n5913) );
	xnor2_1 U5753( .A(n7695), .B(n5935), .Y(n5912) );
	o22ai_1 U5754( .A1(n5891), .A2(n5570), .B1(n5936), .B2(n5937), .Y(n5252) );
	o22ai_1 U5755( .A1(n5893), .A2(n5938), .B1(n5936), .B2(n5939), .Y(n5251) );
	o22ai_1 U5756( .A1(n5895), .A2(n5448), .B1(n5936), .B2(n5803), .Y(n5250) );
	or2_0 U5757( .A(n5940), .B(n5357), .X(n5936) );
	o22ai_1 U5758( .A1(n5891), .A2(n5605), .B1(n5937), .B2(n5941), .Y(n5249) );
	o21ai_0 U5759( .A1(n5357), .A2(n5942), .B1(n5765), .Y(n5891) );
	o22ai_1 U5760( .A1(n5893), .A2(n5910), .B1(n5939), .B2(n5941), .Y(n5248) );
	inv_1 U5761( .A(n5301), .Y(n5939) );
	nor2_1 U5762( .A(n5943), .B(RST), .Y(n5301) );
	inv_1 U5763( .A(n7447), .Y(n5910) );
	o22ai_1 U5764( .A1(n5895), .A2(n5390), .B1(n5803), .B2(n5941), .Y(n5247) );
	or2_0 U5765( .A(n5944), .B(n5357), .X(n5941) );
	nand2_1 U5766( .A(g7425), .B(n5750), .Y(n5803) );
	o21ai_0 U5767( .A1(n5357), .A2(n5945), .B1(n5757), .Y(n5895) );
	o22ai_1 U5768( .A1(n5896), .A2(n5946), .B1(n10041), .B2(n5899), .Y(n5246) );
	inv_1 U5769( .A(n7477), .Y(n5946) );
	o22ai_1 U5770( .A1(n5900), .A2(n5947), .B1(n10041), .B2(n5902), .Y(n5245) );
	inv_1 U5771( .A(n7476), .Y(n5947) );
	o22ai_1 U5772( .A1(n5903), .A2(n5443), .B1(n10041), .B2(n5905), .Y(n5244) );
	o22ai_1 U5773( .A1(n5896), .A2(n5948), .B1(n10042), .B2(n5899), .Y(n5243) );
	inv_1 U5774( .A(n7479), .Y(n5948) );
	o22ai_1 U5775( .A1(n5900), .A2(n5949), .B1(n10042), .B2(n5902), .Y(n5242) );
	inv_1 U5776( .A(n7478), .Y(n5949) );
	o22ai_1 U5777( .A1(n5903), .A2(n5446), .B1(n10042), .B2(n5905), .Y(n5241) );
	o22ai_1 U5778( .A1(n5896), .A2(n5950), .B1(n7695), .B2(n5899), .Y(n5240) );
	inv_1 U5779( .A(n7488), .Y(n5950) );
	o22ai_1 U5780( .A1(n5900), .A2(n5951), .B1(n7695), .B2(n5902), .Y(n5239) );
	inv_1 U5781( .A(n7487), .Y(n5951) );
	o22ai_1 U5782( .A1(n5903), .A2(n5452), .B1(n7695), .B2(n5905), .Y(n5238) );
	o22ai_1 U5783( .A1(n5896), .A2(n5952), .B1(n10038), .B2(n5899), .Y(n5237) );
	inv_1 U5784( .A(n7490), .Y(n5952) );
	o22ai_1 U5785( .A1(n5900), .A2(n5953), .B1(n10038), .B2(n5902), .Y(n5236) );
	inv_1 U5786( .A(n7489), .Y(n5953) );
	o22ai_1 U5787( .A1(n5903), .A2(n5450), .B1(n10038), .B2(n5905), .Y(n5235) );
	o22ai_1 U5788( .A1(n5896), .A2(n5954), .B1(n7295), .B2(n5899), .Y(n5234) );
	inv_1 U5789( .A(n7492), .Y(n5954) );
	o22ai_1 U5790( .A1(n5900), .A2(n5955), .B1(n7295), .B2(n5902), .Y(n5233) );
	inv_1 U5791( .A(n7491), .Y(n5955) );
	o22ai_1 U5792( .A1(n5903), .A2(n5449), .B1(n7295), .B2(n5905), .Y(n5232) );
	o22ai_1 U5793( .A1(n5896), .A2(n5956), .B1(n10040), .B2(n5899), .Y(n5231) );
	inv_1 U5794( .A(n7494), .Y(n5956) );
	o22ai_1 U5795( .A1(n5900), .A2(n5957), .B1(n10040), .B2(n5902), .Y(n5230) );
	inv_1 U5796( .A(n7493), .Y(n5957) );
	o22ai_1 U5797( .A1(n5903), .A2(n5447), .B1(n10040), .B2(n5905), .Y(n5229) );
	o22ai_1 U5798( .A1(n5896), .A2(n5958), .B1(n7299), .B2(n5899), .Y(n5228) );
	inv_1 U5799( .A(n7485), .Y(n5958) );
	o22ai_1 U5800( .A1(n5900), .A2(n5959), .B1(n7299), .B2(n5902), .Y(n5227) );
	inv_1 U5801( .A(n7484), .Y(n5959) );
	o22ai_1 U5802( .A1(n5903), .A2(n5445), .B1(n7299), .B2(n5905), .Y(n5226) );
	o22ai_1 U5803( .A1(n5896), .A2(n5960), .B1(n9951), .B2(n5899), .Y(n5225) );
	o22ai_1 U5804( .A1(n5900), .A2(n5961), .B1(n9951), .B2(n5902), .Y(n5224) );
	o22ai_1 U5805( .A1(n5903), .A2(n5606), .B1(n9951), .B2(n5905), .Y(n5223) );
	o22ai_1 U5806( .A1(n5896), .A2(n5962), .B1(n7689), .B2(n5899), .Y(n5222) );
	inv_1 U5807( .A(n7483), .Y(n5962) );
	o22ai_1 U5808( .A1(n5900), .A2(n5963), .B1(n7689), .B2(n5902), .Y(n5221) );
	inv_1 U5809( .A(n7482), .Y(n5963) );
	o22ai_1 U5810( .A1(n5903), .A2(n5444), .B1(n7689), .B2(n5905), .Y(n5220) );
	o22ai_1 U5811( .A1(n5896), .A2(n5964), .B1(n9957), .B2(n5899), .Y(n5219) );
	or2_0 U5812( .A(n5890), .B(RST), .X(n5899) );
	inv_1 U5813( .A(n7496), .Y(n5964) );
	nand2_1 U5814( .A(n5755), .B(n5890), .Y(n5896) );
	nand3_1 U5815( .A(n9959), .B(n5965), .C(n9872), .Y(n5890) );
	o22ai_1 U5816( .A1(n5900), .A2(n5966), .B1(n9957), .B2(n5902), .Y(n5218) );
	or2_0 U5817( .A(n5892), .B(RST), .X(n5902) );
	inv_1 U5818( .A(n7495), .Y(n5966) );
	nand2_1 U5819( .A(n5755), .B(n5892), .Y(n5900) );
	nand2_1 U5820( .A(n5967), .B(g7487), .Y(n5892) );
	o22ai_1 U5821( .A1(n5903), .A2(n5451), .B1(n9957), .B2(n5905), .Y(n5217) );
	or2_0 U5822( .A(n5894), .B(RST), .X(n5905) );
	nand2_1 U5823( .A(n5757), .B(n5894), .Y(n5903) );
	nand2_1 U5824( .A(n5967), .B(g7425), .Y(n5894) );
	and3_1 U5825( .A(n9959), .B(n5968), .C(n9872), .X(n5967) );
	nor2_1 U5826( .A(n5969), .B(n5893), .Y(n5216) );
	xnor2_1 U5827( .A(n5970), .B(n10041), .Y(n5969) );
	a211oi_1 U5828( .A1(n5365), .A2(n5971), .B1(n5893), .C1(n5970), .Y(n5215) );
	nor2_1 U5829( .A(n5971), .B(n5365), .Y(n5970) );
	nor3_1 U5830( .A(n5893), .B(n5972), .C(n5973), .Y(n5214) );
	a21oi_1 U5831( .A1(n5974), .A2(n10038), .B1(n7695), .Y(n5973) );
	inv_1 U5832( .A(n5971), .Y(n5972) );
	nand3_1 U5833( .A(n7695), .B(n10038), .C(n5974), .Y(n5971) );
	nor2_1 U5834( .A(n5975), .B(n5893), .Y(n5213) );
	xnor2_1 U5835( .A(n5974), .B(n10038), .Y(n5975) );
	nor3_1 U5836( .A(n5893), .B(n5974), .C(n5976), .Y(n5212) );
	a21oi_1 U5837( .A1(n5977), .A2(n10040), .B1(n7295), .Y(n5976) );
	and3_1 U5838( .A(n7295), .B(n10040), .C(n5977), .X(n5974) );
	nor2_1 U5839( .A(n5978), .B(n5893), .Y(n5211) );
	xnor2_1 U5840( .A(n10040), .B(n5977), .Y(n5978) );
	a211oi_1 U5841( .A1(n5933), .A2(n5802), .B1(n5893), .C1(n5977), .Y(n5210) );
	nor2_1 U5842( .A(n5802), .B(n5933), .Y(n5977) );
	nand2_1 U5843( .A(n9951), .B(n5800), .Y(n5802) );
	inv_1 U5844( .A(n7299), .Y(n5933) );
	nor3_1 U5845( .A(n5893), .B(n5800), .C(n5979), .Y(n5209) );
	a21oi_1 U5846( .A1(n9957), .A2(n5965), .B1(n7689), .Y(n5979) );
	and3_1 U5847( .A(n7689), .B(n5965), .C(n9957), .X(n5800) );
	nor2_1 U5848( .A(n5980), .B(n5893), .Y(n5208) );
	inv_1 U5849( .A(n5801), .Y(n5893) );
	a21oi_1 U5850( .A1(g7487), .A2(n9958), .B1(RST), .Y(n5801) );
	xnor2_1 U5851( .A(n5965), .B(n9957), .Y(n5980) );
	nor2_1 U5852( .A(n5942), .B(n7275), .Y(n5965) );
	o32ai_1 U5853( .A1(n5968), .A2(n7236), .A3(RST), .B1(n5937), .B2(n5981), .Y(n5207) );
	inv_1 U5854( .A(n7275), .Y(n5968) );
	o32ai_1 U5855( .A1(n5357), .A2(n7236), .A3(RST), .B1(n5937), .B2(n5982), .Y(n5206) );
	nand2_1 U5856( .A(n7236), .B(n5749), .Y(n5937) );
	o22ai_1 U5857( .A1(n5786), .A2(n5983), .B1(n5984), .B2(n5985), .Y(n5205) );
	inv_1 U5858( .A(n7632), .Y(n5985) );
	nand2_1 U5859( .A(n5755), .B(DFF_1503_D), .Y(n5786) );
	o22ai_1 U5860( .A1(n5566), .A2(n5986), .B1(n5987), .B2(n5988), .Y(n5204) );
	o22ai_1 U5861( .A1(n5719), .A2(n5989), .B1(n5988), .B2(n5990), .Y(n5203) );
	o22ai_1 U5862( .A1(n5991), .A2(n5992), .B1(n5988), .B2(n5993), .Y(n5202) );
	or3_1 U5863( .A(n5982), .B(n5944), .C(n5994), .X(n5988) );
	inv_1 U5864( .A(n7636), .Y(n5991) );
	o22ai_1 U5865( .A1(n5561), .A2(n5986), .B1(n5995), .B2(n5987), .Y(n5201) );
	o22ai_1 U5866( .A1(n5351), .A2(n5989), .B1(n5995), .B2(n5990), .Y(n5200) );
	inv_1 U5867( .A(n5996), .Y(n52) );
	o22ai_1 U5868( .A1(n5995), .A2(n5993), .B1(n5997), .B2(n5992), .Y(n5199) );
	inv_1 U5869( .A(n7659), .Y(n5997) );
	mux2i_1 U5870( .A0(n5998), .A1(n5940), .S(n5999), .Y(n5995) );
	nor2_1 U5871( .A(n6000), .B(n6001), .Y(n5998) );
	mux2i_1 U5872( .A0(n6002), .A1(n6003), .S(n6004), .Y(n6000) );
	inv_1 U5873( .A(n6005), .Y(n6003) );
	o22ai_1 U5874( .A1(n5560), .A2(n5986), .B1(n6006), .B2(n5987), .Y(n5198) );
	o22ai_1 U5875( .A1(n5350), .A2(n5989), .B1(n6006), .B2(n5990), .Y(n5197) );
	o22ai_1 U5876( .A1(n6006), .A2(n5993), .B1(n6007), .B2(n5992), .Y(n5196) );
	inv_1 U5877( .A(n7658), .Y(n6007) );
	mux2i_1 U5878( .A0(n6008), .A1(n5944), .S(n5999), .Y(n6006) );
	nor2_1 U5879( .A(n6009), .B(n6002), .Y(n6008) );
	nand2_1 U5880( .A(n6010), .B(n6011), .Y(n6002) );
	mux2i_1 U5881( .A0(n6012), .A1(n6013), .S(n6014), .Y(n6011) );
	nor2_1 U5882( .A(n6015), .B(n6016), .Y(n6013) );
	nor2_1 U5883( .A(n6017), .B(n6018), .Y(n6012) );
	mux2i_1 U5884( .A0(n6019), .A1(n6020), .S(n6021), .Y(n6010) );
	o22ai_1 U5885( .A1(n6022), .A2(n6023), .B1(n6024), .B2(n6014), .Y(n6020) );
	a211oi_1 U5886( .A1(n6025), .A2(n6026), .B1(n6027), .C1(n6028), .Y(n6024) );
	nor3_1 U5887( .A(n6029), .B(n6030), .C(n6031), .Y(n6028) );
	o32ai_1 U5888( .A1(n6017), .A2(n6032), .A3(n6033), .B1(n6034), .B2(n6035), .Y(n6019) );
	a21oi_1 U5889( .A1(n6025), .A2(n6033), .B1(n6036), .Y(n6035) );
	mux2i_1 U5890( .A0(n6030), .A1(n6037), .S(n6017), .Y(n6036) );
	or2_0 U5891( .A(n6023), .B(n6031), .X(n6037) );
	inv_1 U5892( .A(n6014), .Y(n6034) );
	mux2i_1 U5893( .A0(n6001), .A1(n6038), .S(n6005), .Y(n6009) );
	inv_1 U5894( .A(n6004), .Y(n6038) );
	nand2_1 U5895( .A(n6039), .B(n6040), .Y(n6001) );
	nand3_1 U5896( .A(n6031), .B(n6041), .C(n6042), .Y(n6040) );
	inv_1 U5897( .A(n6022), .Y(n6031) );
	mux2i_1 U5898( .A0(n6043), .A1(n6044), .S(n6014), .Y(n6039) );
	o221ai_1 U5899( .A1(n6045), .A2(n15037), .B1(n5353), .B2(n15036), .C1(n6046), .Y(n6014) );
	nand2_1 U5900( .A(g2424), .B(g5747), .Y(n6046) );
	o221ai_1 U5901( .A1(n6047), .A2(n6018), .B1(n6029), .B2(n6048), .C1(n6049), .Y(n6044) );
	mux2i_1 U5902( .A0(n6050), .A1(n6051), .S(n6021), .Y(n6049) );
	nor2_1 U5903( .A(n6052), .B(n6017), .Y(n6051) );
	a21oi_1 U5904( .A1(n6015), .A2(n6047), .B1(n6041), .Y(n6052) );
	nor2_1 U5905( .A(n6022), .B(n6053), .Y(n6050) );
	a211oi_1 U5906( .A1(n6054), .A2(n6022), .B1(n6027), .C1(n6055), .Y(n6048) );
	nor3_1 U5907( .A(n6021), .B(n6030), .C(n6033), .Y(n6055) );
	o221ai_1 U5908( .A1(n6015), .A2(n6056), .B1(n6023), .B2(n6057), .C1(n6058), .Y(n6043) );
	mux2i_1 U5909( .A0(n6059), .A1(n6060), .S(n6021), .Y(n6058) );
	nor3_1 U5910( .A(n6017), .B(n6027), .C(n6054), .Y(n6060) );
	nor2_1 U5911( .A(n6047), .B(n6032), .Y(n6027) );
	nor2_1 U5912( .A(n6061), .B(n6016), .Y(n6059) );
	inv_1 U5913( .A(n6026), .Y(n6016) );
	nor2_1 U5914( .A(n6033), .B(n6029), .Y(n6026) );
	inv_1 U5915( .A(n6017), .Y(n6029) );
	nand2_1 U5916( .A(n6033), .B(n6017), .Y(n6057) );
	o221ai_1 U5917( .A1(n6045), .A2(n15043), .B1(n5353), .B2(n15041), .C1(n6062), .Y(n6017) );
	nand2_1 U5918( .A(g2439), .B(g5747), .Y(n6062) );
	a21oi_1 U5919( .A1(n6022), .A2(n6021), .B1(n6033), .Y(n6056) );
	inv_1 U5920( .A(n6047), .Y(n6033) );
	o221ai_1 U5921( .A1(n6045), .A2(n15039), .B1(n5353), .B2(n15038), .C1(n6063), .Y(n6047) );
	nand2_1 U5922( .A(g2454), .B(g5747), .Y(n6063) );
	o221ai_1 U5923( .A1(n6045), .A2(n15035), .B1(n5353), .B2(n15034), .C1(n6064), .Y(n6022) );
	nand2_1 U5924( .A(g5747), .B(g2469), .Y(n6064) );
	o22ai_1 U5925( .A1(n5986), .A2(n5607), .B1(n5987), .B2(n6065), .Y(n5195) );
	o22ai_1 U5926( .A1(n5989), .A2(n5593), .B1(n5990), .B2(n6065), .Y(n5194) );
	o22ai_1 U5927( .A1(n5992), .A2(n5402), .B1(n5993), .B2(n6065), .Y(n5193) );
	nand2_1 U5928( .A(n6005), .B(n5999), .Y(n6065) );
	o211ai_1 U5929( .A1(n6066), .A2(n5402), .B1(n6067), .C1(n6068), .Y(n6005) );
	a22oi_1 U5930( .A1(n9874), .A2(g7390), .B1(n9873), .B2(n7224), .Y(n6068) );
	nand3_1 U5931( .A(n7256), .B(n6069), .C(g2616), .Y(n6067) );
	o22ai_1 U5932( .A1(n5986), .A2(n5608), .B1(n5987), .B2(n6070), .Y(n5192) );
	o22ai_1 U5933( .A1(n5989), .A2(n5594), .B1(n5990), .B2(n6070), .Y(n5191) );
	inv_1 U5934( .A(n59), .Y(n5990) );
	nand2_1 U5935( .A(n6071), .B(n5749), .Y(n5989) );
	o22ai_1 U5936( .A1(n5992), .A2(n5403), .B1(n5993), .B2(n6070), .Y(n5190) );
	nand2_1 U5937( .A(n6004), .B(n5999), .Y(n6070) );
	o211ai_1 U5938( .A1(n6066), .A2(n5403), .B1(n6072), .C1(n6073), .Y(n6004) );
	a22oi_1 U5939( .A1(n9876), .A2(g7390), .B1(n9875), .B2(n7224), .Y(n6073) );
	nand3_1 U5940( .A(g2598), .B(n6074), .C(n7256), .Y(n6072) );
	inv_1 U5941( .A(n58), .Y(n5993) );
	nor2_1 U5942( .A(n6066), .B(RST), .Y(n58) );
	nand2_1 U5943( .A(n5755), .B(n6066), .Y(n5992) );
	o22ai_1 U5944( .A1(n6075), .A2(n6076), .B1(n6077), .B2(n6078), .Y(n5189) );
	inv_1 U5945( .A(n7349), .Y(n6078) );
	o22ai_1 U5946( .A1(n6075), .A2(n6079), .B1(n6080), .B2(n6081), .Y(n5188) );
	inv_1 U5947( .A(n7350), .Y(n6081) );
	o22ai_1 U5948( .A1(n6075), .A2(n6082), .B1(n6083), .B2(n5504), .Y(n5187) );
	o21ai_0 U5949( .A1(n6023), .A2(n6084), .B1(n5753), .Y(n6075) );
	nand2_1 U5950( .A(n6030), .B(n6032), .Y(n6023) );
	o22ai_1 U5951( .A1(n6076), .A2(n6085), .B1(n6077), .B2(n6086), .Y(n5186) );
	inv_1 U5952( .A(n7343), .Y(n6086) );
	o22ai_1 U5953( .A1(n6079), .A2(n6085), .B1(n6080), .B2(n6087), .Y(n5185) );
	inv_1 U5954( .A(n7344), .Y(n6087) );
	o22ai_1 U5955( .A1(n6082), .A2(n6085), .B1(n6083), .B2(n5503), .Y(n5184) );
	o221ai_1 U5956( .A1(n6032), .A2(n6088), .B1(n6089), .B2(n6090), .C1(n5743), .Y(n6085) );
	inv_1 U5957( .A(n6025), .Y(n6090) );
	nor2_1 U5958( .A(n6053), .B(n6061), .Y(n6025) );
	mux2i_1 U5959( .A0(n5984), .A1(n5983), .S(n6021), .Y(n6088) );
	o22ai_1 U5960( .A1(n6076), .A2(n6091), .B1(n6077), .B2(n6092), .Y(n5183) );
	inv_1 U5961( .A(n7345), .Y(n6092) );
	o22ai_1 U5962( .A1(n6079), .A2(n6091), .B1(n6080), .B2(n6093), .Y(n5182) );
	inv_1 U5963( .A(n7346), .Y(n6093) );
	o22ai_1 U5964( .A1(n6082), .A2(n6091), .B1(n6083), .B2(n5502), .Y(n5181) );
	o211ai_1 U5965( .A1(n6030), .A2(n6089), .B1(n6018), .C1(n5740), .Y(n6091) );
	inv_1 U5966( .A(n6084), .Y(n6089) );
	xnor2_1 U5967( .A(n6042), .B(n5983), .Y(n6084) );
	inv_1 U5968( .A(n6021), .Y(n6042) );
	o22ai_1 U5969( .A1(n6076), .A2(n6094), .B1(n6077), .B2(n6095), .Y(n5180) );
	inv_1 U5970( .A(n7347), .Y(n6095) );
	nand2_1 U5971( .A(n6076), .B(n5748), .Y(n6077) );
	nand2_1 U5972( .A(n7224), .B(n6096), .Y(n6076) );
	o22ai_1 U5973( .A1(n6079), .A2(n6094), .B1(n6080), .B2(n6097), .Y(n5179) );
	inv_1 U5974( .A(n7348), .Y(n6097) );
	nand2_1 U5975( .A(n6079), .B(n5748), .Y(n6080) );
	nand2_1 U5976( .A(g7390), .B(n6096), .Y(n6079) );
	o22ai_1 U5977( .A1(n6082), .A2(n6094), .B1(n6083), .B2(n5501), .Y(n5178) );
	nand2_1 U5978( .A(n6082), .B(n5748), .Y(n6083) );
	o221ai_1 U5979( .A1(n6098), .A2(n6015), .B1(g3229), .B2(n6018), .C1(n6099), .Y(n6094) );
	a21oi_1 U5980( .A1(n6100), .A2(n6021), .B1(RST), .Y(n6099) );
	o221ai_1 U5981( .A1(n7348), .A2(n6071), .B1(n7347), .B2(n6101), .C1(n6102), .Y(n6021) );
	nand2_1 U5982( .A(g7302), .B(n5501), .Y(n6102) );
	o22ai_1 U5983( .A1(n6030), .A2(n5983), .B1(n6103), .B2(n6053), .Y(n6100) );
	nor2_1 U5984( .A(n6032), .B(n5983), .Y(n6103) );
	inv_1 U5985( .A(n6041), .Y(n6030) );
	inv_1 U5986( .A(n6054), .Y(n6018) );
	nor2_1 U5987( .A(n6041), .B(n6032), .Y(n6054) );
	inv_1 U5988( .A(n6061), .Y(n6032) );
	o221ai_1 U5989( .A1(n7346), .A2(n6071), .B1(n7345), .B2(n6101), .C1(n6104), .Y(n6061) );
	nand2_1 U5990( .A(g7302), .B(n5502), .Y(n6104) );
	o221ai_1 U5991( .A1(n7344), .A2(n6071), .B1(n7343), .B2(n6101), .C1(n6105), .Y(n6041) );
	nand2_1 U5992( .A(g7302), .B(n5503), .Y(n6105) );
	inv_1 U5993( .A(n6053), .Y(n6015) );
	o221ai_1 U5994( .A1(n7350), .A2(n6071), .B1(n7349), .B2(n6101), .C1(n6106), .Y(n6053) );
	nand2_1 U5995( .A(g7302), .B(n5504), .Y(n6106) );
	nand2_1 U5996( .A(g7302), .B(n6096), .Y(n6082) );
	and2_0 U5997( .A(g2632), .B(n5759), .X(n5177) );
	and2_0 U5998( .A(g2617), .B(n5759), .X(n5176) );
	o22ai_1 U5999( .A1(n6107), .A2(n6108), .B1(n6109), .B2(n5643), .Y(n5175) );
	o22ai_1 U6000( .A1(n6107), .A2(n5787), .B1(n6110), .B2(n6111), .Y(n5174) );
	inv_1 U6001( .A(n7459), .Y(n6111) );
	o22ai_1 U6002( .A1(n6107), .A2(n5788), .B1(n6112), .B2(n5416), .Y(n5173) );
	o22ai_1 U6003( .A1(n6108), .A2(n6113), .B1(n6109), .B2(n5644), .Y(n5172) );
	o22ai_1 U6004( .A1(n5787), .A2(n6113), .B1(n6110), .B2(n6114), .Y(n5171) );
	inv_1 U6005( .A(n7453), .Y(n6114) );
	o22ai_1 U6006( .A1(n5788), .A2(n6113), .B1(n6112), .B2(n5417), .Y(n5170) );
	o22ai_1 U6007( .A1(n6115), .A2(n6108), .B1(n6109), .B2(n5645), .Y(n5169) );
	or2_0 U6008( .A(RST), .B(n7260), .X(n6109) );
	o22ai_1 U6009( .A1(n6115), .A2(n5787), .B1(n6110), .B2(n6116), .Y(n5168) );
	inv_1 U6010( .A(n7451), .Y(n6116) );
	or2_0 U6011( .A(RST), .B(g8167), .X(n6110) );
	o22ai_1 U6012( .A1(n6115), .A2(n5788), .B1(n6112), .B2(n5415), .Y(n5167) );
	or2_0 U6013( .A(RST), .B(g8087), .X(n6112) );
	and2_0 U6014( .A(g2642), .B(n5759), .X(n5166) );
	and2_0 U6015( .A(g2648), .B(n5744), .X(n5165) );
	and2_0 U6016( .A(g2646), .B(n5759), .X(n5164) );
	and2_0 U6017( .A(g2638), .B(n5759), .X(n5163) );
	o22ai_1 U6018( .A1(n5982), .A2(n5986), .B1(n5987), .B2(n6117), .Y(n5162) );
	o22ai_1 U6019( .A1(n5986), .A2(n6117), .B1(n9960), .B2(n5987), .Y(n5161) );
	inv_1 U6020( .A(n7290), .Y(n6117) );
	o22ai_1 U6021( .A1(n5986), .A2(n5589), .B1(n6118), .B2(n5987), .Y(n5160) );
	nand2_1 U6022( .A(n7224), .B(n5748), .Y(n5987) );
	nand2_1 U6023( .A(n6101), .B(n5748), .Y(n5986) );
	nor2_1 U6024( .A(RST), .B(n6045), .Y(n5159) );
	inv_1 U6025( .A(g5796), .Y(n6045) );
	and2_0 U6026( .A(g2472), .B(n5758), .X(n5158) );
	and2_0 U6027( .A(g2470), .B(n5758), .X(n5157) );
	and2_0 U6028( .A(g2457), .B(n5758), .X(n5156) );
	and2_0 U6029( .A(g2455), .B(n5758), .X(n5155) );
	and2_0 U6030( .A(g2442), .B(n5758), .X(n5154) );
	and2_0 U6031( .A(g2440), .B(n5758), .X(n5153) );
	and2_0 U6032( .A(g2427), .B(n5750), .X(n5152) );
	and2_0 U6033( .A(g2425), .B(n5743), .X(n5151) );
	a221oi_1 U6034( .A1(n6119), .A2(n6120), .B1(n6121), .B2(n6122), .C1(RST), .Y(n5150) );
	nor4_1 U6035( .A(n6123), .B(n6124), .C(n6125), .D(n6126), .Y(n6120) );
	xnor2_1 U6036( .A(n7709), .B(n6127), .Y(n6126) );
	xnor2_1 U6037( .A(n10051), .B(n6128), .Y(n6125) );
	xnor2_1 U6038( .A(n7705), .B(n6129), .Y(n6124) );
	nand3_1 U6039( .A(n6130), .B(n6131), .C(n6132), .Y(n6123) );
	xor2_1 U6040( .A(n10059), .B(n6133), .X(n6132) );
	nor4_1 U6041( .A(n6134), .B(n6135), .C(n6136), .D(n6137), .Y(n6119) );
	xnor2_1 U6042( .A(n7307), .B(n6138), .Y(n6137) );
	xnor2_1 U6043( .A(n7699), .B(n6139), .Y(n6136) );
	xnor2_1 U6044( .A(n10062), .B(n6140), .Y(n6135) );
	nand3_1 U6045( .A(n6141), .B(n6142), .C(n6143), .Y(n6134) );
	xnor2_1 U6046( .A(n10060), .B(n6144), .Y(n6143) );
	xnor2_1 U6047( .A(n10061), .B(n6145), .Y(n6142) );
	xnor2_1 U6048( .A(n7696), .B(n6146), .Y(n6141) );
	mux2i_1 U6049( .A0(n6147), .A1(n6148), .S(n7743), .Y(n5149) );
	a22oi_1 U6050( .A1(n6149), .A2(n7632), .B1(n48), .B2(n6150), .Y(n6148) );
	nand2_1 U6051( .A(n5756), .B(n14920), .Y(n6147) );
	nor2_1 U6052( .A(RST), .B(n6151), .Y(n5148) );
	and2_0 U6053( .A(g2365), .B(n5744), .X(n5147) );
	o22ai_1 U6054( .A1(n6152), .A2(n6153), .B1(n6154), .B2(n6155), .Y(n5146) );
	inv_1 U6055( .A(n7382), .Y(n6155) );
	nor2_1 U6056( .A(n6156), .B(n6157), .Y(n6154) );
	o22ai_1 U6057( .A1(n6158), .A2(n6153), .B1(n6159), .B2(n6160), .Y(n5145) );
	inv_1 U6058( .A(n7381), .Y(n6160) );
	nor2_1 U6059( .A(n6156), .B(n6149), .Y(n6159) );
	o22ai_1 U6060( .A1(n6153), .A2(n6161), .B1(n6162), .B2(n6163), .Y(n5144) );
	nor2_1 U6061( .A(n6156), .B(n6164), .Y(n6162) );
	and2_0 U6062( .A(n6165), .B(n5749), .X(n6156) );
	nand2_1 U6063( .A(n7264), .B(n6165), .Y(n6153) );
	or3_1 U6064( .A(n6166), .B(n6167), .C(n6168), .X(n6165) );
	o22ai_1 U6065( .A1(n6152), .A2(n6169), .B1(n6170), .B2(n6171), .Y(n5143) );
	nor2_1 U6066( .A(n6172), .B(n6157), .Y(n6170) );
	o22ai_1 U6067( .A1(n6158), .A2(n6169), .B1(n6173), .B2(n6174), .Y(n5142) );
	nor2_1 U6068( .A(n6172), .B(n6149), .Y(n6173) );
	o22ai_1 U6069( .A1(n6161), .A2(n6169), .B1(n6175), .B2(n6176), .Y(n5141) );
	inv_1 U6070( .A(n7726), .Y(n6176) );
	nor2_1 U6071( .A(n6172), .B(n6164), .Y(n6175) );
	a21oi_1 U6072( .A1(n6177), .A2(n6178), .B1(RST), .Y(n6172) );
	inv_1 U6073( .A(n6179), .Y(n6177) );
	o21ai_0 U6074( .A1(n6179), .A2(n6166), .B1(n6180), .Y(n6169) );
	mux2i_1 U6075( .A0(n6168), .A1(n6181), .S(n6113), .Y(n6180) );
	a21oi_1 U6076( .A1(n6182), .A2(n7264), .B1(n6183), .Y(n6179) );
	and4_1 U6077( .A(n6184), .B(n6185), .C(n6186), .D(n6187), .X(n6183) );
	o22ai_1 U6078( .A1(n6188), .A2(n6189), .B1(n6152), .B2(n6190), .Y(n5140) );
	o22ai_1 U6079( .A1(n6191), .A2(n6192), .B1(n6158), .B2(n6190), .Y(n5139) );
	inv_1 U6080( .A(n7573), .Y(n6192) );
	o22ai_1 U6081( .A1(n6193), .A2(n5609), .B1(n6161), .B2(n6190), .Y(n5138) );
	nand2_1 U6082( .A(n6194), .B(n6195), .Y(n6190) );
	mux2i_1 U6083( .A0(n6196), .A1(n6197), .S(n6198), .Y(n6194) );
	nand2_1 U6084( .A(n6187), .B(n6197), .Y(n6196) );
	o211ai_1 U6085( .A1(n6184), .A2(n6199), .B1(n6187), .C1(n6200), .Y(n6197) );
	mux2i_1 U6086( .A0(n6201), .A1(n6202), .S(n6203), .Y(n6200) );
	a21oi_1 U6087( .A1(n6204), .A2(n6205), .B1(n6206), .Y(n6202) );
	nand2_1 U6088( .A(n6184), .B(n6186), .Y(n6205) );
	nand3_1 U6089( .A(n6184), .B(n6185), .C(n7264), .Y(n6201) );
	inv_1 U6090( .A(n6181), .Y(n6199) );
	nand2_1 U6091( .A(n6204), .B(n6186), .Y(n6181) );
	o22ai_1 U6092( .A1(n6188), .A2(n6207), .B1(n6152), .B2(n6208), .Y(n5137) );
	o22ai_1 U6093( .A1(n6191), .A2(n6209), .B1(n6158), .B2(n6208), .Y(n5136) );
	inv_1 U6094( .A(n7575), .Y(n6209) );
	o22ai_1 U6095( .A1(n6193), .A2(n5610), .B1(n6161), .B2(n6208), .Y(n5135) );
	nand2_1 U6096( .A(n6210), .B(n6195), .Y(n6208) );
	xnor2_1 U6097( .A(n6211), .B(n6212), .Y(n6210) );
	a21oi_1 U6098( .A1(n6213), .A2(n6187), .B1(n6121), .Y(n6212) );
	o22ai_1 U6099( .A1(n6214), .A2(n6215), .B1(n6216), .B2(n6203), .Y(n6213) );
	a21oi_1 U6100( .A1(n6217), .A2(n6178), .B1(n6206), .Y(n6216) );
	a21oi_1 U6101( .A1(n6218), .A2(n6184), .B1(n6219), .Y(n6217) );
	inv_1 U6102( .A(n6185), .Y(n6218) );
	mux2i_1 U6103( .A0(n6220), .A1(n6221), .S(n6203), .Y(n6215) );
	o21ai_0 U6104( .A1(n6198), .A2(n6222), .B1(n6223), .Y(n6221) );
	inv_1 U6105( .A(n6224), .Y(n6223) );
	and2_0 U6106( .A(n6222), .B(n6184), .X(n6220) );
	nand2_1 U6107( .A(n6225), .B(n6186), .Y(n6222) );
	nand4_1 U6108( .A(n6226), .B(n6227), .C(n6228), .D(n6229), .Y(n6186) );
	nor3_1 U6109( .A(n6230), .B(n6231), .C(n6232), .Y(n6229) );
	or3_1 U6110( .A(n6233), .B(n6234), .C(n6235), .X(n6230) );
	nor3_1 U6111( .A(n6236), .B(n6237), .C(n6238), .Y(n6228) );
	inv_1 U6112( .A(n6239), .Y(n6225) );
	o22ai_1 U6113( .A1(n6188), .A2(n6240), .B1(n6152), .B2(n6241), .Y(n5134) );
	o22ai_1 U6114( .A1(n6191), .A2(n6242), .B1(n6158), .B2(n6241), .Y(n5133) );
	inv_1 U6115( .A(n7571), .Y(n6242) );
	o22ai_1 U6116( .A1(n6193), .A2(n5611), .B1(n6161), .B2(n6241), .Y(n5132) );
	o21ai_0 U6117( .A1(n6243), .A2(n6244), .B1(n6195), .Y(n6241) );
	nor3_1 U6118( .A(n6185), .B(n6245), .C(n6182), .Y(n6244) );
	o22ai_1 U6119( .A1(n6152), .A2(n6246), .B1(n6247), .B2(n6248), .Y(n5131) );
	inv_1 U6120( .A(n7310), .Y(n6248) );
	nor2_1 U6121( .A(n6249), .B(n6157), .Y(n6247) );
	o22ai_1 U6122( .A1(n6158), .A2(n6246), .B1(n6250), .B2(n6251), .Y(n5130) );
	inv_1 U6123( .A(n7309), .Y(n6251) );
	nor2_1 U6124( .A(n6249), .B(n6149), .Y(n6250) );
	o22ai_1 U6125( .A1(n6161), .A2(n6246), .B1(n6252), .B2(n6253), .Y(n5129) );
	nor2_1 U6126( .A(n6249), .B(n6164), .Y(n6252) );
	a21oi_1 U6127( .A1(n6254), .A2(n6255), .B1(RST), .Y(n6249) );
	inv_1 U6128( .A(n6256), .Y(n6255) );
	o211ai_1 U6129( .A1(n6115), .A2(n6257), .B1(n7264), .C1(n6258), .Y(n6246) );
	mux2i_1 U6130( .A0(n6115), .A1(n6257), .S(n6259), .Y(n6258) );
	o22ai_1 U6131( .A1(n5548), .A2(n6188), .B1(n6152), .B2(n6260), .Y(n5128) );
	o22ai_1 U6132( .A1(n5338), .A2(n6191), .B1(n6158), .B2(n6260), .Y(n5127) );
	o22ai_1 U6133( .A1(n6261), .A2(n6193), .B1(n6161), .B2(n6260), .Y(n5126) );
	xnor2_1 U6134( .A(n6262), .B(n6115), .Y(n6260) );
	inv_1 U6135( .A(n6263), .Y(n6115) );
	nand2_1 U6136( .A(n6254), .B(n6256), .Y(n6262) );
	o221ai_1 U6137( .A1(n7309), .A2(n6264), .B1(n7310), .B2(n6265), .C1(n6266), .Y(n6256) );
	nand2_1 U6138( .A(g5555), .B(n6253), .Y(n6266) );
	inv_1 U6139( .A(n7713), .Y(n6253) );
	and2_0 U6140( .A(n6267), .B(n7264), .X(n6254) );
	mux2i_1 U6141( .A0(n6268), .A1(n6269), .S(n6259), .Y(n6267) );
	nand2_1 U6142( .A(n6257), .B(n6263), .Y(n6269) );
	or2_0 U6143( .A(n6263), .B(n6257), .X(n6268) );
	o221ai_1 U6144( .A1(n6264), .A2(n5338), .B1(n6265), .B2(n5548), .C1(n6270), .Y(n6263) );
	nand2_1 U6145( .A(n7617), .B(g5555), .Y(n6270) );
	inv_1 U6146( .A(n7617), .Y(n6261) );
	o22ai_1 U6147( .A1(n6188), .A2(n5612), .B1(n6152), .B2(n6271), .Y(n5125) );
	o22ai_1 U6148( .A1(n6191), .A2(n5380), .B1(n6158), .B2(n6271), .Y(n5124) );
	o22ai_1 U6149( .A1(n6193), .A2(n6272), .B1(n6161), .B2(n6271), .Y(n5123) );
	mux2_1 U6150( .A0(n6259), .A1(n6257), .S(n7264), .X(n6271) );
	o21ai_0 U6151( .A1(n6273), .A2(n6274), .B1(n6275), .Y(n6257) );
	inv_1 U6152( .A(n6276), .Y(n6275) );
	o22ai_1 U6153( .A1(n9961), .A2(n6277), .B1(n7383), .B2(n6278), .Y(n6274) );
	nor2_1 U6154( .A(n7384), .B(n6279), .Y(n6273) );
	a21oi_1 U6155( .A1(n7780), .A2(n10052), .B1(n6280), .Y(n6259) );
	o22ai_1 U6156( .A1(n6272), .A2(n6281), .B1(n5380), .B2(n6264), .Y(n6280) );
	inv_1 U6157( .A(n7628), .Y(n6272) );
	o22ai_1 U6158( .A1(n6152), .A2(n6282), .B1(n6283), .B2(n6284), .Y(n5122) );
	inv_1 U6159( .A(n7336), .Y(n6284) );
	nor2_1 U6160( .A(n6285), .B(n6157), .Y(n6283) );
	o22ai_1 U6161( .A1(n6158), .A2(n6282), .B1(n6286), .B2(n6287), .Y(n5121) );
	inv_1 U6162( .A(n7335), .Y(n6287) );
	nor2_1 U6163( .A(n6285), .B(n6149), .Y(n6286) );
	o22ai_1 U6164( .A1(n6161), .A2(n6282), .B1(n6288), .B2(n6289), .Y(n5120) );
	nor2_1 U6165( .A(n6285), .B(n6164), .Y(n6288) );
	a21oi_1 U6166( .A1(n6290), .A2(n6291), .B1(RST), .Y(n6285) );
	o22ai_1 U6167( .A1(n5549), .A2(n6188), .B1(n6292), .B2(n6152), .Y(n5119) );
	o22ai_1 U6168( .A1(n5339), .A2(n6191), .B1(n6292), .B2(n6158), .Y(n5118) );
	o22ai_1 U6169( .A1(n6293), .A2(n6193), .B1(n6292), .B2(n6161), .Y(n5117) );
	xnor2_1 U6170( .A(n6151), .B(n6294), .Y(n6292) );
	a21oi_1 U6171( .A1(n6206), .A2(n6295), .B1(n6296), .Y(n6294) );
	nor4_1 U6172( .A(n6297), .B(n6291), .C(n6168), .D(n6298), .Y(n6296) );
	inv_1 U6173( .A(n6299), .Y(n6291) );
	inv_1 U6174( .A(n7677), .Y(n6293) );
	o22ai_1 U6175( .A1(n6300), .A2(n6152), .B1(n6188), .B2(n5666), .Y(n5116) );
	inv_1 U6176( .A(n6157), .Y(n6188) );
	nor2_1 U6177( .A(n7780), .B(RST), .Y(n6157) );
	nand2_1 U6178( .A(n7780), .B(n5747), .Y(n6152) );
	o22ai_1 U6179( .A1(n6300), .A2(n6158), .B1(n6191), .B2(n5667), .Y(n5115) );
	inv_1 U6180( .A(n6149), .Y(n6191) );
	nor2_1 U6181( .A(g7264), .B(RST), .Y(n6149) );
	inv_1 U6182( .A(n48), .Y(n6158) );
	o22ai_1 U6183( .A1(n6300), .A2(n6161), .B1(n6193), .B2(n6301), .Y(n5114) );
	inv_1 U6184( .A(n6164), .Y(n6193) );
	nor2_1 U6185( .A(g5555), .B(RST), .Y(n6164) );
	inv_1 U6186( .A(n3960), .Y(n6161) );
	xnor2_1 U6187( .A(n6297), .B(n6302), .Y(n6300) );
	a21oi_1 U6188( .A1(n6303), .A2(n7264), .B1(n6304), .Y(n6302) );
	inv_1 U6189( .A(n6282), .Y(n6304) );
	nand2_1 U6190( .A(n6297), .B(n6290), .Y(n6282) );
	o32ai_1 U6191( .A1(n6168), .A2(n6151), .A3(n6305), .B1(n6206), .B2(n6306), .Y(n6290) );
	inv_1 U6192( .A(n6295), .Y(n6306) );
	nor3_1 U6193( .A(n6168), .B(n6107), .C(n6307), .Y(n6295) );
	inv_1 U6194( .A(n6305), .Y(n6307) );
	inv_1 U6195( .A(n7264), .Y(n6168) );
	a21oi_1 U6196( .A1(n6308), .A2(n6309), .B1(n6297), .Y(n6303) );
	inv_1 U6197( .A(n6298), .Y(n6309) );
	xnor2_1 U6198( .A(n6305), .B(n6107), .Y(n6298) );
	nor3_1 U6199( .A(n6310), .B(n6311), .C(n6276), .Y(n6305) );
	a21oi_1 U6200( .A1(n6206), .A2(n6151), .B1(n6299), .Y(n6308) );
	o221ai_1 U6201( .A1(n7335), .A2(n6264), .B1(n7336), .B2(n6265), .C1(n6312), .Y(n6299) );
	nand2_1 U6202( .A(g5555), .B(n6289), .Y(n6312) );
	inv_1 U6203( .A(n7732), .Y(n6289) );
	inv_1 U6204( .A(n6107), .Y(n6151) );
	o221ai_1 U6205( .A1(n6264), .A2(n5339), .B1(n6265), .B2(n5549), .C1(n6313), .Y(n6107) );
	nand2_1 U6206( .A(n7677), .B(g5555), .Y(n6313) );
	a221oi_1 U6207( .A1(g7264), .A2(n9889), .B1(n7780), .B2(n10058), .C1(n6314), .Y(n6297) );
	nor2_1 U6208( .A(n6301), .B(n6281), .Y(n6314) );
	inv_1 U6209( .A(n7624), .Y(n6301) );
	and2_0 U6210( .A(g5637), .B(n5759), .X(n5113) );
	nor2_1 U6211( .A(n6315), .B(n6316), .Y(n5112) );
	xnor2_1 U6212( .A(n10059), .B(n6317), .Y(n6315) );
	nor2_1 U6213( .A(n6318), .B(n6319), .Y(n6317) );
	nor2_1 U6214( .A(n6320), .B(n6316), .Y(n5111) );
	xnor2_1 U6215( .A(n6319), .B(n6318), .Y(n6320) );
	inv_1 U6216( .A(n7307), .Y(n6318) );
	nand2_1 U6217( .A(n6321), .B(n7705), .Y(n6319) );
	nor2_1 U6218( .A(n6322), .B(n6316), .Y(n5110) );
	xnor2_1 U6219( .A(n7705), .B(n6321), .Y(n6322) );
	a211oi_1 U6220( .A1(n5371), .A2(n6323), .B1(n6316), .C1(n6321), .Y(n5109) );
	nor2_1 U6221( .A(n6323), .B(n5371), .Y(n6321) );
	nor3_1 U6222( .A(n6316), .B(n6324), .C(n6325), .Y(n5108) );
	a21oi_1 U6223( .A1(n6326), .A2(n10061), .B1(n7696), .Y(n6325) );
	inv_1 U6224( .A(n6323), .Y(n6324) );
	nand3_1 U6225( .A(n7696), .B(n10061), .C(n6326), .Y(n6323) );
	nor2_1 U6226( .A(n6327), .B(n6316), .Y(n5107) );
	xnor2_1 U6227( .A(n10061), .B(n6326), .Y(n6327) );
	a211oi_1 U6228( .A1(n6328), .A2(n6329), .B1(n6316), .C1(n6326), .Y(n5106) );
	nor2_1 U6229( .A(n6329), .B(n6328), .Y(n6326) );
	inv_1 U6230( .A(n6330), .Y(n6329) );
	inv_1 U6231( .A(n7709), .Y(n6328) );
	a211oi_1 U6232( .A1(n5372), .A2(n6331), .B1(n6316), .C1(n6330), .Y(n5105) );
	nor2_1 U6233( .A(n6331), .B(n5372), .Y(n6330) );
	nor3_1 U6234( .A(n6316), .B(n6332), .C(n6333), .Y(n5104) );
	a21oi_1 U6235( .A1(n6334), .A2(n10051), .B1(n7699), .Y(n6333) );
	inv_1 U6236( .A(n6331), .Y(n6332) );
	nand3_1 U6237( .A(n7699), .B(n10051), .C(n6334), .Y(n6331) );
	nor2_1 U6238( .A(n6335), .B(n6316), .Y(n5103) );
	o21ai_0 U6239( .A1(n6336), .A2(n6131), .B1(n5746), .Y(n6316) );
	xnor2_1 U6240( .A(n6334), .B(n10051), .Y(n6335) );
	nor2_1 U6241( .A(n6277), .B(n6337), .Y(n6334) );
	o22ai_1 U6242( .A1(n6338), .A2(n6339), .B1(n6340), .B2(n6341), .Y(n5102) );
	inv_1 U6243( .A(n7673), .Y(n6338) );
	o22ai_1 U6244( .A1(n5331), .A2(n6342), .B1(n6340), .B2(n6343), .Y(n5101) );
	o22ai_1 U6245( .A1(n5547), .A2(n6344), .B1(n6340), .B2(n6345), .Y(n5100) );
	o221ai_1 U6246( .A1(n6346), .A2(n6347), .B1(n6348), .B2(n6349), .C1(n6350), .Y(n6340) );
	xor2_1 U6247( .A(n6351), .B(n6133), .X(n6346) );
	nand2_1 U6248( .A(n6352), .B(n6353), .Y(n6351) );
	xnor2_1 U6249( .A(n6138), .B(n6354), .Y(n6353) );
	inv_1 U6250( .A(n6355), .Y(n51) );
	o22ai_1 U6251( .A1(n6356), .A2(n6339), .B1(n6357), .B2(n6341), .Y(n5099) );
	o22ai_1 U6252( .A1(n5519), .A2(n6342), .B1(n6357), .B2(n6343), .Y(n5098) );
	o22ai_1 U6253( .A1(n5693), .A2(n6344), .B1(n6357), .B2(n6345), .Y(n5097) );
	a221oi_1 U6254( .A1(n6358), .A2(n6359), .B1(n6354), .B2(n6360), .C1(n6361), .Y(n6357) );
	nor2_1 U6255( .A(n6362), .B(n6347), .Y(n6361) );
	xnor2_1 U6256( .A(n6352), .B(n6363), .Y(n6362) );
	and2_0 U6257( .A(n6364), .B(n6365), .X(n6352) );
	mux2i_1 U6258( .A0(n6366), .A1(n6367), .S(n6144), .Y(n6364) );
	nand2_1 U6259( .A(n6243), .B(n6368), .Y(n6367) );
	nand2_1 U6260( .A(n6129), .B(n6354), .Y(n6366) );
	o22ai_1 U6261( .A1(n6369), .A2(n6339), .B1(n6370), .B2(n6341), .Y(n5096) );
	o22ai_1 U6262( .A1(n5521), .A2(n6342), .B1(n6370), .B2(n6343), .Y(n5095) );
	o22ai_1 U6263( .A1(n5694), .A2(n6344), .B1(n6370), .B2(n6345), .Y(n5094) );
	inv_1 U6264( .A(n6371), .Y(n6370) );
	o22ai_1 U6265( .A1(n5836), .A2(n6349), .B1(n6347), .B2(n6372), .Y(n6371) );
	xnor2_1 U6266( .A(n6129), .B(n6373), .Y(n6372) );
	nand2_1 U6267( .A(n6365), .B(n6374), .Y(n6373) );
	xnor2_1 U6268( .A(n6144), .B(n6243), .Y(n6374) );
	o22ai_1 U6269( .A1(n6375), .A2(n6339), .B1(n6376), .B2(n6341), .Y(n5093) );
	o22ai_1 U6270( .A1(n5522), .A2(n6342), .B1(n6376), .B2(n6343), .Y(n5092) );
	o22ai_1 U6271( .A1(n5695), .A2(n6344), .B1(n6376), .B2(n6345), .Y(n5091) );
	inv_1 U6272( .A(n6377), .Y(n6376) );
	o22ai_1 U6273( .A1(n5834), .A2(n6349), .B1(n6347), .B2(n6378), .Y(n6377) );
	xnor2_1 U6274( .A(n6365), .B(n6144), .Y(n6378) );
	and2_0 U6275( .A(n6379), .B(n6380), .X(n6365) );
	xnor2_1 U6276( .A(n6146), .B(n6243), .Y(n6380) );
	o22ai_1 U6277( .A1(n6381), .A2(n6339), .B1(n6341), .B2(n6382), .Y(n5090) );
	o22ai_1 U6278( .A1(n5720), .A2(n6342), .B1(n6343), .B2(n6382), .Y(n5089) );
	o22ai_1 U6279( .A1(n5679), .A2(n6344), .B1(n6345), .B2(n6382), .Y(n5088) );
	nand2_1 U6280( .A(n6383), .B(n6384), .Y(n6382) );
	mux2i_1 U6281( .A0(n6385), .A1(n5832), .S(n6347), .Y(n6383) );
	xnor2_1 U6282( .A(n6146), .B(n6379), .Y(n6385) );
	nor2_1 U6283( .A(n6386), .B(n6387), .Y(n6379) );
	xnor2_1 U6284( .A(n6145), .B(n6354), .Y(n6386) );
	o22ai_1 U6285( .A1(n6388), .A2(n6339), .B1(n6389), .B2(n6341), .Y(n5087) );
	o22ai_1 U6286( .A1(n5721), .A2(n6342), .B1(n6389), .B2(n6343), .Y(n5086) );
	o22ai_1 U6287( .A1(n5680), .A2(n6344), .B1(n6389), .B2(n6345), .Y(n5085) );
	inv_1 U6288( .A(n6390), .Y(n6389) );
	o22ai_1 U6289( .A1(n5830), .A2(n6349), .B1(n6391), .B2(n6347), .Y(n6390) );
	xor2_1 U6290( .A(n6145), .B(n6387), .X(n6391) );
	a22oi_1 U6291( .A1(n6392), .A2(n6393), .B1(n6127), .B2(n6394), .Y(n6387) );
	o22ai_1 U6292( .A1(n6395), .A2(n6339), .B1(n6341), .B2(n6396), .Y(n5084) );
	inv_1 U6293( .A(n7667), .Y(n6395) );
	o22ai_1 U6294( .A1(n5738), .A2(n6342), .B1(n6343), .B2(n6396), .Y(n5083) );
	o22ai_1 U6295( .A1(n5542), .A2(n6344), .B1(n6345), .B2(n6396), .Y(n5082) );
	o221ai_1 U6296( .A1(n6347), .A2(n6397), .B1(n7235), .B2(n6349), .C1(n6350), .Y(n6396) );
	xor2_1 U6297( .A(n6127), .B(n6398), .X(n6397) );
	a21oi_1 U6298( .A1(n6399), .A2(n6393), .B1(n6394), .Y(n6398) );
	nor3_1 U6299( .A(n6400), .B(n6243), .C(n6401), .Y(n6394) );
	inv_1 U6300( .A(n6401), .Y(n6393) );
	nor2_1 U6301( .A(n6140), .B(n6354), .Y(n6399) );
	o22ai_1 U6302( .A1(n6402), .A2(n6339), .B1(n6403), .B2(n6341), .Y(n5081) );
	o22ai_1 U6303( .A1(n5523), .A2(n6342), .B1(n6403), .B2(n6343), .Y(n5080) );
	o22ai_1 U6304( .A1(n5696), .A2(n6344), .B1(n6403), .B2(n6345), .Y(n5079) );
	inv_1 U6305( .A(n6404), .Y(n6403) );
	o221ai_1 U6306( .A1(n6347), .A2(n6405), .B1(n6243), .B2(n6384), .C1(n6406), .Y(n6404) );
	nand2_1 U6307( .A(n6359), .B(n7250), .Y(n6406) );
	inv_1 U6308( .A(n6349), .Y(n6359) );
	xnor2_1 U6309( .A(n6140), .B(n6401), .Y(n6405) );
	o211ai_1 U6310( .A1(n6128), .A2(n6407), .B1(n6408), .C1(n6409), .Y(n6401) );
	mux2i_1 U6311( .A0(n6128), .A1(n6407), .S(n6354), .Y(n6409) );
	o22ai_1 U6312( .A1(n6410), .A2(n6339), .B1(n6341), .B2(n6411), .Y(n5078) );
	o22ai_1 U6313( .A1(n5520), .A2(n6342), .B1(n6343), .B2(n6411), .Y(n5077) );
	o22ai_1 U6314( .A1(n5697), .A2(n6344), .B1(n6345), .B2(n6411), .Y(n5076) );
	o221ai_1 U6315( .A1(n6412), .A2(n6347), .B1(n7586), .B2(n6349), .C1(n6350), .Y(n6411) );
	nand2_1 U6316( .A(n6360), .B(n6243), .Y(n6350) );
	inv_1 U6317( .A(n6384), .Y(n6360) );
	xnor2_1 U6318( .A(n6413), .B(n6407), .Y(n6412) );
	nand2_1 U6319( .A(n6414), .B(n6408), .Y(n6413) );
	xnor2_1 U6320( .A(n6128), .B(n6354), .Y(n6414) );
	o22ai_1 U6321( .A1(n6415), .A2(n6339), .B1(n6416), .B2(n6341), .Y(n5075) );
	nand2_1 U6322( .A(n7228), .B(n5746), .Y(n6341) );
	nand2_1 U6323( .A(n6277), .B(n5746), .Y(n6339) );
	o22ai_1 U6324( .A1(n6416), .A2(n6343), .B1(n5395), .B2(n6342), .Y(n5074) );
	nand2_1 U6325( .A(n6278), .B(n5746), .Y(n6342) );
	inv_1 U6326( .A(n37), .Y(n6343) );
	o22ai_1 U6327( .A1(n5698), .A2(n6344), .B1(n6416), .B2(n6345), .Y(n5073) );
	inv_1 U6328( .A(n36), .Y(n6345) );
	inv_1 U6329( .A(n6417), .Y(n6416) );
	o22ai_1 U6330( .A1(n5821), .A2(n6349), .B1(n6418), .B2(n6347), .Y(n6417) );
	xnor2_1 U6331( .A(n6419), .B(n6128), .Y(n6418) );
	nand2_1 U6332( .A(n6384), .B(n6347), .Y(n6349) );
	o221ai_1 U6333( .A1(n6419), .A2(n6420), .B1(n6245), .B2(n6421), .C1(n6422), .Y(n6347) );
	a21oi_1 U6334( .A1(n6423), .A2(n6178), .B1(n6424), .Y(n6422) );
	inv_1 U6335( .A(n6195), .Y(n6424) );
	a21oi_1 U6336( .A1(n6113), .A2(n6425), .B1(n6219), .Y(n6423) );
	a221oi_1 U6337( .A1(n6174), .A2(g7264), .B1(n6171), .B2(n7780), .C1(n6426), .Y(n6219) );
	nor2_1 U6338( .A(n6281), .B(n7726), .Y(n6426) );
	inv_1 U6339( .A(n7327), .Y(n6171) );
	inv_1 U6340( .A(n7328), .Y(n6174) );
	nand3_1 U6341( .A(n6185), .B(n6187), .C(n6211), .Y(n6425) );
	o21ai_0 U6342( .A1(n6224), .A2(n6239), .B1(n6204), .Y(n6185) );
	o221ai_1 U6343( .A1(n6427), .A2(n6428), .B1(n6429), .B2(n6430), .C1(n6431), .Y(n6239) );
	o221ai_1 U6344( .A1(n6238), .A2(n6432), .B1(n6236), .B2(n6232), .C1(n6237), .Y(n6431) );
	o22ai_1 U6345( .A1(n6237), .A2(n6236), .B1(n6432), .B2(n6232), .Y(n6430) );
	o22ai_1 U6346( .A1(n6238), .A2(n6236), .B1(n6237), .B2(n6432), .Y(n6428) );
	inv_1 U6347( .A(n6227), .Y(n6432) );
	xor2_1 U6348( .A(n7235), .B(n6127), .X(n6227) );
	xnor2_1 U6349( .A(n7586), .B(n6139), .Y(n6237) );
	xnor2_1 U6350( .A(n7267), .B(n6129), .Y(n6236) );
	inv_1 U6351( .A(n6429), .Y(n6238) );
	xor2_1 U6352( .A(n6146), .B(n5832), .X(n6429) );
	inv_1 U6353( .A(n6232), .Y(n6427) );
	xor2_1 U6354( .A(n6310), .B(n6133), .X(n6232) );
	o221ai_1 U6355( .A1(n6433), .A2(n6434), .B1(n6435), .B2(n6436), .C1(n6437), .Y(n6224) );
	o221ai_1 U6356( .A1(n6233), .A2(n6231), .B1(n6438), .B2(n6234), .C1(n6235), .Y(n6437) );
	o22ai_1 U6357( .A1(n6233), .A2(n6235), .B1(n6438), .B2(n6231), .Y(n6436) );
	o22ai_1 U6358( .A1(n6234), .A2(n6233), .B1(n6438), .B2(n6235), .Y(n6434) );
	xnor2_1 U6359( .A(n5821), .B(n6439), .Y(n6235) );
	inv_1 U6360( .A(n6226), .Y(n6438) );
	xnor2_1 U6361( .A(n7250), .B(n6400), .Y(n6226) );
	xor2_1 U6362( .A(n7232), .B(n6144), .X(n6233) );
	inv_1 U6363( .A(n6435), .Y(n6234) );
	xor2_1 U6364( .A(n6145), .B(n5830), .X(n6435) );
	inv_1 U6365( .A(n6231), .Y(n6433) );
	xnor2_1 U6366( .A(n6311), .B(n6363), .Y(n6231) );
	inv_1 U6367( .A(n6182), .Y(n6113) );
	nor3_1 U6368( .A(n6245), .B(n6184), .C(n6203), .Y(n6182) );
	inv_1 U6369( .A(n6198), .Y(n6184) );
	inv_1 U6370( .A(n6206), .Y(n6421) );
	nor2_1 U6371( .A(n6440), .B(n6441), .Y(n6206) );
	inv_1 U6372( .A(n7720), .Y(n6441) );
	a21oi_1 U6373( .A1(n6122), .A2(n6354), .B1(n6442), .Y(n6420) );
	o211ai_1 U6374( .A1(n6442), .A2(n6122), .B1(n6195), .C1(n6408), .Y(n6384) );
	inv_1 U6375( .A(n6419), .Y(n6408) );
	nor2_1 U6376( .A(n6243), .B(n6121), .Y(n6419) );
	nand2_1 U6377( .A(n6178), .B(n6167), .Y(n6195) );
	o221ai_1 U6378( .A1(n7381), .A2(n6264), .B1(n7382), .B2(n6265), .C1(n6443), .Y(n6167) );
	nand2_1 U6379( .A(g5555), .B(n6163), .Y(n6443) );
	inv_1 U6380( .A(n7737), .Y(n6163) );
	inv_1 U6381( .A(n6166), .Y(n6178) );
	nand2_1 U6382( .A(n6444), .B(n6445), .Y(n6166) );
	nor4_1 U6383( .A(n6446), .B(n6447), .C(n6448), .D(n6449), .Y(n6445) );
	xnor2_1 U6384( .A(n6450), .B(n6348), .Y(n6449) );
	a222oi_1 U6385( .A1(g7084), .A2(n6451), .B1(n7228), .B2(n5427), .C1(g6837), .C2(n6452), .Y(n6450) );
	xnor2_1 U6386( .A(n6453), .B(n6358), .Y(n6448) );
	a222oi_1 U6387( .A1(g7084), .A2(n6454), .B1(n7228), .B2(n5428), .C1(g6837), .C2(n6455), .Y(n6453) );
	mux2i_1 U6388( .A0(n6456), .A1(n6457), .S(n5832), .Y(n6447) );
	nand2_1 U6389( .A(n10063), .B(n6457), .Y(n6456) );
	nand3_1 U6390( .A(n6458), .B(n6459), .C(n6204), .Y(n6446) );
	inv_1 U6391( .A(n6214), .Y(n6204) );
	nand2_1 U6392( .A(n7720), .B(n6440), .Y(n6214) );
	o21ai_0 U6393( .A1(n10064), .A2(n6277), .B1(n6460), .Y(n6440) );
	a22oi_1 U6394( .A1(g6837), .A2(n6461), .B1(g7084), .B2(n6462), .Y(n6460) );
	xnor2_1 U6395( .A(n5821), .B(n6463), .Y(n6459) );
	a222oi_1 U6396( .A1(g7084), .A2(n6464), .B1(n7228), .B2(n5438), .C1(g6837), .C2(n6465), .Y(n6463) );
	xnor2_1 U6397( .A(n5824), .B(n6466), .Y(n6458) );
	a222oi_1 U6398( .A1(g7084), .A2(n6467), .B1(n7228), .B2(n5437), .C1(g6837), .C2(n6468), .Y(n6466) );
	nor4_1 U6399( .A(n6469), .B(n6470), .C(n6471), .D(n6472), .Y(n6444) );
	mux2i_1 U6400( .A0(n6473), .A1(n6474), .S(n5828), .Y(n6472) );
	nand2_1 U6401( .A(n7287), .B(n6474), .Y(n6473) );
	mux2i_1 U6402( .A0(n6475), .A1(n6476), .S(n5834), .Y(n6471) );
	nand2_1 U6403( .A(n7284), .B(n6476), .Y(n6475) );
	mux2i_1 U6404( .A0(n6477), .A1(n6478), .S(n5836), .Y(n6470) );
	nand2_1 U6405( .A(n7609), .B(n6478), .Y(n6477) );
	nand3_1 U6406( .A(n6479), .B(n6480), .C(n6481), .Y(n6469) );
	mux2i_1 U6407( .A0(n6482), .A1(n6483), .S(n5826), .Y(n6481) );
	nor2_1 U6408( .A(n6483), .B(n5359), .Y(n6482) );
	mux2i_1 U6409( .A0(n6484), .A1(n6485), .S(n6277), .Y(n6480) );
	nand2_1 U6410( .A(n6486), .B(n6487), .Y(n6485) );
	a222oi_1 U6411( .A1(n6478), .A2(n7267), .B1(n6457), .B2(n7261), .C1(n6474), .C2(n7235), .Y(n6487) );
	a22oi_1 U6412( .A1(n5487), .A2(g7084), .B1(n5318), .B2(g6837), .Y(n6474) );
	a22oi_1 U6413( .A1(n5486), .A2(g7084), .B1(n5317), .B2(g6837), .Y(n6457) );
	a22oi_1 U6414( .A1(n5484), .A2(g7084), .B1(n5315), .B2(g6837), .Y(n6478) );
	a222oi_1 U6415( .A1(n6488), .A2(n7250), .B1(n6476), .B2(n7232), .C1(n6489), .C2(n7273), .Y(n6486) );
	inv_1 U6416( .A(n6490), .Y(n6489) );
	a22oi_1 U6417( .A1(n5485), .A2(g7084), .B1(n5316), .B2(g6837), .Y(n6476) );
	inv_1 U6418( .A(n6483), .Y(n6488) );
	o22ai_1 U6419( .A1(n9909), .A2(n6278), .B1(n9910), .B2(n6279), .Y(n6483) );
	nand2_1 U6420( .A(n6491), .B(n6492), .Y(n6484) );
	a222oi_1 U6421( .A1(n5826), .A2(n5359), .B1(n5834), .B2(n6493), .C1(n5828), .C2(n6494), .Y(n6492) );
	a222oi_1 U6422( .A1(n5830), .A2(n5305), .B1(n5832), .B2(n5379), .C1(n5836), .C2(n6495), .Y(n6491) );
	mux2i_1 U6423( .A0(n6496), .A1(n6490), .S(n5830), .Y(n6479) );
	nor2_1 U6424( .A(n6490), .B(n5305), .Y(n6496) );
	o22ai_1 U6425( .A1(n9907), .A2(n6278), .B1(n9908), .B2(n6279), .Y(n6490) );
	and4_1 U6426( .A(n6133), .B(n6497), .C(n6127), .D(n6498), .X(n6122) );
	nor3_1 U6427( .A(n6407), .B(n6363), .C(n6400), .Y(n6498) );
	and3_1 U6428( .A(n6392), .B(n6497), .C(n6499), .X(n6442) );
	nor3_1 U6429( .A(n6133), .B(n6139), .C(n6138), .Y(n6499) );
	inv_1 U6430( .A(n6363), .Y(n6138) );
	o221ai_1 U6431( .A1(n6278), .A2(n5519), .B1(n6277), .B2(n6356), .C1(n6500), .Y(n6363) );
	nand2_1 U6432( .A(n9903), .B(g6837), .Y(n6500) );
	inv_1 U6433( .A(n7676), .Y(n6356) );
	inv_1 U6434( .A(n6407), .Y(n6139) );
	o221ai_1 U6435( .A1(n6278), .A2(n5520), .B1(n6277), .B2(n6410), .C1(n6501), .Y(n6407) );
	nand2_1 U6436( .A(n9905), .B(g6837), .Y(n6501) );
	inv_1 U6437( .A(n7671), .Y(n6410) );
	a21oi_1 U6438( .A1(n7228), .A2(n7673), .B1(n6502), .Y(n6133) );
	o22ai_1 U6439( .A1(n5547), .A2(n6279), .B1(n5331), .B2(n6278), .Y(n6502) );
	nor4_1 U6440( .A(n6145), .B(n6144), .C(n6503), .D(n6146), .Y(n6497) );
	o21ai_0 U6441( .A1(n6277), .A2(n6381), .B1(n6504), .Y(n6146) );
	a22oi_1 U6442( .A1(n9899), .A2(g6837), .B1(n9898), .B2(g7084), .Y(n6504) );
	inv_1 U6443( .A(n7668), .Y(n6381) );
	nand2_1 U6444( .A(n6129), .B(n6128), .Y(n6503) );
	inv_1 U6445( .A(n6439), .Y(n6128) );
	o221ai_1 U6446( .A1(n6278), .A2(n5395), .B1(n6277), .B2(n6415), .C1(n6505), .Y(n6439) );
	nand2_1 U6447( .A(n9897), .B(g6837), .Y(n6505) );
	inv_1 U6448( .A(n7670), .Y(n6415) );
	inv_1 U6449( .A(n6368), .Y(n6129) );
	o221ai_1 U6450( .A1(n6278), .A2(n5521), .B1(n6277), .B2(n6369), .C1(n6506), .Y(n6368) );
	nand2_1 U6451( .A(n9896), .B(g6837), .Y(n6506) );
	inv_1 U6452( .A(n7674), .Y(n6369) );
	o221ai_1 U6453( .A1(n6278), .A2(n5522), .B1(n6277), .B2(n6375), .C1(n6507), .Y(n6144) );
	nand2_1 U6454( .A(n9900), .B(g6837), .Y(n6507) );
	inv_1 U6455( .A(n7669), .Y(n6375) );
	o21ai_0 U6456( .A1(n6277), .A2(n6388), .B1(n6508), .Y(n6145) );
	a22oi_1 U6457( .A1(n9902), .A2(g6837), .B1(n9901), .B2(g7084), .Y(n6508) );
	inv_1 U6458( .A(n7672), .Y(n6388) );
	nor3_1 U6459( .A(n6127), .B(n6140), .C(n6354), .Y(n6392) );
	inv_1 U6460( .A(n6243), .Y(n6354) );
	nor3_1 U6461( .A(n6187), .B(n6211), .C(n6198), .Y(n6243) );
	inv_1 U6462( .A(n6203), .Y(n6211) );
	inv_1 U6463( .A(n6400), .Y(n6140) );
	o221ai_1 U6464( .A1(n6278), .A2(n5523), .B1(n6277), .B2(n6402), .C1(n6509), .Y(n6400) );
	nand2_1 U6465( .A(n9904), .B(g6837), .Y(n6509) );
	inv_1 U6466( .A(n7675), .Y(n6402) );
	a221oi_1 U6467( .A1(g7084), .A2(n9895), .B1(n7228), .B2(n7667), .C1(n6510), .Y(n6127) );
	nor2_1 U6468( .A(n5542), .B(n6279), .Y(n6510) );
	nand2_1 U6469( .A(n6279), .B(n5746), .Y(n6344) );
	o22ai_1 U6470( .A1(n6511), .A2(n5601), .B1(n6512), .B2(n6513), .Y(n5072) );
	o22ai_1 U6471( .A1(n6514), .A2(n6515), .B1(n6513), .B2(n6516), .Y(n5071) );
	inv_1 U6472( .A(n7383), .Y(n6515) );
	o22ai_1 U6473( .A1(n6517), .A2(n6518), .B1(n6513), .B2(n6519), .Y(n5070) );
	nand2_1 U6474( .A(n6276), .B(n5746), .Y(n6513) );
	nand2_1 U6475( .A(n6520), .B(n6521), .Y(n6276) );
	nor4_1 U6476( .A(n5821), .B(n5824), .C(n5826), .D(n5828), .Y(n6521) );
	inv_1 U6477( .A(n7235), .Y(n5828) );
	inv_1 U6478( .A(n7250), .Y(n5826) );
	inv_1 U6479( .A(n7586), .Y(n5824) );
	inv_1 U6480( .A(n7242), .Y(n5821) );
	nor4_1 U6481( .A(n5830), .B(n5832), .C(n5834), .D(n5836), .Y(n6520) );
	inv_1 U6482( .A(n7267), .Y(n5836) );
	inv_1 U6483( .A(n7232), .Y(n5834) );
	inv_1 U6484( .A(n7273), .Y(n5830) );
	inv_1 U6485( .A(n7384), .Y(n6518) );
	o22ai_1 U6486( .A1(n6512), .A2(n6522), .B1(n6511), .B2(n6523), .Y(n5069) );
	inv_1 U6487( .A(n7414), .Y(n6523) );
	o22ai_1 U6488( .A1(n6516), .A2(n6522), .B1(n6514), .B2(n5410), .Y(n5068) );
	o22ai_1 U6489( .A1(n6519), .A2(n6522), .B1(n6517), .B2(n6524), .Y(n5067) );
	o22ai_1 U6490( .A1(n6512), .A2(n6525), .B1(n6511), .B2(n6526), .Y(n5066) );
	inv_1 U6491( .A(n7406), .Y(n6526) );
	o22ai_1 U6492( .A1(n6516), .A2(n6525), .B1(n6514), .B2(n6527), .Y(n5065) );
	o22ai_1 U6493( .A1(n6519), .A2(n6525), .B1(n6517), .B2(n5398), .Y(n5064) );
	o22ai_1 U6494( .A1(n6512), .A2(n6528), .B1(n6511), .B2(n5675), .Y(n5063) );
	nand2_1 U6495( .A(n6512), .B(n5746), .Y(n6511) );
	nand2_1 U6496( .A(n6529), .B(n7228), .Y(n6512) );
	o22ai_1 U6497( .A1(n6516), .A2(n6528), .B1(n6514), .B2(n6462), .Y(n5062) );
	inv_1 U6498( .A(n7388), .Y(n6462) );
	nand2_1 U6499( .A(n6516), .B(n5746), .Y(n6514) );
	nand2_1 U6500( .A(n6529), .B(g7084), .Y(n6516) );
	o22ai_1 U6501( .A1(n6519), .A2(n6528), .B1(n6517), .B2(n6461), .Y(n5061) );
	inv_1 U6502( .A(n7391), .Y(n6461) );
	nand2_1 U6503( .A(n6519), .B(n5746), .Y(n6517) );
	nand4_1 U6504( .A(n45), .B(n7267), .C(n7273), .D(n5832), .Y(n6528) );
	inv_1 U6505( .A(n7261), .Y(n5832) );
	nand2_1 U6506( .A(n6529), .B(g6837), .Y(n6519) );
	o22ai_1 U6507( .A1(n6530), .A2(n5427), .B1(n6336), .B2(n6531), .Y(n5060) );
	o22ai_1 U6508( .A1(n6532), .A2(n6451), .B1(n6531), .B2(n6533), .Y(n5059) );
	inv_1 U6509( .A(n7400), .Y(n6451) );
	o22ai_1 U6510( .A1(n6534), .A2(n6452), .B1(n6531), .B2(n6535), .Y(n5058) );
	nand2_1 U6511( .A(n6310), .B(n5745), .Y(n6531) );
	inv_1 U6512( .A(n6348), .Y(n6310) );
	o21ai_0 U6513( .A1(n7406), .A2(n6277), .B1(n6536), .Y(n6348) );
	a22oi_1 U6514( .A1(g6837), .A2(n5398), .B1(g7084), .B2(n6527), .Y(n6536) );
	inv_1 U6515( .A(n7405), .Y(n6527) );
	inv_1 U6516( .A(n7404), .Y(n6452) );
	o22ai_1 U6517( .A1(n6530), .A2(n5428), .B1(n6336), .B2(n6537), .Y(n5057) );
	o22ai_1 U6518( .A1(n6532), .A2(n6454), .B1(n6533), .B2(n6537), .Y(n5056) );
	inv_1 U6519( .A(n7407), .Y(n6454) );
	o22ai_1 U6520( .A1(n6534), .A2(n6455), .B1(n6535), .B2(n6537), .Y(n5055) );
	nand2_1 U6521( .A(n6311), .B(n5745), .Y(n6537) );
	inv_1 U6522( .A(n6358), .Y(n6311) );
	o21ai_0 U6523( .A1(n7414), .A2(n6277), .B1(n6538), .Y(n6358) );
	a22oi_1 U6524( .A1(g6837), .A2(n6524), .B1(g7084), .B2(n5410), .Y(n6538) );
	inv_1 U6525( .A(n7415), .Y(n6524) );
	inv_1 U6526( .A(n7228), .Y(n6277) );
	inv_1 U6527( .A(n7413), .Y(n6455) );
	o22ai_1 U6528( .A1(n6336), .A2(n6539), .B1(n6495), .B2(n6530), .Y(n5054) );
	inv_1 U6529( .A(n7609), .Y(n6495) );
	o22ai_1 U6530( .A1(n6533), .A2(n6539), .B1(n6532), .B2(n5484), .Y(n5053) );
	o22ai_1 U6531( .A1(n6535), .A2(n6539), .B1(n6534), .B2(n5315), .Y(n5052) );
	inv_1 U6532( .A(n46), .Y(n6539) );
	o22ai_1 U6533( .A1(n6336), .A2(n6540), .B1(n6493), .B2(n6530), .Y(n5051) );
	inv_1 U6534( .A(n7284), .Y(n6493) );
	o22ai_1 U6535( .A1(n6540), .A2(n6533), .B1(n6532), .B2(n5485), .Y(n5050) );
	o22ai_1 U6536( .A1(n6540), .A2(n6535), .B1(n6534), .B2(n5316), .Y(n5049) );
	inv_1 U6537( .A(n45), .Y(n6540) );
	o22ai_1 U6538( .A1(n6336), .A2(n6541), .B1(n5379), .B2(n6530), .Y(n5048) );
	o22ai_1 U6539( .A1(n6533), .A2(n6541), .B1(n6532), .B2(n5486), .Y(n5047) );
	o22ai_1 U6540( .A1(n6535), .A2(n6541), .B1(n6534), .B2(n5317), .Y(n5046) );
	inv_1 U6541( .A(n43), .Y(n6541) );
	o22ai_1 U6542( .A1(n6336), .A2(n6542), .B1(n5305), .B2(n6530), .Y(n5045) );
	o22ai_1 U6543( .A1(n6533), .A2(n6542), .B1(n6532), .B2(n5646), .Y(n5044) );
	o22ai_1 U6544( .A1(n6535), .A2(n6542), .B1(n6534), .B2(n5635), .Y(n5043) );
	inv_1 U6545( .A(n42), .Y(n6542) );
	o22ai_1 U6546( .A1(n6336), .A2(n6543), .B1(n6494), .B2(n6530), .Y(n5042) );
	inv_1 U6547( .A(n7287), .Y(n6494) );
	o22ai_1 U6548( .A1(n6533), .A2(n6543), .B1(n6532), .B2(n5487), .Y(n5041) );
	o22ai_1 U6549( .A1(n6535), .A2(n6543), .B1(n6534), .B2(n5318), .Y(n5040) );
	inv_1 U6550( .A(n41), .Y(n6543) );
	o22ai_1 U6551( .A1(n6336), .A2(n6544), .B1(n5359), .B2(n6530), .Y(n5039) );
	o22ai_1 U6552( .A1(n6533), .A2(n6544), .B1(n6532), .B2(n5647), .Y(n5038) );
	o22ai_1 U6553( .A1(n6535), .A2(n6544), .B1(n6534), .B2(n5636), .Y(n5037) );
	inv_1 U6554( .A(n40), .Y(n6544) );
	o22ai_1 U6555( .A1(n6336), .A2(n6525), .B1(n6530), .B2(n5437), .Y(n5036) );
	o22ai_1 U6556( .A1(n6525), .A2(n6533), .B1(n6532), .B2(n6467), .Y(n5035) );
	inv_1 U6557( .A(n7399), .Y(n6467) );
	o22ai_1 U6558( .A1(n6525), .A2(n6535), .B1(n6534), .B2(n6468), .Y(n5034) );
	inv_1 U6559( .A(n7401), .Y(n6468) );
	inv_1 U6560( .A(n39), .Y(n6525) );
	o22ai_1 U6561( .A1(n6336), .A2(n6522), .B1(n6530), .B2(n5438), .Y(n5033) );
	nand2_1 U6562( .A(n5756), .B(n6336), .Y(n6530) );
	nand2_1 U6563( .A(n7720), .B(n7228), .Y(n6336) );
	o22ai_1 U6564( .A1(n6522), .A2(n6533), .B1(n6532), .B2(n6464), .Y(n5032) );
	inv_1 U6565( .A(n7402), .Y(n6464) );
	nand2_1 U6566( .A(n5756), .B(n6533), .Y(n6532) );
	nand2_1 U6567( .A(n7720), .B(g7084), .Y(n6533) );
	o22ai_1 U6568( .A1(n6522), .A2(n6535), .B1(n6534), .B2(n6465), .Y(n5031) );
	inv_1 U6569( .A(n7408), .Y(n6465) );
	nand2_1 U6570( .A(n5756), .B(n6535), .Y(n6534) );
	nand2_1 U6571( .A(n7720), .B(g6837), .Y(n6535) );
	inv_1 U6572( .A(n38), .Y(n6522) );
	a21oi_1 U6573( .A1(n6545), .A2(n6546), .B1(n6547), .Y(n5030) );
	a21oi_1 U6574( .A1(n5337), .A2(n6548), .B1(n6549), .Y(n5029) );
	a21oi_1 U6575( .A1(n5546), .A2(n6550), .B1(n6551), .Y(n5028) );
	o22ai_1 U6576( .A1(n6552), .A2(n6553), .B1(n6554), .B2(n6555), .Y(n5027) );
	inv_1 U6577( .A(n7499), .Y(n6553) );
	o22ai_1 U6578( .A1(n6556), .A2(n6557), .B1(n6554), .B2(n6558), .Y(n5026) );
	inv_1 U6579( .A(n7522), .Y(n6557) );
	o22ai_1 U6580( .A1(n6559), .A2(n6560), .B1(n6554), .B2(n6561), .Y(n5025) );
	nand4_1 U6581( .A(n6562), .B(n6563), .C(n6564), .D(n6565), .Y(n6554) );
	a222oi_1 U6582( .A1(g7357), .A2(n6566), .B1(n7237), .B2(n6567), .C1(g7229), .C2(n5391), .Y(n6565) );
	nand2_1 U6583( .A(n9911), .B(n10067), .Y(n6567) );
	nand4_1 U6584( .A(n6568), .B(n6569), .C(n6570), .D(n6571), .Y(n6564) );
	nor3_1 U6585( .A(n6572), .B(n6573), .C(n6574), .Y(n6571) );
	xor2_1 U6586( .A(n6575), .B(n10070), .X(n6574) );
	xor2_1 U6587( .A(n6576), .B(n7690), .X(n6573) );
	nand3_1 U6588( .A(n6577), .B(n6578), .C(n6579), .Y(n6572) );
	xor2_1 U6589( .A(n9952), .B(n6580), .X(n6579) );
	xnor2_1 U6590( .A(n10071), .B(n6581), .Y(n6578) );
	xnor2_1 U6591( .A(n10072), .B(n6582), .Y(n6577) );
	nor3_1 U6592( .A(n6583), .B(n6584), .C(n6585), .Y(n6570) );
	xor2_1 U6593( .A(n6586), .B(n9962), .X(n6585) );
	xor2_1 U6594( .A(n6587), .B(n10068), .X(n6584) );
	xor2_1 U6595( .A(n6588), .B(n7296), .X(n6583) );
	xnor2_1 U6596( .A(n7300), .B(n6589), .Y(n6569) );
	xnor2_1 U6597( .A(n7692), .B(n6590), .Y(n6568) );
	o22ai_1 U6598( .A1(n6547), .A2(n5571), .B1(n6591), .B2(n6592), .Y(n5024) );
	o22ai_1 U6599( .A1(n6549), .A2(n6593), .B1(n6591), .B2(n6594), .Y(n5023) );
	o22ai_1 U6600( .A1(n6551), .A2(n5478), .B1(n6591), .B2(n5809), .Y(n5022) );
	nand2_1 U6601( .A(n6595), .B(n9963), .Y(n6591) );
	o22ai_1 U6602( .A1(n6547), .A2(n5613), .B1(n6592), .B2(n6596), .Y(n5021) );
	o21ai_0 U6603( .A1(n5362), .A2(n6597), .B1(n5762), .Y(n6547) );
	o22ai_1 U6604( .A1(n6549), .A2(n6566), .B1(n6594), .B2(n6596), .Y(n5020) );
	inv_1 U6605( .A(n5298), .Y(n6594) );
	nor2_1 U6606( .A(n6598), .B(RST), .Y(n5298) );
	inv_1 U6607( .A(n7448), .Y(n6566) );
	o22ai_1 U6608( .A1(n6551), .A2(n5391), .B1(n5809), .B2(n6596), .Y(n5019) );
	nand2_1 U6609( .A(n6599), .B(n9963), .Y(n6596) );
	nand2_1 U6610( .A(g7229), .B(n5744), .Y(n5809) );
	o21ai_0 U6611( .A1(n5362), .A2(n6600), .B1(n5740), .Y(n6551) );
	o22ai_1 U6612( .A1(n6552), .A2(n6601), .B1(n10071), .B2(n6555), .Y(n5018) );
	inv_1 U6613( .A(n7501), .Y(n6601) );
	o22ai_1 U6614( .A1(n6556), .A2(n6602), .B1(n10071), .B2(n6558), .Y(n5017) );
	inv_1 U6615( .A(n7500), .Y(n6602) );
	o22ai_1 U6616( .A1(n6559), .A2(n5473), .B1(n10071), .B2(n6561), .Y(n5016) );
	o22ai_1 U6617( .A1(n6552), .A2(n6603), .B1(n10072), .B2(n6555), .Y(n5015) );
	inv_1 U6618( .A(n7503), .Y(n6603) );
	o22ai_1 U6619( .A1(n6556), .A2(n6604), .B1(n10072), .B2(n6558), .Y(n5014) );
	inv_1 U6620( .A(n7502), .Y(n6604) );
	o22ai_1 U6621( .A1(n6559), .A2(n5476), .B1(n10072), .B2(n6561), .Y(n5013) );
	o22ai_1 U6622( .A1(n6552), .A2(n6605), .B1(n7692), .B2(n6555), .Y(n5012) );
	inv_1 U6623( .A(n7512), .Y(n6605) );
	o22ai_1 U6624( .A1(n6556), .A2(n6606), .B1(n7692), .B2(n6558), .Y(n5011) );
	inv_1 U6625( .A(n7511), .Y(n6606) );
	o22ai_1 U6626( .A1(n6559), .A2(n5482), .B1(n7692), .B2(n6561), .Y(n5010) );
	o22ai_1 U6627( .A1(n6552), .A2(n6607), .B1(n10068), .B2(n6555), .Y(n5009) );
	inv_1 U6628( .A(n7514), .Y(n6607) );
	o22ai_1 U6629( .A1(n6556), .A2(n6608), .B1(n10068), .B2(n6558), .Y(n5008) );
	inv_1 U6630( .A(n7513), .Y(n6608) );
	o22ai_1 U6631( .A1(n6559), .A2(n5479), .B1(n10068), .B2(n6561), .Y(n5007) );
	o22ai_1 U6632( .A1(n6552), .A2(n6609), .B1(n7296), .B2(n6555), .Y(n5006) );
	inv_1 U6633( .A(n7516), .Y(n6609) );
	o22ai_1 U6634( .A1(n6556), .A2(n6610), .B1(n7296), .B2(n6558), .Y(n5005) );
	inv_1 U6635( .A(n7515), .Y(n6610) );
	o22ai_1 U6636( .A1(n6559), .A2(n5480), .B1(n7296), .B2(n6561), .Y(n5004) );
	o22ai_1 U6637( .A1(n6552), .A2(n6611), .B1(n10070), .B2(n6555), .Y(n5003) );
	inv_1 U6638( .A(n7518), .Y(n6611) );
	o22ai_1 U6639( .A1(n6556), .A2(n6612), .B1(n10070), .B2(n6558), .Y(n5002) );
	inv_1 U6640( .A(n7517), .Y(n6612) );
	o22ai_1 U6641( .A1(n6559), .A2(n5477), .B1(n10070), .B2(n6561), .Y(n5001) );
	o22ai_1 U6642( .A1(n6552), .A2(n6613), .B1(n7300), .B2(n6555), .Y(n5000) );
	inv_1 U6643( .A(n7509), .Y(n6613) );
	inv_1 U6644( .A(n6614), .Y(n50) );
	o22ai_1 U6645( .A1(n6556), .A2(n6615), .B1(n7300), .B2(n6558), .Y(n4999) );
	inv_1 U6646( .A(n7508), .Y(n6615) );
	o22ai_1 U6647( .A1(n6559), .A2(n5475), .B1(n7300), .B2(n6561), .Y(n4998) );
	o22ai_1 U6648( .A1(n6552), .A2(n6616), .B1(n9952), .B2(n6555), .Y(n4997) );
	o22ai_1 U6649( .A1(n6556), .A2(n6617), .B1(n9952), .B2(n6558), .Y(n4996) );
	o22ai_1 U6650( .A1(n6559), .A2(n5614), .B1(n9952), .B2(n6561), .Y(n4995) );
	o22ai_1 U6651( .A1(n6552), .A2(n6618), .B1(n7690), .B2(n6555), .Y(n4994) );
	inv_1 U6652( .A(n7507), .Y(n6618) );
	o22ai_1 U6653( .A1(n6556), .A2(n6619), .B1(n7690), .B2(n6558), .Y(n4993) );
	inv_1 U6654( .A(n7506), .Y(n6619) );
	o22ai_1 U6655( .A1(n6559), .A2(n5474), .B1(n7690), .B2(n6561), .Y(n4992) );
	o22ai_1 U6656( .A1(n6552), .A2(n6620), .B1(n9962), .B2(n6555), .Y(n4991) );
	or2_0 U6657( .A(n6546), .B(RST), .X(n6555) );
	inv_1 U6658( .A(n7520), .Y(n6620) );
	nand2_1 U6659( .A(n5756), .B(n6546), .Y(n6552) );
	nand3_1 U6660( .A(n9964), .B(n6621), .C(n9914), .Y(n6546) );
	o22ai_1 U6661( .A1(n6556), .A2(n6622), .B1(n9962), .B2(n6558), .Y(n4990) );
	or2_0 U6662( .A(n6548), .B(RST), .X(n6558) );
	inv_1 U6663( .A(n7519), .Y(n6622) );
	nand2_1 U6664( .A(n5757), .B(n6548), .Y(n6556) );
	nand2_1 U6665( .A(n6623), .B(g7357), .Y(n6548) );
	o22ai_1 U6666( .A1(n6559), .A2(n5481), .B1(n9962), .B2(n6561), .Y(n4989) );
	or2_0 U6667( .A(n6550), .B(RST), .X(n6561) );
	nand2_1 U6668( .A(n5757), .B(n6550), .Y(n6559) );
	nand2_1 U6669( .A(n6623), .B(g7229), .Y(n6550) );
	and3_1 U6670( .A(n9964), .B(n6624), .C(n9914), .X(n6623) );
	nor2_1 U6671( .A(n6625), .B(n6549), .Y(n4988) );
	xnor2_1 U6672( .A(n6626), .B(n10071), .Y(n6625) );
	a211oi_1 U6673( .A1(n5366), .A2(n6627), .B1(n6549), .C1(n6626), .Y(n4987) );
	nor2_1 U6674( .A(n6627), .B(n5366), .Y(n6626) );
	nor3_1 U6675( .A(n6549), .B(n6628), .C(n6629), .Y(n4986) );
	a21oi_1 U6676( .A1(n6630), .A2(n10068), .B1(n7692), .Y(n6629) );
	inv_1 U6677( .A(n6627), .Y(n6628) );
	nand3_1 U6678( .A(n7692), .B(n10068), .C(n6630), .Y(n6627) );
	nor2_1 U6679( .A(n6631), .B(n6549), .Y(n4985) );
	xnor2_1 U6680( .A(n6630), .B(n10068), .Y(n6631) );
	nor3_1 U6681( .A(n6549), .B(n6630), .C(n6632), .Y(n4984) );
	a21oi_1 U6682( .A1(n6633), .A2(n10070), .B1(n7296), .Y(n6632) );
	and3_1 U6683( .A(n7296), .B(n10070), .C(n6633), .X(n6630) );
	nor2_1 U6684( .A(n6634), .B(n6549), .Y(n4983) );
	xnor2_1 U6685( .A(n10070), .B(n6633), .Y(n6634) );
	a211oi_1 U6686( .A1(n6635), .A2(n5808), .B1(n6549), .C1(n6633), .Y(n4982) );
	nor2_1 U6687( .A(n5808), .B(n6635), .Y(n6633) );
	nand2_1 U6688( .A(n9952), .B(n5806), .Y(n5808) );
	inv_1 U6689( .A(n7300), .Y(n6635) );
	nor3_1 U6690( .A(n6549), .B(n5806), .C(n6636), .Y(n4981) );
	a21oi_1 U6691( .A1(n9962), .A2(n6621), .B1(n7690), .Y(n6636) );
	and3_1 U6692( .A(n7690), .B(n6621), .C(n9962), .X(n5806) );
	nor2_1 U6693( .A(n6637), .B(n6549), .Y(n4980) );
	inv_1 U6694( .A(n5807), .Y(n6549) );
	a21oi_1 U6695( .A1(g7357), .A2(n9963), .B1(RST), .Y(n5807) );
	xnor2_1 U6696( .A(n6621), .B(n9962), .Y(n6637) );
	nor2_1 U6697( .A(n6597), .B(n7276), .Y(n6621) );
	o32ai_1 U6698( .A1(n6624), .A2(n7237), .A3(RST), .B1(n5981), .B2(n6592), .Y(n4979) );
	inv_1 U6699( .A(n7276), .Y(n6624) );
	o32ai_1 U6700( .A1(n5362), .A2(n7237), .A3(RST), .B1(n6592), .B2(n6638), .Y(n4978) );
	nand2_1 U6701( .A(n7237), .B(n5744), .Y(n6592) );
	o22ai_1 U6702( .A1(n5983), .A2(n6639), .B1(n5984), .B2(n5674), .Y(n4977) );
	and2_0 U6703( .A(n5749), .B(g16399), .X(n4976) );
	and2_0 U6704( .A(n5752), .B(n6640), .X(n4975) );
	o22ai_1 U6705( .A1(n5563), .A2(n6641), .B1(n6642), .B2(n6643), .Y(n4974) );
	o22ai_1 U6706( .A1(n5722), .A2(n6644), .B1(n6643), .B2(n6645), .Y(n4973) );
	o22ai_1 U6707( .A1(n6646), .A2(n6647), .B1(n6643), .B2(n6648), .Y(n4972) );
	nand3_1 U6708( .A(n7589), .B(n6599), .C(n6649), .Y(n6643) );
	inv_1 U6709( .A(n7637), .Y(n6646) );
	o22ai_1 U6710( .A1(n5559), .A2(n6641), .B1(n6650), .B2(n6642), .Y(n4971) );
	o22ai_1 U6711( .A1(n5349), .A2(n6644), .B1(n6650), .B2(n6645), .Y(n4970) );
	o22ai_1 U6712( .A1(n6650), .A2(n6648), .B1(n6651), .B2(n6647), .Y(n4969) );
	inv_1 U6713( .A(n7661), .Y(n6651) );
	mux2i_1 U6714( .A0(n6652), .A1(n6653), .S(n5999), .Y(n6650) );
	nor2_1 U6715( .A(n6654), .B(n6655), .Y(n6652) );
	mux2_1 U6716( .A0(n6656), .A1(n6657), .S(n6658), .X(n6654) );
	o22ai_1 U6717( .A1(n5554), .A2(n6641), .B1(n6659), .B2(n6642), .Y(n4968) );
	o22ai_1 U6718( .A1(n5344), .A2(n6644), .B1(n6659), .B2(n6645), .Y(n4967) );
	o22ai_1 U6719( .A1(n6659), .A2(n6648), .B1(n6660), .B2(n6647), .Y(n4966) );
	inv_1 U6720( .A(n7660), .Y(n6660) );
	mux2i_1 U6721( .A0(n6661), .A1(n6662), .S(n5999), .Y(n6659) );
	nor2_1 U6722( .A(n6663), .B(n6664), .Y(n6661) );
	inv_1 U6723( .A(n6657), .Y(n6664) );
	a222oi_1 U6724( .A1(n6665), .A2(n6666), .B1(n6667), .B2(n6668), .C1(n6669), .C2(n6670), .Y(n6657) );
	o22ai_1 U6725( .A1(n6665), .A2(n6671), .B1(n6672), .B2(n6673), .Y(n6670) );
	o22ai_1 U6726( .A1(n6674), .A2(n6675), .B1(n6676), .B2(n6665), .Y(n6668) );
	a21oi_1 U6727( .A1(n6677), .A2(n6678), .B1(n6679), .Y(n6676) );
	o22ai_1 U6728( .A1(n6680), .A2(n6681), .B1(n6682), .B2(n6683), .Y(n6677) );
	o32ai_1 U6729( .A1(n6669), .A2(n6684), .A3(n6682), .B1(n6685), .B2(n6667), .Y(n6666) );
	a21oi_1 U6730( .A1(n6686), .A2(n6682), .B1(n6687), .Y(n6685) );
	mux2i_1 U6731( .A0(n6680), .A1(n6688), .S(n6678), .Y(n6687) );
	or2_0 U6732( .A(n6675), .B(n6681), .X(n6688) );
	mux2i_1 U6733( .A0(n6655), .A1(n6658), .S(n6656), .Y(n6663) );
	inv_1 U6734( .A(n6689), .Y(n6658) );
	nand2_1 U6735( .A(n6690), .B(n6691), .Y(n6655) );
	nand3_1 U6736( .A(n6681), .B(n6692), .C(n6693), .Y(n6691) );
	inv_1 U6737( .A(n6674), .Y(n6681) );
	mux2i_1 U6738( .A0(n6694), .A1(n6695), .S(n6665), .Y(n6690) );
	o221ai_1 U6739( .A1(n6696), .A2(n15047), .B1(n5354), .B2(n15046), .C1(n6697), .Y(n6665) );
	nand2_1 U6740( .A(g1730), .B(g5695), .Y(n6697) );
	o221ai_1 U6741( .A1(n6698), .A2(n6671), .B1(n6669), .B2(n6699), .C1(n6700), .Y(n6695) );
	mux2i_1 U6742( .A0(n6701), .A1(n6702), .S(n6667), .Y(n6700) );
	nor2_1 U6743( .A(n6703), .B(n6678), .Y(n6702) );
	a21oi_1 U6744( .A1(n6684), .A2(n6698), .B1(n6692), .Y(n6703) );
	nor2_1 U6745( .A(n6674), .B(n6704), .Y(n6701) );
	a221oi_1 U6746( .A1(n6705), .A2(n6674), .B1(n6706), .B2(n6692), .C1(n6679), .Y(n6699) );
	inv_1 U6747( .A(n6678), .Y(n6669) );
	o21ai_0 U6748( .A1(n6684), .A2(n6707), .B1(n6708), .Y(n6694) );
	mux2i_1 U6749( .A0(n6709), .A1(n6710), .S(n6678), .Y(n6708) );
	o221ai_1 U6750( .A1(n6696), .A2(n15053), .B1(n5354), .B2(n15051), .C1(n6711), .Y(n6678) );
	nand2_1 U6751( .A(g1745), .B(g5695), .Y(n6711) );
	o22ai_1 U6752( .A1(n6698), .A2(n6675), .B1(n6712), .B2(n6673), .Y(n6710) );
	inv_1 U6753( .A(n6706), .Y(n6673) );
	nor2_1 U6754( .A(n6667), .B(n6682), .Y(n6706) );
	nor3_1 U6755( .A(n6705), .B(n6679), .C(n6693), .Y(n6709) );
	nor2_1 U6756( .A(n6698), .B(n6672), .Y(n6679) );
	a21oi_1 U6757( .A1(n6674), .A2(n6667), .B1(n6682), .Y(n6707) );
	inv_1 U6758( .A(n6698), .Y(n6682) );
	o221ai_1 U6759( .A1(n6696), .A2(n15049), .B1(n5354), .B2(n15048), .C1(n6713), .Y(n6698) );
	nand2_1 U6760( .A(g1760), .B(g5695), .Y(n6713) );
	o221ai_1 U6761( .A1(n6696), .A2(n15045), .B1(n5354), .B2(n15044), .C1(n6714), .Y(n6674) );
	nand2_1 U6762( .A(g5695), .B(g1775), .Y(n6714) );
	o22ai_1 U6763( .A1(n6641), .A2(n5615), .B1(n6642), .B2(n6715), .Y(n4965) );
	o22ai_1 U6764( .A1(n6644), .A2(n5595), .B1(n6645), .B2(n6715), .Y(n4964) );
	o22ai_1 U6765( .A1(n6647), .A2(n5404), .B1(n6648), .B2(n6715), .Y(n4963) );
	nand2_1 U6766( .A(n6656), .B(n5999), .Y(n6715) );
	o211ai_1 U6767( .A1(n6716), .A2(n5404), .B1(n6717), .C1(n6718), .Y(n6656) );
	a22oi_1 U6768( .A1(n9918), .A2(g7194), .B1(n9917), .B2(n7225), .Y(n6718) );
	nand3_1 U6769( .A(n7256), .B(n6719), .C(g1922), .Y(n6717) );
	o22ai_1 U6770( .A1(n6641), .A2(n5616), .B1(n6642), .B2(n6720), .Y(n4962) );
	o22ai_1 U6771( .A1(n6644), .A2(n5596), .B1(n6645), .B2(n6720), .Y(n4961) );
	inv_1 U6772( .A(n21), .Y(n6645) );
	nand2_1 U6773( .A(n6721), .B(n5744), .Y(n6644) );
	o22ai_1 U6774( .A1(n6647), .A2(n5405), .B1(n6648), .B2(n6720), .Y(n4960) );
	nand2_1 U6775( .A(n6689), .B(n5999), .Y(n6720) );
	o211ai_1 U6776( .A1(n6716), .A2(n5405), .B1(n6722), .C1(n6723), .Y(n6689) );
	a22oi_1 U6777( .A1(n9920), .A2(g7194), .B1(n9919), .B2(n7225), .Y(n6723) );
	nand3_1 U6778( .A(n7256), .B(n6724), .C(g1904), .Y(n6722) );
	inv_1 U6779( .A(n20), .Y(n6648) );
	nand2_1 U6780( .A(n5757), .B(n6716), .Y(n6647) );
	o22ai_1 U6781( .A1(n6725), .A2(n6726), .B1(n6727), .B2(n6728), .Y(n4959) );
	inv_1 U6782( .A(n7357), .Y(n6728) );
	o22ai_1 U6783( .A1(n6725), .A2(n6729), .B1(n6730), .B2(n6731), .Y(n4958) );
	inv_1 U6784( .A(n7358), .Y(n6731) );
	o22ai_1 U6785( .A1(n6725), .A2(n6732), .B1(n6733), .B2(n5508), .Y(n4957) );
	o21ai_0 U6786( .A1(n6675), .A2(n6734), .B1(n5759), .Y(n6725) );
	nand2_1 U6787( .A(n6672), .B(n6680), .Y(n6675) );
	o22ai_1 U6788( .A1(n6726), .A2(n6735), .B1(n6727), .B2(n6736), .Y(n4956) );
	inv_1 U6789( .A(n7351), .Y(n6736) );
	o22ai_1 U6790( .A1(n6729), .A2(n6735), .B1(n6730), .B2(n6737), .Y(n4955) );
	inv_1 U6791( .A(n7352), .Y(n6737) );
	o22ai_1 U6792( .A1(n6732), .A2(n6735), .B1(n6733), .B2(n5507), .Y(n4954) );
	o221ai_1 U6793( .A1(n6672), .A2(n6738), .B1(n6739), .B2(n6683), .C1(n5749), .Y(n6735) );
	inv_1 U6794( .A(n6686), .Y(n6683) );
	nor2_1 U6795( .A(n6704), .B(n6712), .Y(n6686) );
	mux2i_1 U6796( .A0(n5984), .A1(n5983), .S(n6667), .Y(n6738) );
	o22ai_1 U6797( .A1(n6726), .A2(n6740), .B1(n6727), .B2(n6741), .Y(n4953) );
	inv_1 U6798( .A(n7353), .Y(n6741) );
	o22ai_1 U6799( .A1(n6729), .A2(n6740), .B1(n6730), .B2(n6742), .Y(n4952) );
	inv_1 U6800( .A(n7354), .Y(n6742) );
	o22ai_1 U6801( .A1(n6732), .A2(n6740), .B1(n6733), .B2(n5506), .Y(n4951) );
	o211ai_1 U6802( .A1(n6680), .A2(n6739), .B1(n6671), .C1(n5740), .Y(n6740) );
	inv_1 U6803( .A(n6734), .Y(n6739) );
	xnor2_1 U6804( .A(n6693), .B(n5983), .Y(n6734) );
	inv_1 U6805( .A(n6667), .Y(n6693) );
	o22ai_1 U6806( .A1(n6726), .A2(n6743), .B1(n6727), .B2(n6744), .Y(n4950) );
	inv_1 U6807( .A(n7355), .Y(n6744) );
	nand2_1 U6808( .A(n6726), .B(n5744), .Y(n6727) );
	nand2_1 U6809( .A(n7225), .B(n6640), .Y(n6726) );
	o22ai_1 U6810( .A1(n6729), .A2(n6743), .B1(n6730), .B2(n6745), .Y(n4949) );
	inv_1 U6811( .A(n7356), .Y(n6745) );
	nand2_1 U6812( .A(n6729), .B(n5743), .Y(n6730) );
	nand2_1 U6813( .A(g7194), .B(n6640), .Y(n6729) );
	o22ai_1 U6814( .A1(n6732), .A2(n6743), .B1(n6733), .B2(n5505), .Y(n4948) );
	nand2_1 U6815( .A(n6732), .B(n5743), .Y(n6733) );
	o221ai_1 U6816( .A1(n6098), .A2(n6684), .B1(g3229), .B2(n6671), .C1(n6746), .Y(n6743) );
	a21oi_1 U6817( .A1(n6747), .A2(n6667), .B1(RST), .Y(n6746) );
	o221ai_1 U6818( .A1(n7356), .A2(n6721), .B1(n7355), .B2(n6748), .C1(n6749), .Y(n6667) );
	nand2_1 U6819( .A(g7052), .B(n5505), .Y(n6749) );
	o22ai_1 U6820( .A1(n6680), .A2(n5983), .B1(n6750), .B2(n6704), .Y(n6747) );
	nor2_1 U6821( .A(n6672), .B(n5983), .Y(n6750) );
	inv_1 U6822( .A(n6692), .Y(n6680) );
	inv_1 U6823( .A(n6705), .Y(n6671) );
	nor2_1 U6824( .A(n6692), .B(n6672), .Y(n6705) );
	inv_1 U6825( .A(n6712), .Y(n6672) );
	o221ai_1 U6826( .A1(n7354), .A2(n6721), .B1(n7353), .B2(n6748), .C1(n6751), .Y(n6712) );
	nand2_1 U6827( .A(g7052), .B(n5506), .Y(n6751) );
	o221ai_1 U6828( .A1(n7352), .A2(n6721), .B1(n7351), .B2(n6748), .C1(n6752), .Y(n6692) );
	nand2_1 U6829( .A(g7052), .B(n5507), .Y(n6752) );
	inv_1 U6830( .A(n6704), .Y(n6684) );
	o221ai_1 U6831( .A1(n7358), .A2(n6721), .B1(n7357), .B2(n6748), .C1(n6753), .Y(n6704) );
	nand2_1 U6832( .A(g7052), .B(n5508), .Y(n6753) );
	nand2_1 U6833( .A(g7052), .B(n6640), .Y(n6732) );
	o32ai_1 U6834( .A1(n6754), .A2(n6599), .A3(n6638), .B1(n6755), .B2(n6756), .Y(n6640) );
	nor2_1 U6835( .A(n6649), .B(n6595), .Y(n6756) );
	inv_1 U6836( .A(n6653), .Y(n6595) );
	inv_1 U6837( .A(n6754), .Y(n6649) );
	inv_1 U6838( .A(n6662), .Y(n6599) );
	o21ai_0 U6839( .A1(n6748), .A2(n5563), .B1(n6757), .Y(n6754) );
	a22oi_1 U6840( .A1(n7637), .A2(g7052), .B1(n9921), .B2(g7194), .Y(n6757) );
	and2_0 U6841( .A(g1938), .B(n5754), .X(n4947) );
	inv_1 U6842( .A(n6758), .Y(n4946) );
	and2_0 U6843( .A(g1923), .B(n5758), .X(n4945) );
	o22ai_1 U6844( .A1(n6759), .A2(n6760), .B1(n6761), .B2(n5648), .Y(n4944) );
	o22ai_1 U6845( .A1(n6759), .A2(n6762), .B1(n6763), .B2(n6764), .Y(n4943) );
	inv_1 U6846( .A(n7460), .Y(n6764) );
	o22ai_1 U6847( .A1(n6759), .A2(n6765), .B1(n6766), .B2(n5419), .Y(n4942) );
	o22ai_1 U6848( .A1(n6760), .A2(n6767), .B1(n6761), .B2(n5649), .Y(n4941) );
	o22ai_1 U6849( .A1(n6762), .A2(n6767), .B1(n6763), .B2(n6768), .Y(n4940) );
	inv_1 U6850( .A(n7455), .Y(n6768) );
	o22ai_1 U6851( .A1(n6765), .A2(n6767), .B1(n6766), .B2(n5420), .Y(n4939) );
	o22ai_1 U6852( .A1(n6769), .A2(n6760), .B1(n6761), .B2(n5650), .Y(n4938) );
	or2_0 U6853( .A(RST), .B(n7257), .X(n6761) );
	o22ai_1 U6854( .A1(n6769), .A2(n6762), .B1(n6763), .B2(n6770), .Y(n4937) );
	inv_1 U6855( .A(n7452), .Y(n6770) );
	or2_0 U6856( .A(RST), .B(g8082), .X(n6763) );
	o22ai_1 U6857( .A1(n6769), .A2(n6765), .B1(n6766), .B2(n5418), .Y(n4936) );
	or2_0 U6858( .A(RST), .B(g8012), .X(n6766) );
	and2_0 U6859( .A(g1948), .B(n5753), .X(n4935) );
	and2_0 U6860( .A(g1954), .B(n5748), .X(n4934) );
	and2_0 U6861( .A(g1952), .B(n5758), .X(n4933) );
	and2_0 U6862( .A(g1944), .B(n5747), .X(n4932) );
	o22ai_1 U6863( .A1(n6638), .A2(n6641), .B1(n6642), .B2(n6771), .Y(n4931) );
	o22ai_1 U6864( .A1(n6641), .A2(n6771), .B1(n9965), .B2(n6642), .Y(n4930) );
	o22ai_1 U6865( .A1(n6641), .A2(n5590), .B1(n6118), .B2(n6642), .Y(n4929) );
	nand2_1 U6866( .A(n7225), .B(n5743), .Y(n6642) );
	nand2_1 U6867( .A(n6748), .B(n5743), .Y(n6641) );
	nor2_1 U6868( .A(RST), .B(n6696), .Y(n4928) );
	inv_1 U6869( .A(g5738), .Y(n6696) );
	and2_0 U6870( .A(g1778), .B(n5758), .X(n4927) );
	and2_0 U6871( .A(g1776), .B(n5759), .X(n4926) );
	and2_0 U6872( .A(g1763), .B(n5759), .X(n4925) );
	and2_0 U6873( .A(g1761), .B(n5759), .X(n4924) );
	and2_0 U6874( .A(g1748), .B(n5759), .X(n4923) );
	and2_0 U6875( .A(g1746), .B(n5746), .X(n4922) );
	and2_0 U6876( .A(g1733), .B(n5759), .X(n4921) );
	and2_0 U6877( .A(g1731), .B(n5759), .X(n4920) );
	and2_0 U6878( .A(n5760), .B(n6150), .X(n4919) );
	mux2i_1 U6879( .A0(g1679), .A1(n6772), .S(n7731), .Y(n6150) );
	mux2i_1 U6880( .A0(n6773), .A1(n9966), .S(n6774), .Y(n6772) );
	nor2_1 U6881( .A(RST), .B(n6775), .Y(n4918) );
	and2_0 U6882( .A(g1671), .B(n5742), .X(n4917) );
	o22ai_1 U6883( .A1(n6776), .A2(n6777), .B1(n6778), .B2(n6779), .Y(n4916) );
	inv_1 U6884( .A(n7376), .Y(n6779) );
	nor2_1 U6885( .A(n6780), .B(n6781), .Y(n6778) );
	o22ai_1 U6886( .A1(n6777), .A2(n6782), .B1(n6783), .B2(n6784), .Y(n4915) );
	inv_1 U6887( .A(n7375), .Y(n6784) );
	nor2_1 U6888( .A(n6780), .B(n6785), .Y(n6783) );
	o22ai_1 U6889( .A1(n6777), .A2(n6786), .B1(n6787), .B2(n6788), .Y(n4914) );
	nor2_1 U6890( .A(n6780), .B(n6789), .Y(n6787) );
	and2_0 U6891( .A(n6790), .B(n5740), .X(n6780) );
	nand2_1 U6892( .A(n7265), .B(n6790), .Y(n6777) );
	or3_1 U6893( .A(n6791), .B(n6792), .C(n6793), .X(n6790) );
	o22ai_1 U6894( .A1(n6776), .A2(n6794), .B1(n6795), .B2(n6796), .Y(n4913) );
	nor2_1 U6895( .A(n6797), .B(n6781), .Y(n6795) );
	o22ai_1 U6896( .A1(n6782), .A2(n6794), .B1(n6798), .B2(n6799), .Y(n4912) );
	nor2_1 U6897( .A(n6797), .B(n6785), .Y(n6798) );
	o22ai_1 U6898( .A1(n6786), .A2(n6794), .B1(n6800), .B2(n6801), .Y(n4911) );
	inv_1 U6899( .A(n7727), .Y(n6801) );
	nor2_1 U6900( .A(n6797), .B(n6789), .Y(n6800) );
	a21oi_1 U6901( .A1(n6802), .A2(n6803), .B1(RST), .Y(n6797) );
	inv_1 U6902( .A(n6804), .Y(n6802) );
	o21ai_0 U6903( .A1(n6804), .A2(n6791), .B1(n6805), .Y(n6794) );
	mux2i_1 U6904( .A0(n6793), .A1(n6806), .S(n6767), .Y(n6805) );
	a21oi_1 U6905( .A1(n6807), .A2(n7265), .B1(n6808), .Y(n6804) );
	and4_1 U6906( .A(n6809), .B(n6810), .C(n6811), .D(n6812), .X(n6808) );
	o22ai_1 U6907( .A1(n6813), .A2(n6814), .B1(n6776), .B2(n6815), .Y(n4910) );
	o22ai_1 U6908( .A1(n6816), .A2(n6817), .B1(n6782), .B2(n6815), .Y(n4909) );
	inv_1 U6909( .A(n7579), .Y(n6817) );
	o22ai_1 U6910( .A1(n6818), .A2(n5617), .B1(n6786), .B2(n6815), .Y(n4908) );
	nand2_1 U6911( .A(n6819), .B(n6820), .Y(n6815) );
	mux2i_1 U6912( .A0(n6821), .A1(n6822), .S(n6823), .Y(n6819) );
	nand2_1 U6913( .A(n6812), .B(n6822), .Y(n6821) );
	o211ai_1 U6914( .A1(n6809), .A2(n6824), .B1(n6812), .C1(n6825), .Y(n6822) );
	mux2i_1 U6915( .A0(n6826), .A1(n6827), .S(n6828), .Y(n6825) );
	a21oi_1 U6916( .A1(n6829), .A2(n6830), .B1(n6831), .Y(n6827) );
	nand2_1 U6917( .A(n6809), .B(n6811), .Y(n6830) );
	nand3_1 U6918( .A(n7265), .B(n6810), .C(n6809), .Y(n6826) );
	inv_1 U6919( .A(n6806), .Y(n6824) );
	nand2_1 U6920( .A(n6829), .B(n6811), .Y(n6806) );
	o22ai_1 U6921( .A1(n6813), .A2(n6832), .B1(n6776), .B2(n6833), .Y(n4907) );
	o22ai_1 U6922( .A1(n6816), .A2(n6834), .B1(n6782), .B2(n6833), .Y(n4906) );
	inv_1 U6923( .A(n7581), .Y(n6834) );
	o22ai_1 U6924( .A1(n6818), .A2(n5618), .B1(n6786), .B2(n6833), .Y(n4905) );
	nand2_1 U6925( .A(n6835), .B(n6820), .Y(n6833) );
	xnor2_1 U6926( .A(n6836), .B(n6837), .Y(n6835) );
	a21oi_1 U6927( .A1(n6838), .A2(n6812), .B1(n6839), .Y(n6837) );
	o22ai_1 U6928( .A1(n6840), .A2(n6841), .B1(n6842), .B2(n6828), .Y(n6838) );
	a21oi_1 U6929( .A1(n6843), .A2(n6803), .B1(n6831), .Y(n6842) );
	a21oi_1 U6930( .A1(n6844), .A2(n6809), .B1(n6845), .Y(n6843) );
	inv_1 U6931( .A(n6810), .Y(n6844) );
	a22oi_1 U6932( .A1(n6809), .A2(n6846), .B1(n6847), .B2(n6828), .Y(n6840) );
	xnor2_1 U6933( .A(n6836), .B(n6848), .Y(n6846) );
	nand2_1 U6934( .A(n6849), .B(n6811), .Y(n6848) );
	nand4_1 U6935( .A(n6850), .B(n6851), .C(n6852), .D(n6853), .Y(n6811) );
	nor3_1 U6936( .A(n6854), .B(n6855), .C(n6856), .Y(n6853) );
	or3_1 U6937( .A(n6857), .B(n6858), .C(n6859), .X(n6854) );
	nor3_1 U6938( .A(n6860), .B(n6861), .C(n6862), .Y(n6852) );
	inv_1 U6939( .A(n6863), .Y(n6849) );
	o22ai_1 U6940( .A1(n6813), .A2(n6864), .B1(n6776), .B2(n6865), .Y(n4904) );
	o22ai_1 U6941( .A1(n6816), .A2(n6866), .B1(n6782), .B2(n6865), .Y(n4903) );
	inv_1 U6942( .A(n7577), .Y(n6866) );
	o22ai_1 U6943( .A1(n6818), .A2(n5619), .B1(n6786), .B2(n6865), .Y(n4902) );
	o21ai_0 U6944( .A1(n6867), .A2(n6868), .B1(n6820), .Y(n6865) );
	nor3_1 U6945( .A(n6810), .B(n6869), .C(n6807), .Y(n6868) );
	o22ai_1 U6946( .A1(n6776), .A2(n6870), .B1(n6871), .B2(n6872), .Y(n4901) );
	inv_1 U6947( .A(n7312), .Y(n6872) );
	nor2_1 U6948( .A(n6873), .B(n6781), .Y(n6871) );
	o22ai_1 U6949( .A1(n6782), .A2(n6870), .B1(n6874), .B2(n6875), .Y(n4900) );
	inv_1 U6950( .A(n7311), .Y(n6875) );
	nor2_1 U6951( .A(n6873), .B(n6785), .Y(n6874) );
	inv_1 U6952( .A(n6876), .Y(n49) );
	o22ai_1 U6953( .A1(n6786), .A2(n6870), .B1(n6877), .B2(n6878), .Y(n4899) );
	nor2_1 U6954( .A(n6873), .B(n6789), .Y(n6877) );
	a21oi_1 U6955( .A1(n6879), .A2(n6880), .B1(RST), .Y(n6873) );
	inv_1 U6956( .A(n6881), .Y(n6880) );
	o211ai_1 U6957( .A1(n6769), .A2(n6882), .B1(n7265), .C1(n6883), .Y(n6870) );
	mux2i_1 U6958( .A0(n6882), .A1(n6769), .S(n6884), .Y(n6883) );
	o22ai_1 U6959( .A1(n5550), .A2(n6813), .B1(n6776), .B2(n6885), .Y(n4898) );
	o22ai_1 U6960( .A1(n5340), .A2(n6816), .B1(n6782), .B2(n6885), .Y(n4897) );
	o22ai_1 U6961( .A1(n6886), .A2(n6818), .B1(n6786), .B2(n6885), .Y(n4896) );
	xnor2_1 U6962( .A(n6887), .B(n6769), .Y(n6885) );
	nand2_1 U6963( .A(n6879), .B(n6881), .Y(n6887) );
	o221ai_1 U6964( .A1(n7311), .A2(n6774), .B1(n7312), .B2(n6888), .C1(n6889), .Y(n6881) );
	nand2_1 U6965( .A(g5511), .B(n6878), .Y(n6889) );
	inv_1 U6966( .A(n7714), .Y(n6878) );
	and2_0 U6967( .A(n6890), .B(n7265), .X(n6879) );
	mux2i_1 U6968( .A0(n6891), .A1(n6892), .S(n6884), .Y(n6890) );
	nand2_1 U6969( .A(n6769), .B(n6893), .Y(n6892) );
	inv_1 U6970( .A(n6894), .Y(n6769) );
	nand2_1 U6971( .A(n6882), .B(n6894), .Y(n6891) );
	o221ai_1 U6972( .A1(n6774), .A2(n5340), .B1(n6888), .B2(n5550), .C1(n6895), .Y(n6894) );
	nand2_1 U6973( .A(n7633), .B(g5511), .Y(n6895) );
	inv_1 U6974( .A(n7633), .Y(n6886) );
	o22ai_1 U6975( .A1(n6813), .A2(n5562), .B1(n6896), .B2(n6776), .Y(n4895) );
	o22ai_1 U6976( .A1(n6816), .A2(n5620), .B1(n6896), .B2(n6782), .Y(n4894) );
	o22ai_1 U6977( .A1(n6818), .A2(n6897), .B1(n6896), .B2(n6786), .Y(n4893) );
	mux2i_1 U6978( .A0(n6893), .A1(n6884), .S(n6793), .Y(n6896) );
	o21ai_0 U6979( .A1(n6888), .A2(n5562), .B1(n6898), .Y(n6884) );
	a22oi_1 U6980( .A1(n7629), .A2(g5511), .B1(n9792), .B2(g7014), .Y(n6898) );
	inv_1 U6981( .A(n6882), .Y(n6893) );
	o21ai_0 U6982( .A1(n6899), .A2(n6900), .B1(n6901), .Y(n6882) );
	inv_1 U6983( .A(n6902), .Y(n6901) );
	o22ai_1 U6984( .A1(n9968), .A2(n6903), .B1(n7385), .B2(n6904), .Y(n6900) );
	nor2_1 U6985( .A(n7386), .B(n6905), .Y(n6899) );
	inv_1 U6986( .A(n7629), .Y(n6897) );
	o22ai_1 U6987( .A1(n6776), .A2(n6906), .B1(n6907), .B2(n6908), .Y(n4892) );
	inv_1 U6988( .A(n7338), .Y(n6908) );
	nor2_1 U6989( .A(n6909), .B(n6781), .Y(n6907) );
	o22ai_1 U6990( .A1(n6782), .A2(n6906), .B1(n6910), .B2(n6911), .Y(n4891) );
	inv_1 U6991( .A(n7337), .Y(n6911) );
	nor2_1 U6992( .A(n6909), .B(n6785), .Y(n6910) );
	o22ai_1 U6993( .A1(n6786), .A2(n6906), .B1(n6912), .B2(n6913), .Y(n4890) );
	nor2_1 U6994( .A(n6909), .B(n6789), .Y(n6912) );
	a21oi_1 U6995( .A1(n6914), .A2(n6915), .B1(RST), .Y(n6909) );
	o22ai_1 U6996( .A1(n5551), .A2(n6813), .B1(n6916), .B2(n6776), .Y(n4889) );
	o22ai_1 U6997( .A1(n5341), .A2(n6816), .B1(n6916), .B2(n6782), .Y(n4888) );
	o22ai_1 U6998( .A1(n6917), .A2(n6818), .B1(n6916), .B2(n6786), .Y(n4887) );
	xnor2_1 U6999( .A(n6775), .B(n6918), .Y(n6916) );
	a21oi_1 U7000( .A1(n6831), .A2(n6919), .B1(n6920), .Y(n6918) );
	nor4_1 U7001( .A(n6921), .B(n6915), .C(n6793), .D(n6922), .Y(n6920) );
	inv_1 U7002( .A(n6923), .Y(n6915) );
	inv_1 U7003( .A(n7623), .Y(n6917) );
	o22ai_1 U7004( .A1(n6924), .A2(n6776), .B1(n6813), .B2(n5668), .Y(n4886) );
	inv_1 U7005( .A(n6781), .Y(n6813) );
	nor2_1 U7006( .A(n7782), .B(RST), .Y(n6781) );
	nand2_1 U7007( .A(n7782), .B(n5741), .Y(n6776) );
	o22ai_1 U7008( .A1(n6924), .A2(n6782), .B1(n6816), .B2(n5669), .Y(n4885) );
	inv_1 U7009( .A(n6785), .Y(n6816) );
	nor2_1 U7010( .A(g7014), .B(RST), .Y(n6785) );
	inv_1 U7011( .A(n172), .Y(n6782) );
	o22ai_1 U7012( .A1(n6924), .A2(n6786), .B1(n6818), .B2(n6925), .Y(n4884) );
	inv_1 U7013( .A(n6789), .Y(n6818) );
	nor2_1 U7014( .A(g5511), .B(RST), .Y(n6789) );
	inv_1 U7015( .A(n3959), .Y(n6786) );
	xnor2_1 U7016( .A(n6921), .B(n6926), .Y(n6924) );
	a21oi_1 U7017( .A1(n6927), .A2(n7265), .B1(n6928), .Y(n6926) );
	inv_1 U7018( .A(n6906), .Y(n6928) );
	nand2_1 U7019( .A(n6921), .B(n6914), .Y(n6906) );
	o32ai_1 U7020( .A1(n6793), .A2(n6775), .A3(n6929), .B1(n6831), .B2(n6930), .Y(n6914) );
	inv_1 U7021( .A(n6919), .Y(n6930) );
	nor3_1 U7022( .A(n6793), .B(n6759), .C(n6931), .Y(n6919) );
	inv_1 U7023( .A(n6929), .Y(n6931) );
	inv_1 U7024( .A(n7265), .Y(n6793) );
	a21oi_1 U7025( .A1(n6932), .A2(n6933), .B1(n6921), .Y(n6927) );
	inv_1 U7026( .A(n6922), .Y(n6933) );
	xnor2_1 U7027( .A(n6929), .B(n6759), .Y(n6922) );
	nor3_1 U7028( .A(n6934), .B(n6935), .C(n6902), .Y(n6929) );
	a21oi_1 U7029( .A1(n6831), .A2(n6775), .B1(n6923), .Y(n6932) );
	o221ai_1 U7030( .A1(n7337), .A2(n6774), .B1(n7338), .B2(n6888), .C1(n6936), .Y(n6923) );
	nand2_1 U7031( .A(g5511), .B(n6913), .Y(n6936) );
	inv_1 U7032( .A(n7733), .Y(n6913) );
	inv_1 U7033( .A(n6759), .Y(n6775) );
	o221ai_1 U7034( .A1(n6774), .A2(n5341), .B1(n6888), .B2(n5551), .C1(n6937), .Y(n6759) );
	nand2_1 U7035( .A(n7623), .B(g5511), .Y(n6937) );
	a221oi_1 U7036( .A1(g7014), .A2(n9793), .B1(n7782), .B2(n9986), .C1(n6938), .Y(n6921) );
	nor2_1 U7037( .A(n6925), .B(n6939), .Y(n6938) );
	inv_1 U7038( .A(n7625), .Y(n6925) );
	and2_0 U7039( .A(g5612), .B(n5759), .X(n4883) );
	nor2_1 U7040( .A(n6940), .B(n6941), .Y(n4882) );
	xnor2_1 U7041( .A(n10088), .B(n6942), .Y(n6940) );
	nor2_1 U7042( .A(n6943), .B(n6944), .Y(n6942) );
	nor2_1 U7043( .A(n6945), .B(n6941), .Y(n4881) );
	xnor2_1 U7044( .A(n6943), .B(n6944), .Y(n6945) );
	inv_1 U7045( .A(n7308), .Y(n6944) );
	nand2_1 U7046( .A(n7706), .B(n6946), .Y(n6943) );
	nor2_1 U7047( .A(n6947), .B(n6941), .Y(n4880) );
	xnor2_1 U7048( .A(n7706), .B(n6946), .Y(n6947) );
	a211oi_1 U7049( .A1(n5377), .A2(n6948), .B1(n6941), .C1(n6946), .Y(n4879) );
	nor2_1 U7050( .A(n5377), .B(n6948), .Y(n6946) );
	nor3_1 U7051( .A(n6941), .B(n6949), .C(n6950), .Y(n4878) );
	a21oi_1 U7052( .A1(n10086), .A2(n6951), .B1(n7697), .Y(n6950) );
	inv_1 U7053( .A(n6948), .Y(n6949) );
	nand3_1 U7054( .A(n7697), .B(n6951), .C(n10086), .Y(n6948) );
	nor2_1 U7055( .A(n6952), .B(n6941), .Y(n4877) );
	xnor2_1 U7056( .A(n10086), .B(n6951), .Y(n6952) );
	a211oi_1 U7057( .A1(n6953), .A2(n6954), .B1(n6941), .C1(n6951), .Y(n4876) );
	nor2_1 U7058( .A(n6953), .B(n6954), .Y(n6951) );
	inv_1 U7059( .A(n7710), .Y(n6953) );
	inv_1 U7060( .A(n6955), .Y(n4875) );
	o211ai_1 U7061( .A1(n10085), .A2(n6956), .B1(n6957), .C1(n6954), .Y(n6955) );
	nand2_1 U7062( .A(n10085), .B(n6956), .Y(n6954) );
	inv_1 U7063( .A(n6941), .Y(n6957) );
	nor3_1 U7064( .A(n6941), .B(n6956), .C(n6958), .Y(n4874) );
	a21oi_1 U7065( .A1(n9967), .A2(n6959), .B1(n7700), .Y(n6958) );
	and3_1 U7066( .A(n7700), .B(n6959), .C(n9967), .X(n6956) );
	nor2_1 U7067( .A(n6960), .B(n6941), .Y(n4873) );
	o21ai_0 U7068( .A1(n6131), .A2(n6961), .B1(n5741), .Y(n6941) );
	xnor2_1 U7069( .A(n6959), .B(n9967), .Y(n6960) );
	nor2_1 U7070( .A(n6903), .B(n6337), .Y(n6959) );
	o22ai_1 U7071( .A1(n6962), .A2(n6963), .B1(n6964), .B2(n6965), .Y(n4872) );
	o22ai_1 U7072( .A1(n5723), .A2(n6966), .B1(n6964), .B2(n6967), .Y(n4871) );
	o22ai_1 U7073( .A1(n5681), .A2(n6968), .B1(n6964), .B2(n6969), .Y(n4870) );
	o221ai_1 U7074( .A1(n6970), .A2(n6971), .B1(n6972), .B2(n6973), .C1(n6974), .Y(n6964) );
	xnor2_1 U7075( .A(n6975), .B(n6976), .Y(n6970) );
	nand2_1 U7076( .A(n6977), .B(n6978), .Y(n6975) );
	xnor2_1 U7077( .A(n6979), .B(n6980), .Y(n6978) );
	o22ai_1 U7078( .A1(n6981), .A2(n6963), .B1(n6982), .B2(n6965), .Y(n4869) );
	o22ai_1 U7079( .A1(n5533), .A2(n6966), .B1(n6982), .B2(n6967), .Y(n4868) );
	o22ai_1 U7080( .A1(n5699), .A2(n6968), .B1(n6982), .B2(n6969), .Y(n4867) );
	inv_1 U7081( .A(n6983), .Y(n6982) );
	o221ai_1 U7082( .A1(n6971), .A2(n6984), .B1(n6867), .B2(n6985), .C1(n6986), .Y(n6983) );
	nand2_1 U7083( .A(n6987), .B(n6988), .Y(n6986) );
	xnor2_1 U7084( .A(n6977), .B(n6989), .Y(n6984) );
	nor2_1 U7085( .A(n6990), .B(n6991), .Y(n6977) );
	mux2_1 U7086( .A0(n6992), .A1(n6993), .S(n6994), .X(n6990) );
	nand2_1 U7087( .A(n6867), .B(n6995), .Y(n6993) );
	nand2_1 U7088( .A(n6996), .B(n6980), .Y(n6992) );
	o22ai_1 U7089( .A1(n6997), .A2(n6963), .B1(n6998), .B2(n6965), .Y(n4866) );
	o22ai_1 U7090( .A1(n5724), .A2(n6966), .B1(n6998), .B2(n6967), .Y(n4865) );
	o22ai_1 U7091( .A1(n5682), .A2(n6968), .B1(n6998), .B2(n6969), .Y(n4864) );
	inv_1 U7092( .A(n6999), .Y(n6998) );
	o22ai_1 U7093( .A1(n5852), .A2(n6973), .B1(n6971), .B2(n7000), .Y(n6999) );
	xnor2_1 U7094( .A(n6994), .B(n7001), .Y(n7000) );
	nor2_1 U7095( .A(n7002), .B(n6991), .Y(n7001) );
	xnor2_1 U7096( .A(n6867), .B(n6996), .Y(n7002) );
	o22ai_1 U7097( .A1(n7003), .A2(n6963), .B1(n7004), .B2(n6965), .Y(n4863) );
	o22ai_1 U7098( .A1(n5534), .A2(n6966), .B1(n7004), .B2(n6967), .Y(n4862) );
	o22ai_1 U7099( .A1(n5700), .A2(n6968), .B1(n7004), .B2(n6969), .Y(n4861) );
	inv_1 U7100( .A(n7005), .Y(n7004) );
	o22ai_1 U7101( .A1(n5850), .A2(n6973), .B1(n6971), .B2(n7006), .Y(n7005) );
	xnor2_1 U7102( .A(n6991), .B(n6996), .Y(n7006) );
	nand2_1 U7103( .A(n7007), .B(n7008), .Y(n6991) );
	xnor2_1 U7104( .A(n7009), .B(n6867), .Y(n7008) );
	o22ai_1 U7105( .A1(n7010), .A2(n6963), .B1(n6965), .B2(n7011), .Y(n4860) );
	o22ai_1 U7106( .A1(n5725), .A2(n6966), .B1(n6967), .B2(n7011), .Y(n4859) );
	o22ai_1 U7107( .A1(n5683), .A2(n6968), .B1(n6969), .B2(n7011), .Y(n4858) );
	nand2_1 U7108( .A(n7012), .B(n6985), .Y(n7011) );
	mux2i_1 U7109( .A0(n7013), .A1(n5848), .S(n6971), .Y(n7012) );
	xnor2_1 U7110( .A(n7009), .B(n7007), .Y(n7013) );
	nor2_1 U7111( .A(n7014), .B(n7015), .Y(n7007) );
	xnor2_1 U7112( .A(n7016), .B(n6980), .Y(n7014) );
	o22ai_1 U7113( .A1(n7017), .A2(n6963), .B1(n7018), .B2(n6965), .Y(n4857) );
	o22ai_1 U7114( .A1(n5726), .A2(n6966), .B1(n7018), .B2(n6967), .Y(n4856) );
	o22ai_1 U7115( .A1(n5684), .A2(n6968), .B1(n7018), .B2(n6969), .Y(n4855) );
	inv_1 U7116( .A(n7019), .Y(n7018) );
	o22ai_1 U7117( .A1(n5846), .A2(n6973), .B1(n7020), .B2(n6971), .Y(n7019) );
	xnor2_1 U7118( .A(n7021), .B(n7015), .Y(n7020) );
	a22oi_1 U7119( .A1(n7022), .A2(n7023), .B1(n7024), .B2(n7025), .Y(n7015) );
	o22ai_1 U7120( .A1(n7026), .A2(n6963), .B1(n6965), .B2(n7027), .Y(n4854) );
	o22ai_1 U7121( .A1(n5531), .A2(n6966), .B1(n6967), .B2(n7027), .Y(n4853) );
	o22ai_1 U7122( .A1(n5701), .A2(n6968), .B1(n6969), .B2(n7027), .Y(n4852) );
	o221ai_1 U7123( .A1(n6971), .A2(n7028), .B1(n7271), .B2(n6973), .C1(n6974), .Y(n7027) );
	xnor2_1 U7124( .A(n7029), .B(n7030), .Y(n7028) );
	nor2_1 U7125( .A(n7031), .B(n7025), .Y(n7030) );
	nor3_1 U7126( .A(n7032), .B(n6867), .C(n7033), .Y(n7025) );
	nor3_1 U7127( .A(n7033), .B(n7034), .C(n6980), .Y(n7031) );
	o22ai_1 U7128( .A1(n7035), .A2(n6963), .B1(n7036), .B2(n6965), .Y(n4851) );
	o22ai_1 U7129( .A1(n5532), .A2(n6966), .B1(n7036), .B2(n6967), .Y(n4850) );
	o22ai_1 U7130( .A1(n5702), .A2(n6968), .B1(n7036), .B2(n6969), .Y(n4849) );
	inv_1 U7131( .A(n7037), .Y(n7036) );
	o221ai_1 U7132( .A1(n6971), .A2(n7038), .B1(n6867), .B2(n6985), .C1(n7039), .Y(n7037) );
	nand2_1 U7133( .A(n6987), .B(n7246), .Y(n7039) );
	inv_1 U7134( .A(n6973), .Y(n6987) );
	xnor2_1 U7135( .A(n7023), .B(n7032), .Y(n7038) );
	inv_1 U7136( .A(n7033), .Y(n7023) );
	o211ai_1 U7137( .A1(n7040), .A2(n6980), .B1(n7041), .C1(n7042), .Y(n7033) );
	mux2i_1 U7138( .A0(n7040), .A1(n6980), .S(n7043), .Y(n7042) );
	o22ai_1 U7139( .A1(n7044), .A2(n6963), .B1(n6965), .B2(n7045), .Y(n4848) );
	o22ai_1 U7140( .A1(n5530), .A2(n6966), .B1(n6967), .B2(n7045), .Y(n4847) );
	o22ai_1 U7141( .A1(n5703), .A2(n6968), .B1(n6969), .B2(n7045), .Y(n4846) );
	o221ai_1 U7142( .A1(n7046), .A2(n6971), .B1(n7585), .B2(n6973), .C1(n6974), .Y(n7045) );
	or2_0 U7143( .A(n6985), .B(n6980), .X(n6974) );
	xnor2_1 U7144( .A(n7047), .B(n7043), .Y(n7046) );
	nand2_1 U7145( .A(n7048), .B(n7041), .Y(n7047) );
	xnor2_1 U7146( .A(n7049), .B(n6980), .Y(n7048) );
	o22ai_1 U7147( .A1(n7050), .A2(n6963), .B1(n7051), .B2(n6965), .Y(n4845) );
	nand2_1 U7148( .A(n7229), .B(n5741), .Y(n6965) );
	nand2_1 U7149( .A(n6903), .B(n5741), .Y(n6963) );
	o22ai_1 U7150( .A1(n7051), .A2(n6967), .B1(n5396), .B2(n6966), .Y(n4844) );
	nand2_1 U7151( .A(n6904), .B(n5741), .Y(n6966) );
	inv_1 U7152( .A(n170), .Y(n6967) );
	o22ai_1 U7153( .A1(n5704), .A2(n6968), .B1(n7051), .B2(n6969), .Y(n4843) );
	inv_1 U7154( .A(n169), .Y(n6969) );
	inv_1 U7155( .A(n7052), .Y(n7051) );
	o22ai_1 U7156( .A1(n5838), .A2(n6973), .B1(n7053), .B2(n6971), .Y(n7052) );
	xnor2_1 U7157( .A(n7054), .B(n7049), .Y(n7053) );
	nand2_1 U7158( .A(n6985), .B(n6971), .Y(n6973) );
	o221ai_1 U7159( .A1(n7054), .A2(n7055), .B1(n6869), .B2(n7056), .C1(n7057), .Y(n6971) );
	a21oi_1 U7160( .A1(n7058), .A2(n6803), .B1(n7059), .Y(n7057) );
	inv_1 U7161( .A(n6820), .Y(n7059) );
	a21oi_1 U7162( .A1(n6767), .A2(n7060), .B1(n6845), .Y(n7058) );
	a221oi_1 U7163( .A1(n6799), .A2(g7014), .B1(n6796), .B2(n7782), .C1(n7061), .Y(n6845) );
	nor2_1 U7164( .A(n6939), .B(n7727), .Y(n7061) );
	inv_1 U7165( .A(n7329), .Y(n6796) );
	inv_1 U7166( .A(n7330), .Y(n6799) );
	nand3_1 U7167( .A(n6810), .B(n6812), .C(n6836), .Y(n7060) );
	o21ai_0 U7168( .A1(n6847), .A2(n6863), .B1(n6829), .Y(n6810) );
	o221ai_1 U7169( .A1(n7062), .A2(n7063), .B1(n7064), .B2(n7065), .C1(n7066), .Y(n6863) );
	o221ai_1 U7170( .A1(n6858), .A2(n6855), .B1(n6857), .B2(n6859), .C1(n7067), .Y(n7066) );
	o22ai_1 U7171( .A1(n6858), .A2(n6859), .B1(n6855), .B2(n7067), .Y(n7065) );
	o22ai_1 U7172( .A1(n6859), .A2(n7067), .B1(n6857), .B2(n6855), .Y(n7063) );
	xnor2_1 U7173( .A(n7271), .B(n7024), .Y(n6855) );
	inv_1 U7174( .A(n7064), .Y(n6857) );
	xor2_1 U7175( .A(n7009), .B(n5848), .X(n7064) );
	inv_1 U7176( .A(n6850), .Y(n7067) );
	xor2_1 U7177( .A(n6934), .B(n6976), .X(n6850) );
	xnor2_1 U7178( .A(n6994), .B(n5852), .Y(n6859) );
	inv_1 U7179( .A(n6858), .Y(n7062) );
	xor2_1 U7180( .A(n7585), .B(n7043), .X(n6858) );
	o221ai_1 U7181( .A1(n6851), .A2(n7068), .B1(n7069), .B2(n7070), .C1(n7071), .Y(n6847) );
	o221ai_1 U7182( .A1(n6862), .A2(n7072), .B1(n6856), .B2(n6861), .C1(n6860), .Y(n7071) );
	o22ai_1 U7183( .A1(n6862), .A2(n6860), .B1(n6856), .B2(n7072), .Y(n7070) );
	o22ai_1 U7184( .A1(n6861), .A2(n6862), .B1(n6856), .B2(n6860), .Y(n7068) );
	xnor2_1 U7185( .A(n7243), .B(n7049), .Y(n6860) );
	xnor2_1 U7186( .A(n7246), .B(n7034), .Y(n6856) );
	xnor2_1 U7187( .A(n7234), .B(n6996), .Y(n6862) );
	inv_1 U7188( .A(n7069), .Y(n6861) );
	xnor2_1 U7189( .A(n7021), .B(n5846), .Y(n7069) );
	inv_1 U7190( .A(n7072), .Y(n6851) );
	xnor2_1 U7191( .A(n6935), .B(n6989), .Y(n7072) );
	inv_1 U7192( .A(n6807), .Y(n6767) );
	nor3_1 U7193( .A(n6869), .B(n6809), .C(n6828), .Y(n6807) );
	inv_1 U7194( .A(n6831), .Y(n7056) );
	nor2_1 U7195( .A(n7073), .B(n7074), .Y(n6831) );
	inv_1 U7196( .A(n7717), .Y(n7074) );
	inv_1 U7197( .A(n6812), .Y(n6869) );
	a21oi_1 U7198( .A1(n7075), .A2(n6980), .B1(n7076), .Y(n7055) );
	o211ai_1 U7199( .A1(n7075), .A2(n7076), .B1(n6820), .C1(n7041), .Y(n6985) );
	inv_1 U7200( .A(n7054), .Y(n7041) );
	nor2_1 U7201( .A(n6867), .B(n6839), .Y(n7054) );
	nand2_1 U7202( .A(n6803), .B(n6792), .Y(n6820) );
	o221ai_1 U7203( .A1(n7375), .A2(n6774), .B1(n7376), .B2(n6888), .C1(n7077), .Y(n6792) );
	nand2_1 U7204( .A(g5511), .B(n6788), .Y(n7077) );
	inv_1 U7205( .A(n7738), .Y(n6788) );
	inv_1 U7206( .A(n6791), .Y(n6803) );
	nand2_1 U7207( .A(n7078), .B(n7079), .Y(n6791) );
	nor4_1 U7208( .A(n7080), .B(n7081), .C(n7082), .D(n7083), .Y(n7079) );
	xnor2_1 U7209( .A(n7084), .B(n6972), .Y(n7083) );
	a222oi_1 U7210( .A1(g6782), .A2(n7085), .B1(n7229), .B2(n5429), .C1(g6573), .C2(n7086), .Y(n7084) );
	xnor2_1 U7211( .A(n7087), .B(n6988), .Y(n7082) );
	a222oi_1 U7212( .A1(g6782), .A2(n7088), .B1(n7229), .B2(n5430), .C1(g6573), .C2(n7089), .Y(n7087) );
	mux2i_1 U7213( .A0(n7090), .A1(n7091), .S(n5848), .Y(n7081) );
	nand2_1 U7214( .A(n7322), .B(n7091), .Y(n7090) );
	nand3_1 U7215( .A(n7092), .B(n7093), .C(n6829), .Y(n7080) );
	inv_1 U7216( .A(n6841), .Y(n6829) );
	nand2_1 U7217( .A(n7717), .B(n7073), .Y(n6841) );
	o21ai_0 U7218( .A1(n9987), .A2(n6903), .B1(n7094), .Y(n7073) );
	a22oi_1 U7219( .A1(g6573), .A2(n7095), .B1(g6782), .B2(n7096), .Y(n7094) );
	xnor2_1 U7220( .A(n5838), .B(n7097), .Y(n7093) );
	a222oi_1 U7221( .A1(g6782), .A2(n7098), .B1(n7229), .B2(n5439), .C1(g6573), .C2(n7099), .Y(n7097) );
	xnor2_1 U7222( .A(n5840), .B(n7100), .Y(n7092) );
	a222oi_1 U7223( .A1(g6782), .A2(n7101), .B1(n7229), .B2(n5431), .C1(g6573), .C2(n7102), .Y(n7100) );
	nor4_1 U7224( .A(n7103), .B(n7104), .C(n7105), .D(n7106), .Y(n7078) );
	mux2i_1 U7225( .A0(n7107), .A1(n7108), .S(n5844), .Y(n7106) );
	nand2_1 U7226( .A(n7614), .B(n7108), .Y(n7107) );
	mux2i_1 U7227( .A0(n7109), .A1(n7110), .S(n5850), .Y(n7105) );
	nand2_1 U7228( .A(n7611), .B(n7110), .Y(n7109) );
	mux2i_1 U7229( .A0(n7111), .A1(n7112), .S(n5852), .Y(n7104) );
	nand2_1 U7230( .A(n7610), .B(n7112), .Y(n7111) );
	nand3_1 U7231( .A(n7113), .B(n7114), .C(n7115), .Y(n7103) );
	mux2i_1 U7232( .A0(n7116), .A1(n7117), .S(n5842), .Y(n7115) );
	nor2_1 U7233( .A(n7117), .B(n7118), .Y(n7116) );
	mux2i_1 U7234( .A0(n7119), .A1(n7120), .S(n6903), .Y(n7114) );
	nand2_1 U7235( .A(n7121), .B(n7122), .Y(n7120) );
	a222oi_1 U7236( .A1(n7112), .A2(n7268), .B1(n7091), .B2(n7221), .C1(n7108), .C2(n7271), .Y(n7122) );
	a22oi_1 U7237( .A1(n5491), .A2(g6782), .B1(n5322), .B2(g6573), .Y(n7108) );
	a22oi_1 U7238( .A1(n5490), .A2(g6782), .B1(n5321), .B2(g6573), .Y(n7091) );
	a22oi_1 U7239( .A1(n5488), .A2(g6782), .B1(n5319), .B2(g6573), .Y(n7112) );
	a222oi_1 U7240( .A1(n7123), .A2(n7246), .B1(n7110), .B2(n7234), .C1(n7124), .C2(n7274), .Y(n7121) );
	inv_1 U7241( .A(n7125), .Y(n7124) );
	a22oi_1 U7242( .A1(n5489), .A2(g6782), .B1(n5320), .B2(g6573), .Y(n7110) );
	inv_1 U7243( .A(n7117), .Y(n7123) );
	o22ai_1 U7244( .A1(n9796), .A2(n6904), .B1(n9797), .B2(n6905), .Y(n7117) );
	nand2_1 U7245( .A(n7126), .B(n7127), .Y(n7119) );
	a222oi_1 U7246( .A1(n5842), .A2(n7118), .B1(n5848), .B2(n7128), .C1(n5850), .C2(n7129), .Y(n7127) );
	a222oi_1 U7247( .A1(n5846), .A2(n5360), .B1(n5852), .B2(n7130), .C1(n5844), .C2(n7131), .Y(n7126) );
	mux2i_1 U7248( .A0(n7132), .A1(n7125), .S(n5846), .Y(n7113) );
	nor2_1 U7249( .A(n7125), .B(n5360), .Y(n7132) );
	o22ai_1 U7250( .A1(n9794), .A2(n6904), .B1(n9795), .B2(n6905), .Y(n7125) );
	and3_1 U7251( .A(n7022), .B(n7133), .C(n7134), .X(n7076) );
	and3_1 U7252( .A(n6989), .B(n7043), .C(n6976), .X(n7134) );
	nor3_1 U7253( .A(n7034), .B(n7024), .C(n6980), .Y(n7022) );
	inv_1 U7254( .A(n6867), .Y(n6980) );
	nor3_1 U7255( .A(n6823), .B(n6836), .C(n6812), .Y(n6867) );
	nand2_1 U7256( .A(n6905), .B(n5741), .Y(n6968) );
	o22ai_1 U7257( .A1(n7135), .A2(n5602), .B1(n7136), .B2(n7137), .Y(n4842) );
	o22ai_1 U7258( .A1(n7138), .A2(n7139), .B1(n7137), .B2(n7140), .Y(n4841) );
	inv_1 U7259( .A(n7385), .Y(n7139) );
	o22ai_1 U7260( .A1(n7141), .A2(n7142), .B1(n7137), .B2(n7143), .Y(n4840) );
	nand2_1 U7261( .A(n6902), .B(n5742), .Y(n7137) );
	nand2_1 U7262( .A(n7144), .B(n7145), .Y(n6902) );
	nor4_1 U7263( .A(n5838), .B(n5840), .C(n5842), .D(n5844), .Y(n7145) );
	inv_1 U7264( .A(n7271), .Y(n5844) );
	inv_1 U7265( .A(n7246), .Y(n5842) );
	inv_1 U7266( .A(n7585), .Y(n5840) );
	inv_1 U7267( .A(n7243), .Y(n5838) );
	nor4_1 U7268( .A(n5846), .B(n5848), .C(n5850), .D(n5852), .Y(n7144) );
	inv_1 U7269( .A(n7268), .Y(n5852) );
	inv_1 U7270( .A(n7221), .Y(n5848) );
	inv_1 U7271( .A(n7274), .Y(n5846) );
	inv_1 U7272( .A(n7386), .Y(n7142) );
	o22ai_1 U7273( .A1(n7136), .A2(n7146), .B1(n7135), .B2(n7147), .Y(n4839) );
	inv_1 U7274( .A(n7426), .Y(n7147) );
	o22ai_1 U7275( .A1(n7140), .A2(n7146), .B1(n7138), .B2(n5411), .Y(n4838) );
	o22ai_1 U7276( .A1(n7143), .A2(n7146), .B1(n7141), .B2(n7148), .Y(n4837) );
	o22ai_1 U7277( .A1(n7136), .A2(n7149), .B1(n7135), .B2(n7150), .Y(n4836) );
	inv_1 U7278( .A(n7418), .Y(n7150) );
	o22ai_1 U7279( .A1(n7140), .A2(n7149), .B1(n7138), .B2(n7151), .Y(n4835) );
	o22ai_1 U7280( .A1(n7143), .A2(n7149), .B1(n7141), .B2(n5399), .Y(n4834) );
	o22ai_1 U7281( .A1(n7136), .A2(n7152), .B1(n7135), .B2(n5676), .Y(n4833) );
	nand2_1 U7282( .A(n7136), .B(n5743), .Y(n7135) );
	nand2_1 U7283( .A(n7229), .B(n6529), .Y(n7136) );
	o22ai_1 U7284( .A1(n7140), .A2(n7152), .B1(n7138), .B2(n7096), .Y(n4832) );
	inv_1 U7285( .A(n7392), .Y(n7096) );
	nand2_1 U7286( .A(n7140), .B(n5743), .Y(n7138) );
	nand2_1 U7287( .A(g6782), .B(n6529), .Y(n7140) );
	o22ai_1 U7288( .A1(n7143), .A2(n7152), .B1(n7141), .B2(n7095), .Y(n4831) );
	inv_1 U7289( .A(n7394), .Y(n7095) );
	nand2_1 U7290( .A(n7143), .B(n5743), .Y(n7141) );
	nand4_1 U7291( .A(n5), .B(n7268), .C(n7274), .D(n5850), .Y(n7152) );
	inv_1 U7292( .A(n7234), .Y(n5850) );
	nand2_1 U7293( .A(g6573), .B(n6529), .Y(n7143) );
	o22ai_1 U7294( .A1(n7153), .A2(n5429), .B1(n6961), .B2(n7154), .Y(n4830) );
	o22ai_1 U7295( .A1(n7155), .A2(n7085), .B1(n7154), .B2(n7156), .Y(n4829) );
	inv_1 U7296( .A(n7409), .Y(n7085) );
	o22ai_1 U7297( .A1(n7157), .A2(n7086), .B1(n7154), .B2(n7158), .Y(n4828) );
	nand2_1 U7298( .A(n6934), .B(n5743), .Y(n7154) );
	inv_1 U7299( .A(n6972), .Y(n6934) );
	o21ai_0 U7300( .A1(n7418), .A2(n6903), .B1(n7159), .Y(n6972) );
	a22oi_1 U7301( .A1(g6573), .A2(n5399), .B1(g6782), .B2(n7151), .Y(n7159) );
	inv_1 U7302( .A(n7417), .Y(n7151) );
	inv_1 U7303( .A(n7416), .Y(n7086) );
	o22ai_1 U7304( .A1(n7153), .A2(n5430), .B1(n6961), .B2(n7160), .Y(n4827) );
	o22ai_1 U7305( .A1(n7155), .A2(n7088), .B1(n7156), .B2(n7160), .Y(n4826) );
	inv_1 U7306( .A(n7419), .Y(n7088) );
	o22ai_1 U7307( .A1(n7157), .A2(n7089), .B1(n7158), .B2(n7160), .Y(n4825) );
	nand2_1 U7308( .A(n6935), .B(n5743), .Y(n7160) );
	inv_1 U7309( .A(n6988), .Y(n6935) );
	o21ai_0 U7310( .A1(n7426), .A2(n6903), .B1(n7161), .Y(n6988) );
	a22oi_1 U7311( .A1(g6573), .A2(n7148), .B1(g6782), .B2(n5411), .Y(n7161) );
	inv_1 U7312( .A(n7427), .Y(n7148) );
	inv_1 U7313( .A(n7425), .Y(n7089) );
	o22ai_1 U7314( .A1(n6961), .A2(n7162), .B1(n7130), .B2(n7153), .Y(n4824) );
	inv_1 U7315( .A(n7610), .Y(n7130) );
	o22ai_1 U7316( .A1(n7156), .A2(n7162), .B1(n7155), .B2(n5488), .Y(n4823) );
	o22ai_1 U7317( .A1(n7158), .A2(n7162), .B1(n7157), .B2(n5319), .Y(n4822) );
	inv_1 U7318( .A(n171), .Y(n7162) );
	o22ai_1 U7319( .A1(n6961), .A2(n7163), .B1(n7129), .B2(n7153), .Y(n4821) );
	inv_1 U7320( .A(n7611), .Y(n7129) );
	o22ai_1 U7321( .A1(n7156), .A2(n7163), .B1(n7155), .B2(n5489), .Y(n4820) );
	o22ai_1 U7322( .A1(n7158), .A2(n7163), .B1(n7157), .B2(n5320), .Y(n4819) );
	inv_1 U7323( .A(n4), .Y(n7163) );
	o22ai_1 U7324( .A1(n6961), .A2(n7164), .B1(n7128), .B2(n7153), .Y(n4818) );
	inv_1 U7325( .A(n7322), .Y(n7128) );
	o22ai_1 U7326( .A1(n7164), .A2(n7156), .B1(n7155), .B2(n5490), .Y(n4817) );
	o22ai_1 U7327( .A1(n7164), .A2(n7158), .B1(n7157), .B2(n5321), .Y(n4816) );
	inv_1 U7328( .A(n5), .Y(n7164) );
	nor2_1 U7329( .A(RST), .B(n7221), .Y(n5) );
	o22ai_1 U7330( .A1(n6961), .A2(n7165), .B1(n5360), .B2(n7153), .Y(n4815) );
	o22ai_1 U7331( .A1(n7156), .A2(n7165), .B1(n7155), .B2(n5651), .Y(n4814) );
	o22ai_1 U7332( .A1(n7158), .A2(n7165), .B1(n7157), .B2(n5637), .Y(n4813) );
	inv_1 U7333( .A(n6), .Y(n7165) );
	nor2_1 U7334( .A(RST), .B(n7274), .Y(n6) );
	o22ai_1 U7335( .A1(n6961), .A2(n7166), .B1(n7131), .B2(n7153), .Y(n4812) );
	inv_1 U7336( .A(n7614), .Y(n7131) );
	o22ai_1 U7337( .A1(n7156), .A2(n7166), .B1(n7155), .B2(n5491), .Y(n4811) );
	o22ai_1 U7338( .A1(n7158), .A2(n7166), .B1(n7157), .B2(n5322), .Y(n4810) );
	inv_1 U7339( .A(n7), .Y(n7166) );
	nor2_1 U7340( .A(RST), .B(n7271), .Y(n7) );
	o22ai_1 U7341( .A1(n6961), .A2(n7167), .B1(n7118), .B2(n7153), .Y(n4809) );
	inv_1 U7342( .A(n7324), .Y(n7118) );
	o22ai_1 U7343( .A1(n7156), .A2(n7167), .B1(n7155), .B2(n5652), .Y(n4808) );
	o22ai_1 U7344( .A1(n7158), .A2(n7167), .B1(n7157), .B2(n5638), .Y(n4807) );
	inv_1 U7345( .A(n8), .Y(n7167) );
	nor2_1 U7346( .A(RST), .B(n7246), .Y(n8) );
	o22ai_1 U7347( .A1(n7153), .A2(n5431), .B1(n6961), .B2(n7149), .Y(n4806) );
	o22ai_1 U7348( .A1(n7155), .A2(n7101), .B1(n7149), .B2(n7156), .Y(n4805) );
	inv_1 U7349( .A(n7403), .Y(n7101) );
	o22ai_1 U7350( .A1(n7157), .A2(n7102), .B1(n7149), .B2(n7158), .Y(n4804) );
	inv_1 U7351( .A(n9), .Y(n7149) );
	nor2_1 U7352( .A(n7585), .B(RST), .Y(n9) );
	inv_1 U7353( .A(n7410), .Y(n7102) );
	o22ai_1 U7354( .A1(n6961), .A2(n7146), .B1(n7153), .B2(n5439), .Y(n4803) );
	nand2_1 U7355( .A(n5757), .B(n6961), .Y(n7153) );
	nand2_1 U7356( .A(n7717), .B(n7229), .Y(n6961) );
	o22ai_1 U7357( .A1(n7146), .A2(n7156), .B1(n7155), .B2(n7098), .Y(n4802) );
	inv_1 U7358( .A(n7411), .Y(n7098) );
	nand2_1 U7359( .A(n5757), .B(n7156), .Y(n7155) );
	nand2_1 U7360( .A(n7717), .B(g6782), .Y(n7156) );
	o22ai_1 U7361( .A1(n7146), .A2(n7158), .B1(n7157), .B2(n7099), .Y(n4801) );
	inv_1 U7362( .A(n7420), .Y(n7099) );
	nand2_1 U7363( .A(n5757), .B(n7158), .Y(n7157) );
	nand2_1 U7364( .A(n7717), .B(g6573), .Y(n7158) );
	inv_1 U7365( .A(n10), .Y(n7146) );
	a21oi_1 U7366( .A1(n7168), .A2(n7169), .B1(n7170), .Y(n4800) );
	nor2_1 U7367( .A(n6264), .B(RST), .Y(n48) );
	a21oi_1 U7368( .A1(n5335), .A2(n7171), .B1(n7172), .Y(n4799) );
	a21oi_1 U7369( .A1(n5544), .A2(n7173), .B1(n7174), .Y(n4798) );
	o22ai_1 U7370( .A1(n7175), .A2(n7176), .B1(n7177), .B2(n7178), .Y(n4797) );
	inv_1 U7371( .A(n7523), .Y(n7176) );
	o22ai_1 U7372( .A1(n7179), .A2(n7180), .B1(n7177), .B2(n7181), .Y(n4796) );
	inv_1 U7373( .A(n7546), .Y(n7180) );
	o22ai_1 U7374( .A1(n7182), .A2(n7183), .B1(n7177), .B2(n7184), .Y(n4795) );
	nand4_1 U7375( .A(n7185), .B(n7186), .C(n7187), .D(n7188), .Y(n7177) );
	a222oi_1 U7376( .A1(g7161), .A2(n7189), .B1(n7238), .B2(n7190), .C1(g6979), .C2(n5392), .Y(n7188) );
	nand2_1 U7377( .A(n9867), .B(n9988), .Y(n7190) );
	nand4_1 U7378( .A(n7191), .B(n7192), .C(n7193), .D(n7194), .Y(n7187) );
	nor3_1 U7379( .A(n7195), .B(n7196), .C(n7197), .Y(n7194) );
	xor2_1 U7380( .A(n7198), .B(n9990), .X(n7197) );
	xor2_1 U7381( .A(n7199), .B(n7691), .X(n7196) );
	nand3_1 U7382( .A(n7200), .B(n7201), .C(n7202), .Y(n7195) );
	xor2_1 U7383( .A(n9953), .B(n7203), .X(n7202) );
	xnor2_1 U7384( .A(n9991), .B(n7204), .Y(n7201) );
	xnor2_1 U7385( .A(n9992), .B(n7205), .Y(n7200) );
	nor3_1 U7386( .A(n7206), .B(n7207), .C(n7208), .Y(n7193) );
	xor2_1 U7387( .A(n7209), .B(n9969), .X(n7208) );
	xor2_1 U7388( .A(n7210), .B(n9989), .X(n7207) );
	xnor2_1 U7389( .A(n7211), .B(n7212), .Y(n7206) );
	xnor2_1 U7390( .A(n7297), .B(n7213), .Y(n7192) );
	xnor2_1 U7391( .A(n7693), .B(n7214), .Y(n7191) );
	o22ai_1 U7392( .A1(n7170), .A2(n5572), .B1(n7215), .B2(n7216), .Y(n4794) );
	o22ai_1 U7393( .A1(n7172), .A2(n7217), .B1(n7215), .B2(n7218), .Y(n4793) );
	o22ai_1 U7394( .A1(n7174), .A2(n5458), .B1(n7215), .B2(n5814), .Y(n4792) );
	nand2_1 U7395( .A(n7219), .B(n9970), .Y(n7215) );
	o22ai_1 U7396( .A1(n7170), .A2(n5621), .B1(n7216), .B2(n7220), .Y(n4791) );
	o21ai_0 U7397( .A1(n5363), .A2(n7253), .B1(n5742), .Y(n7170) );
	o22ai_1 U7398( .A1(n7172), .A2(n7189), .B1(n7218), .B2(n7220), .Y(n4790) );
	inv_1 U7399( .A(n5295), .Y(n7218) );
	nor2_1 U7400( .A(n7746), .B(RST), .Y(n5295) );
	inv_1 U7401( .A(n7449), .Y(n7189) );
	o22ai_1 U7402( .A1(n7174), .A2(n5392), .B1(n5814), .B2(n7220), .Y(n4789) );
	nand2_1 U7403( .A(n7747), .B(n9970), .Y(n7220) );
	nand2_1 U7404( .A(g6979), .B(n5743), .Y(n5814) );
	o21ai_0 U7405( .A1(n5363), .A2(n7748), .B1(n5758), .Y(n7174) );
	o22ai_1 U7406( .A1(n7175), .A2(n7749), .B1(n9991), .B2(n7178), .Y(n4788) );
	inv_1 U7407( .A(n7525), .Y(n7749) );
	o22ai_1 U7408( .A1(n7179), .A2(n7750), .B1(n9991), .B2(n7181), .Y(n4787) );
	inv_1 U7409( .A(n7524), .Y(n7750) );
	o22ai_1 U7410( .A1(n7182), .A2(n5453), .B1(n9991), .B2(n7184), .Y(n4786) );
	o22ai_1 U7411( .A1(n7175), .A2(n7751), .B1(n9992), .B2(n7178), .Y(n4785) );
	inv_1 U7412( .A(n7527), .Y(n7751) );
	o22ai_1 U7413( .A1(n7179), .A2(n7752), .B1(n9992), .B2(n7181), .Y(n4784) );
	inv_1 U7414( .A(n7526), .Y(n7752) );
	o22ai_1 U7415( .A1(n7182), .A2(n5456), .B1(n9992), .B2(n7184), .Y(n4783) );
	o22ai_1 U7416( .A1(n7175), .A2(n7753), .B1(n7693), .B2(n7178), .Y(n4782) );
	inv_1 U7417( .A(n7536), .Y(n7753) );
	o22ai_1 U7418( .A1(n7179), .A2(n7754), .B1(n7693), .B2(n7181), .Y(n4781) );
	inv_1 U7419( .A(n7535), .Y(n7754) );
	o22ai_1 U7420( .A1(n7182), .A2(n5462), .B1(n7693), .B2(n7184), .Y(n4780) );
	o22ai_1 U7421( .A1(n7175), .A2(n7755), .B1(n9989), .B2(n7178), .Y(n4779) );
	inv_1 U7422( .A(n7538), .Y(n7755) );
	o22ai_1 U7423( .A1(n7179), .A2(n7756), .B1(n9989), .B2(n7181), .Y(n4778) );
	inv_1 U7424( .A(n7537), .Y(n7756) );
	o22ai_1 U7425( .A1(n7182), .A2(n5459), .B1(n9989), .B2(n7184), .Y(n4777) );
	o22ai_1 U7426( .A1(n7175), .A2(n7757), .B1(n7297), .B2(n7178), .Y(n4776) );
	inv_1 U7427( .A(n7540), .Y(n7757) );
	o22ai_1 U7428( .A1(n7179), .A2(n7758), .B1(n7297), .B2(n7181), .Y(n4775) );
	inv_1 U7429( .A(n7539), .Y(n7758) );
	o22ai_1 U7430( .A1(n7182), .A2(n5460), .B1(n7297), .B2(n7184), .Y(n4774) );
	o22ai_1 U7431( .A1(n7175), .A2(n7759), .B1(n9990), .B2(n7178), .Y(n4773) );
	inv_1 U7432( .A(n7542), .Y(n7759) );
	o22ai_1 U7433( .A1(n7179), .A2(n7760), .B1(n9990), .B2(n7181), .Y(n4772) );
	inv_1 U7434( .A(n7541), .Y(n7760) );
	o22ai_1 U7435( .A1(n7182), .A2(n5457), .B1(n9990), .B2(n7184), .Y(n4771) );
	o22ai_1 U7436( .A1(n7175), .A2(n7761), .B1(n7301), .B2(n7178), .Y(n4770) );
	inv_1 U7437( .A(n7533), .Y(n7761) );
	o22ai_1 U7438( .A1(n7179), .A2(n7762), .B1(n7301), .B2(n7181), .Y(n4769) );
	inv_1 U7439( .A(n7532), .Y(n7762) );
	o22ai_1 U7440( .A1(n7182), .A2(n5455), .B1(n7301), .B2(n7184), .Y(n4768) );
	o22ai_1 U7441( .A1(n7175), .A2(n7763), .B1(n9953), .B2(n7178), .Y(n4767) );
	o22ai_1 U7442( .A1(n7179), .A2(n7764), .B1(n9953), .B2(n7181), .Y(n4766) );
	o22ai_1 U7443( .A1(n7182), .A2(n5622), .B1(n9953), .B2(n7184), .Y(n4765) );
	o22ai_1 U7444( .A1(n7175), .A2(n7765), .B1(n7691), .B2(n7178), .Y(n4764) );
	inv_1 U7445( .A(n7531), .Y(n7765) );
	o22ai_1 U7446( .A1(n7179), .A2(n7766), .B1(n7691), .B2(n7181), .Y(n4763) );
	inv_1 U7447( .A(n7530), .Y(n7766) );
	o22ai_1 U7448( .A1(n7182), .A2(n5454), .B1(n7691), .B2(n7184), .Y(n4762) );
	o22ai_1 U7449( .A1(n7175), .A2(n7767), .B1(n9969), .B2(n7178), .Y(n4761) );
	or2_0 U7450( .A(n7169), .B(RST), .X(n7178) );
	inv_1 U7451( .A(n7544), .Y(n7767) );
	nand2_1 U7452( .A(n5757), .B(n7169), .Y(n7175) );
	nand3_1 U7453( .A(n9971), .B(n7768), .C(n9866), .Y(n7169) );
	o22ai_1 U7454( .A1(n7179), .A2(n7769), .B1(n9969), .B2(n7181), .Y(n4760) );
	or2_0 U7455( .A(n7171), .B(RST), .X(n7181) );
	inv_1 U7456( .A(n7543), .Y(n7769) );
	nand2_1 U7457( .A(n5757), .B(n7171), .Y(n7179) );
	nand2_1 U7458( .A(n7770), .B(g7161), .Y(n7171) );
	o22ai_1 U7459( .A1(n7182), .A2(n5461), .B1(n9969), .B2(n7184), .Y(n4759) );
	or2_0 U7460( .A(n7173), .B(RST), .X(n7184) );
	nand2_1 U7461( .A(n5757), .B(n7173), .Y(n7182) );
	nand2_1 U7462( .A(n7770), .B(g6979), .Y(n7173) );
	and3_1 U7463( .A(n9971), .B(n7771), .C(n9866), .X(n7770) );
	nor2_1 U7464( .A(n7772), .B(n7172), .Y(n4758) );
	xnor2_1 U7465( .A(n7773), .B(n9991), .Y(n7772) );
	a211oi_1 U7466( .A1(n5367), .A2(n7774), .B1(n7172), .C1(n7773), .Y(n4757) );
	nor2_1 U7467( .A(n7774), .B(n5367), .Y(n7773) );
	nor3_1 U7468( .A(n7172), .B(n7776), .C(n7777), .Y(n4756) );
	a21oi_1 U7469( .A1(n7778), .A2(n9989), .B1(n7693), .Y(n7777) );
	inv_1 U7470( .A(n7774), .Y(n7776) );
	nand3_1 U7471( .A(n7693), .B(n9989), .C(n7778), .Y(n7774) );
	nor2_1 U7472( .A(n7779), .B(n7172), .Y(n4755) );
	xnor2_1 U7473( .A(n7778), .B(n9989), .Y(n7779) );
	nor3_1 U7474( .A(n7172), .B(n7778), .C(n7781), .Y(n4754) );
	a21oi_1 U7475( .A1(n7783), .A2(n9990), .B1(n7297), .Y(n7781) );
	and3_1 U7476( .A(n7297), .B(n9990), .C(n7783), .X(n7778) );
	nor2_1 U7477( .A(n7785), .B(n7172), .Y(n4753) );
	xnor2_1 U7478( .A(n9990), .B(n7783), .Y(n7785) );
	a211oi_1 U7479( .A1(n7212), .A2(n5813), .B1(n7172), .C1(n7783), .Y(n4752) );
	nor2_1 U7480( .A(n5813), .B(n7212), .Y(n7783) );
	nand2_1 U7481( .A(n9953), .B(n5811), .Y(n5813) );
	inv_1 U7482( .A(n7301), .Y(n7212) );
	nor3_1 U7483( .A(n7172), .B(n5811), .C(n7786), .Y(n4751) );
	a21oi_1 U7484( .A1(n9969), .A2(n7768), .B1(n7691), .Y(n7786) );
	and3_1 U7485( .A(n7691), .B(n7768), .C(n9969), .X(n5811) );
	nor2_1 U7486( .A(n7787), .B(n7172), .Y(n4750) );
	inv_1 U7487( .A(n5812), .Y(n7172) );
	a21oi_1 U7488( .A1(g7161), .A2(n9970), .B1(RST), .Y(n5812) );
	xnor2_1 U7489( .A(n7768), .B(n9969), .Y(n7787) );
	nor2_1 U7490( .A(n7253), .B(n7277), .Y(n7768) );
	o32ai_1 U7491( .A1(n7771), .A2(n7238), .A3(RST), .B1(n5981), .B2(n7216), .Y(n4749) );
	inv_1 U7492( .A(n7277), .Y(n7771) );
	o32ai_1 U7493( .A1(n5363), .A2(n7238), .A3(RST), .B1(n7216), .B2(n7788), .Y(n4748) );
	nand2_1 U7494( .A(n7238), .B(n5743), .Y(n7216) );
	o22ai_1 U7495( .A1(n5983), .A2(n7789), .B1(n5984), .B2(n5568), .Y(n4747) );
	and2_0 U7496( .A(n5757), .B(g16355), .X(n4746) );
	and2_0 U7497( .A(n5758), .B(n7790), .X(n4745) );
	o22ai_1 U7498( .A1(n5564), .A2(n7791), .B1(n7792), .B2(n7793), .Y(n4744) );
	o22ai_1 U7499( .A1(n5727), .A2(n7794), .B1(n7793), .B2(n7795), .Y(n4743) );
	o22ai_1 U7500( .A1(n7796), .A2(n7797), .B1(n7793), .B2(n7798), .Y(n4742) );
	nand3_1 U7501( .A(n7590), .B(n7747), .C(n7799), .Y(n7793) );
	inv_1 U7502( .A(n7638), .Y(n7796) );
	o22ai_1 U7503( .A1(n5556), .A2(n7791), .B1(n7800), .B2(n7792), .Y(n4741) );
	o22ai_1 U7504( .A1(n5346), .A2(n7794), .B1(n7800), .B2(n7795), .Y(n4740) );
	o22ai_1 U7505( .A1(n7800), .A2(n7798), .B1(n7801), .B2(n7797), .Y(n4739) );
	inv_1 U7506( .A(n7663), .Y(n7801) );
	mux2i_1 U7507( .A0(n7802), .A1(n7803), .S(n5999), .Y(n7800) );
	nor2_1 U7508( .A(n7804), .B(n7805), .Y(n7802) );
	mux2_1 U7509( .A0(n7806), .A1(n7807), .S(n7808), .X(n7804) );
	o22ai_1 U7510( .A1(n5555), .A2(n7791), .B1(n7809), .B2(n7792), .Y(n4738) );
	o22ai_1 U7511( .A1(n5345), .A2(n7794), .B1(n7809), .B2(n7795), .Y(n4737) );
	o22ai_1 U7512( .A1(n7809), .A2(n7798), .B1(n7810), .B2(n7797), .Y(n4736) );
	inv_1 U7513( .A(n7662), .Y(n7810) );
	mux2i_1 U7514( .A0(n7811), .A1(n7812), .S(n5999), .Y(n7809) );
	nor2_1 U7515( .A(n7813), .B(n7814), .Y(n7811) );
	inv_1 U7516( .A(n7807), .Y(n7814) );
	a222oi_1 U7517( .A1(n7815), .A2(n7816), .B1(n7817), .B2(n7818), .C1(n7819), .C2(n7820), .Y(n7807) );
	o22ai_1 U7518( .A1(n7815), .A2(n7821), .B1(n7822), .B2(n7823), .Y(n7820) );
	o22ai_1 U7519( .A1(n7824), .A2(n7825), .B1(n7826), .B2(n7815), .Y(n7818) );
	a21oi_1 U7520( .A1(n7827), .A2(n7828), .B1(n7829), .Y(n7826) );
	o22ai_1 U7521( .A1(n7830), .A2(n7831), .B1(n7832), .B2(n7833), .Y(n7827) );
	o32ai_1 U7522( .A1(n7819), .A2(n7834), .A3(n7832), .B1(n7835), .B2(n7817), .Y(n7816) );
	a21oi_1 U7523( .A1(n7836), .A2(n7832), .B1(n7837), .Y(n7835) );
	mux2i_1 U7524( .A0(n7830), .A1(n7838), .S(n7828), .Y(n7837) );
	or2_0 U7525( .A(n7825), .B(n7831), .X(n7838) );
	mux2i_1 U7526( .A0(n7805), .A1(n7808), .S(n7806), .Y(n7813) );
	inv_1 U7527( .A(n7839), .Y(n7808) );
	nand2_1 U7528( .A(n7840), .B(n7841), .Y(n7805) );
	nand3_1 U7529( .A(n7831), .B(n7842), .C(n7843), .Y(n7841) );
	inv_1 U7530( .A(n7824), .Y(n7831) );
	mux2i_1 U7531( .A0(n7844), .A1(n7845), .S(n7815), .Y(n7840) );
	o221ai_1 U7532( .A1(n7846), .A2(n15057), .B1(n5355), .B2(n15056), .C1(n7847), .Y(n7815) );
	nand2_1 U7533( .A(g1036), .B(g5657), .Y(n7847) );
	o221ai_1 U7534( .A1(n7848), .A2(n7821), .B1(n7819), .B2(n7849), .C1(n7850), .Y(n7845) );
	mux2i_1 U7535( .A0(n7851), .A1(n7852), .S(n7817), .Y(n7850) );
	nor2_1 U7536( .A(n7853), .B(n7828), .Y(n7852) );
	a21oi_1 U7537( .A1(n7834), .A2(n7848), .B1(n7842), .Y(n7853) );
	nor2_1 U7538( .A(n7824), .B(n7854), .Y(n7851) );
	a221oi_1 U7539( .A1(n7855), .A2(n7824), .B1(n7856), .B2(n7842), .C1(n7829), .Y(n7849) );
	inv_1 U7540( .A(n7828), .Y(n7819) );
	o21ai_0 U7541( .A1(n7834), .A2(n7857), .B1(n7858), .Y(n7844) );
	mux2i_1 U7542( .A0(n7859), .A1(n7860), .S(n7828), .Y(n7858) );
	o221ai_1 U7543( .A1(n7846), .A2(n15063), .B1(n5355), .B2(n15061), .C1(n7861), .Y(n7828) );
	nand2_1 U7544( .A(g1051), .B(g5657), .Y(n7861) );
	o22ai_1 U7545( .A1(n7848), .A2(n7825), .B1(n7862), .B2(n7823), .Y(n7860) );
	inv_1 U7546( .A(n7856), .Y(n7823) );
	nor2_1 U7547( .A(n7817), .B(n7832), .Y(n7856) );
	nor3_1 U7548( .A(n7855), .B(n7829), .C(n7843), .Y(n7859) );
	nor2_1 U7549( .A(n7848), .B(n7822), .Y(n7829) );
	a21oi_1 U7550( .A1(n7824), .A2(n7817), .B1(n7832), .Y(n7857) );
	inv_1 U7551( .A(n7848), .Y(n7832) );
	o221ai_1 U7552( .A1(n7846), .A2(n15059), .B1(n5355), .B2(n15058), .C1(n7863), .Y(n7848) );
	nand2_1 U7553( .A(g1066), .B(g5657), .Y(n7863) );
	o221ai_1 U7554( .A1(n7846), .A2(n15055), .B1(n5355), .B2(n15054), .C1(n7864), .Y(n7824) );
	nand2_1 U7555( .A(g5657), .B(g1081), .Y(n7864) );
	o22ai_1 U7556( .A1(n7791), .A2(n5623), .B1(n7792), .B2(n7865), .Y(n4735) );
	o22ai_1 U7557( .A1(n7794), .A2(n5597), .B1(n7795), .B2(n7865), .Y(n4734) );
	o22ai_1 U7558( .A1(n7797), .A2(n5406), .B1(n7798), .B2(n7865), .Y(n4733) );
	nand2_1 U7559( .A(n7806), .B(n5999), .Y(n7865) );
	o211ai_1 U7560( .A1(n7866), .A2(n5406), .B1(n7867), .C1(n7868), .Y(n7806) );
	a22oi_1 U7561( .A1(n9799), .A2(g6944), .B1(n9798), .B2(n7226), .Y(n7868) );
	nand3_1 U7562( .A(n7256), .B(n7869), .C(g1228), .Y(n7867) );
	o22ai_1 U7563( .A1(n7791), .A2(n5624), .B1(n7792), .B2(n7870), .Y(n4732) );
	o22ai_1 U7564( .A1(n7794), .A2(n5598), .B1(n7795), .B2(n7870), .Y(n4731) );
	inv_1 U7565( .A(n153), .Y(n7795) );
	nand2_1 U7566( .A(n7871), .B(n5744), .Y(n7794) );
	o22ai_1 U7567( .A1(n7797), .A2(n5407), .B1(n7798), .B2(n7870), .Y(n4730) );
	nand2_1 U7568( .A(n7839), .B(n5999), .Y(n7870) );
	o211ai_1 U7569( .A1(n7866), .A2(n5407), .B1(n7872), .C1(n7873), .Y(n7839) );
	a22oi_1 U7570( .A1(n9801), .A2(g6944), .B1(n9800), .B2(n7226), .Y(n7873) );
	nand3_1 U7571( .A(n7256), .B(n7874), .C(g1210), .Y(n7872) );
	inv_1 U7572( .A(n152), .Y(n7798) );
	nand2_1 U7573( .A(n5756), .B(n7866), .Y(n7797) );
	o22ai_1 U7574( .A1(n7875), .A2(n7876), .B1(n7877), .B2(n7878), .Y(n4729) );
	inv_1 U7575( .A(n7365), .Y(n7878) );
	o22ai_1 U7576( .A1(n7875), .A2(n7879), .B1(n7880), .B2(n7881), .Y(n4728) );
	inv_1 U7577( .A(n7366), .Y(n7881) );
	o22ai_1 U7578( .A1(n7875), .A2(n7882), .B1(n7883), .B2(n5512), .Y(n4727) );
	o21ai_0 U7579( .A1(n7825), .A2(n7884), .B1(n5760), .Y(n7875) );
	nand2_1 U7580( .A(n7822), .B(n7830), .Y(n7825) );
	o22ai_1 U7581( .A1(n7876), .A2(n7885), .B1(n7877), .B2(n7886), .Y(n4726) );
	inv_1 U7582( .A(n7359), .Y(n7886) );
	o22ai_1 U7583( .A1(n7879), .A2(n7885), .B1(n7880), .B2(n7887), .Y(n4725) );
	inv_1 U7584( .A(n7360), .Y(n7887) );
	o22ai_1 U7585( .A1(n7882), .A2(n7885), .B1(n7883), .B2(n5511), .Y(n4724) );
	o221ai_1 U7586( .A1(n7822), .A2(n7888), .B1(n7889), .B2(n7833), .C1(n5747), .Y(n7885) );
	inv_1 U7587( .A(n7836), .Y(n7833) );
	nor2_1 U7588( .A(n7854), .B(n7862), .Y(n7836) );
	mux2i_1 U7589( .A0(n5984), .A1(n5983), .S(n7817), .Y(n7888) );
	o22ai_1 U7590( .A1(n7876), .A2(n7890), .B1(n7877), .B2(n7891), .Y(n4723) );
	inv_1 U7591( .A(n7361), .Y(n7891) );
	o22ai_1 U7592( .A1(n7879), .A2(n7890), .B1(n7880), .B2(n7892), .Y(n4722) );
	inv_1 U7593( .A(n7362), .Y(n7892) );
	o22ai_1 U7594( .A1(n7882), .A2(n7890), .B1(n7883), .B2(n5510), .Y(n4721) );
	o211ai_1 U7595( .A1(n7830), .A2(n7889), .B1(n7821), .C1(n5740), .Y(n7890) );
	inv_1 U7596( .A(n7884), .Y(n7889) );
	xnor2_1 U7597( .A(n7843), .B(n5983), .Y(n7884) );
	inv_1 U7598( .A(n7817), .Y(n7843) );
	o22ai_1 U7599( .A1(n7876), .A2(n7893), .B1(n7877), .B2(n7894), .Y(n4720) );
	inv_1 U7600( .A(n7363), .Y(n7894) );
	nand2_1 U7601( .A(n7876), .B(n5744), .Y(n7877) );
	nand2_1 U7602( .A(n7226), .B(n7790), .Y(n7876) );
	o22ai_1 U7603( .A1(n7879), .A2(n7893), .B1(n7880), .B2(n7895), .Y(n4719) );
	inv_1 U7604( .A(n7364), .Y(n7895) );
	nand2_1 U7605( .A(n7879), .B(n5744), .Y(n7880) );
	nand2_1 U7606( .A(g6944), .B(n7790), .Y(n7879) );
	o22ai_1 U7607( .A1(n7882), .A2(n7893), .B1(n7883), .B2(n5509), .Y(n4718) );
	nand2_1 U7608( .A(n7882), .B(n5747), .Y(n7883) );
	o221ai_1 U7609( .A1(n6098), .A2(n7834), .B1(g3229), .B2(n7821), .C1(n7896), .Y(n7893) );
	a21oi_1 U7610( .A1(n7897), .A2(n7817), .B1(RST), .Y(n7896) );
	o221ai_1 U7611( .A1(n7364), .A2(n7871), .B1(n7363), .B2(n7898), .C1(n7899), .Y(n7817) );
	nand2_1 U7612( .A(g6750), .B(n5509), .Y(n7899) );
	o22ai_1 U7613( .A1(n7830), .A2(n5983), .B1(n7900), .B2(n7854), .Y(n7897) );
	nor2_1 U7614( .A(n7822), .B(n5983), .Y(n7900) );
	inv_1 U7615( .A(n7842), .Y(n7830) );
	inv_1 U7616( .A(n7855), .Y(n7821) );
	nor2_1 U7617( .A(n7842), .B(n7822), .Y(n7855) );
	inv_1 U7618( .A(n7862), .Y(n7822) );
	o221ai_1 U7619( .A1(n7362), .A2(n7871), .B1(n7361), .B2(n7898), .C1(n7901), .Y(n7862) );
	nand2_1 U7620( .A(g6750), .B(n5510), .Y(n7901) );
	o221ai_1 U7621( .A1(n7360), .A2(n7871), .B1(n7359), .B2(n7898), .C1(n7902), .Y(n7842) );
	nand2_1 U7622( .A(g6750), .B(n5511), .Y(n7902) );
	inv_1 U7623( .A(n7854), .Y(n7834) );
	o221ai_1 U7624( .A1(n7366), .A2(n7871), .B1(n7365), .B2(n7898), .C1(n7903), .Y(n7854) );
	nand2_1 U7625( .A(g6750), .B(n5512), .Y(n7903) );
	nand2_1 U7626( .A(g6750), .B(n7790), .Y(n7882) );
	o32ai_1 U7627( .A1(n7904), .A2(n7747), .A3(n7788), .B1(n6755), .B2(n7905), .Y(n7790) );
	nor2_1 U7628( .A(n7799), .B(n7219), .Y(n7905) );
	inv_1 U7629( .A(n7803), .Y(n7219) );
	inv_1 U7630( .A(n7904), .Y(n7799) );
	inv_1 U7631( .A(n7812), .Y(n7747) );
	o21ai_0 U7632( .A1(n7898), .A2(n5564), .B1(n7906), .Y(n7904) );
	a22oi_1 U7633( .A1(n7638), .A2(g6750), .B1(n9802), .B2(g6944), .Y(n7906) );
	and2_0 U7634( .A(g1244), .B(n5758), .X(n4717) );
	and2_0 U7635( .A(g1229), .B(n5758), .X(n4716) );
	o22ai_1 U7636( .A1(n7907), .A2(n7908), .B1(n7909), .B2(n5653), .Y(n4715) );
	o22ai_1 U7637( .A1(n7907), .A2(n7910), .B1(n7911), .B2(n7912), .Y(n4714) );
	inv_1 U7638( .A(n7461), .Y(n7912) );
	o22ai_1 U7639( .A1(n7907), .A2(n7913), .B1(n7914), .B2(n5422), .Y(n4713) );
	o22ai_1 U7640( .A1(n7908), .A2(n7915), .B1(n7909), .B2(n5654), .Y(n4712) );
	o22ai_1 U7641( .A1(n7910), .A2(n7915), .B1(n7911), .B2(n7916), .Y(n4711) );
	inv_1 U7642( .A(n7457), .Y(n7916) );
	o22ai_1 U7643( .A1(n7913), .A2(n7915), .B1(n7914), .B2(n5423), .Y(n4710) );
	o22ai_1 U7644( .A1(n7917), .A2(n7908), .B1(n7909), .B2(n5655), .Y(n4709) );
	or2_0 U7645( .A(RST), .B(n7258), .X(n7909) );
	o22ai_1 U7646( .A1(n7917), .A2(n7910), .B1(n7911), .B2(n7918), .Y(n4708) );
	inv_1 U7647( .A(n7454), .Y(n7918) );
	or2_0 U7648( .A(RST), .B(g8007), .X(n7911) );
	o22ai_1 U7649( .A1(n7917), .A2(n7913), .B1(n7914), .B2(n5421), .Y(n4707) );
	or2_0 U7650( .A(RST), .B(g7961), .X(n7914) );
	and2_0 U7651( .A(g1254), .B(n5758), .X(n4706) );
	and2_0 U7652( .A(g1260), .B(n5758), .X(n4705) );
	and2_0 U7653( .A(g1258), .B(n5759), .X(n4704) );
	and2_0 U7654( .A(g1250), .B(n5758), .X(n4703) );
	o22ai_1 U7655( .A1(n7788), .A2(n7791), .B1(n7792), .B2(n7919), .Y(n4702) );
	o22ai_1 U7656( .A1(n7791), .A2(n7919), .B1(n9972), .B2(n7792), .Y(n4701) );
	o22ai_1 U7657( .A1(n7791), .A2(n5591), .B1(n6118), .B2(n7792), .Y(n4700) );
	nand2_1 U7658( .A(n7226), .B(n5747), .Y(n7792) );
	nand2_1 U7659( .A(n7898), .B(n5748), .Y(n7791) );
	nor2_1 U7660( .A(RST), .B(n7846), .Y(n4699) );
	inv_1 U7661( .A(g5686), .Y(n7846) );
	and2_0 U7662( .A(g1084), .B(n5759), .X(n4698) );
	and2_0 U7663( .A(g1082), .B(n5758), .X(n4697) );
	and2_0 U7664( .A(g1069), .B(n5758), .X(n4696) );
	and2_0 U7665( .A(g1067), .B(n5758), .X(n4695) );
	and2_0 U7666( .A(g1054), .B(n5759), .X(n4694) );
	and2_0 U7667( .A(g1052), .B(n5741), .X(n4693) );
	and2_0 U7668( .A(g1039), .B(n5758), .X(n4692) );
	and2_0 U7669( .A(g1037), .B(n5759), .X(n4691) );
	and2_0 U7670( .A(n5760), .B(n6773), .X(n4690) );
	mux2i_1 U7671( .A0(g985), .A1(n7920), .S(n7742), .Y(n6773) );
	mux2_1 U7672( .A0(n5568), .A1(n7921), .S(g6712), .X(n7920) );
	nor2_1 U7673( .A(RST), .B(n7922), .Y(n4689) );
	and2_0 U7674( .A(g977), .B(n5759), .X(n4688) );
	o22ai_1 U7675( .A1(n7923), .A2(n7924), .B1(n7925), .B2(n7926), .Y(n4687) );
	o21ai_0 U7676( .A1(n7927), .A2(n7928), .B1(n5764), .Y(n7926) );
	inv_1 U7677( .A(n7378), .Y(n7925) );
	o22ai_1 U7678( .A1(n7924), .A2(n7929), .B1(n7930), .B2(n7931), .Y(n4686) );
	o21ai_0 U7679( .A1(n7932), .A2(n7928), .B1(n5761), .Y(n7931) );
	o22ai_1 U7680( .A1(n7924), .A2(n7933), .B1(n7934), .B2(n7935), .Y(n4685) );
	inv_1 U7681( .A(n7377), .Y(n7935) );
	a21oi_1 U7682( .A1(n7928), .A2(n5755), .B1(n7936), .Y(n7934) );
	nand2_1 U7683( .A(n7263), .B(n7928), .Y(n7924) );
	nand3_1 U7684( .A(n7937), .B(n7938), .C(n7263), .Y(n7928) );
	inv_1 U7685( .A(n7939), .Y(n7938) );
	o22ai_1 U7686( .A1(n7923), .A2(n7940), .B1(n7941), .B2(n7942), .Y(n4684) );
	nor2_1 U7687( .A(n7943), .B(n7944), .Y(n7941) );
	o22ai_1 U7688( .A1(n7929), .A2(n7940), .B1(n7945), .B2(n7946), .Y(n4683) );
	inv_1 U7689( .A(n7728), .Y(n7946) );
	nor2_1 U7690( .A(n7943), .B(n7947), .Y(n7945) );
	o22ai_1 U7691( .A1(n7933), .A2(n7940), .B1(n7948), .B2(n7949), .Y(n4682) );
	nor2_1 U7692( .A(n7943), .B(n7936), .Y(n7948) );
	and2_0 U7693( .A(n7950), .B(n5765), .X(n7943) );
	nand2_1 U7694( .A(n7951), .B(n7950), .Y(n7940) );
	nand2_1 U7695( .A(n7937), .B(n7952), .Y(n7950) );
	o21ai_0 U7696( .A1(n7915), .A2(n7953), .B1(n7954), .Y(n7952) );
	nand4_1 U7697( .A(n7955), .B(n7956), .C(n7957), .D(n7958), .Y(n7954) );
	mux2i_1 U7698( .A0(n7953), .A1(n7959), .S(n7915), .Y(n7951) );
	o22ai_1 U7699( .A1(n7923), .A2(n7960), .B1(n7961), .B2(n7962), .Y(n4681) );
	o22ai_1 U7700( .A1(n7929), .A2(n7960), .B1(n7963), .B2(n5663), .Y(n4680) );
	o22ai_1 U7701( .A1(n7964), .A2(n7965), .B1(n7933), .B2(n7960), .Y(n4679) );
	nand2_1 U7702( .A(n7966), .B(n7967), .Y(n7960) );
	mux2i_1 U7703( .A0(n7968), .A1(n7969), .S(n7970), .Y(n7966) );
	nand2_1 U7704( .A(n7958), .B(n7969), .Y(n7968) );
	o211ai_1 U7705( .A1(n7955), .A2(n7971), .B1(n7958), .C1(n7972), .Y(n7969) );
	mux2i_1 U7706( .A0(n7973), .A1(n7974), .S(n7975), .Y(n7972) );
	a21oi_1 U7707( .A1(n7976), .A2(n7977), .B1(n7978), .Y(n7974) );
	nand2_1 U7708( .A(n7955), .B(n7957), .Y(n7977) );
	nand3_1 U7709( .A(n7263), .B(n7956), .C(n7955), .Y(n7973) );
	inv_1 U7710( .A(n7959), .Y(n7971) );
	nand2_1 U7711( .A(n7976), .B(n7957), .Y(n7959) );
	inv_1 U7712( .A(n7465), .Y(n7965) );
	o22ai_1 U7713( .A1(n7923), .A2(n7979), .B1(n7961), .B2(n7980), .Y(n4678) );
	o22ai_1 U7714( .A1(n7929), .A2(n7979), .B1(n7963), .B2(n5664), .Y(n4677) );
	o22ai_1 U7715( .A1(n7964), .A2(n7981), .B1(n7933), .B2(n7979), .Y(n4676) );
	nand2_1 U7716( .A(n7982), .B(n7967), .Y(n7979) );
	xnor2_1 U7717( .A(n7983), .B(n7984), .Y(n7982) );
	a21oi_1 U7718( .A1(n7985), .A2(n7958), .B1(n7986), .Y(n7984) );
	o22ai_1 U7719( .A1(n7987), .A2(n7988), .B1(n7989), .B2(n7975), .Y(n7985) );
	a21oi_1 U7720( .A1(n7990), .A2(n7937), .B1(n7978), .Y(n7989) );
	a21oi_1 U7721( .A1(n7991), .A2(n7955), .B1(n7992), .Y(n7990) );
	mux2i_1 U7722( .A0(n7993), .A1(n7994), .S(n7975), .Y(n7988) );
	o21ai_0 U7723( .A1(n7970), .A2(n7995), .B1(n7996), .Y(n7994) );
	and2_0 U7724( .A(n7995), .B(n7955), .X(n7993) );
	nand2_1 U7725( .A(n7997), .B(n7957), .Y(n7995) );
	nand4_1 U7726( .A(n7998), .B(n7999), .C(n8000), .D(n8001), .Y(n7957) );
	nor3_1 U7727( .A(n8002), .B(n8003), .C(n8004), .Y(n8001) );
	nand3_1 U7728( .A(n8005), .B(n8006), .C(n8007), .Y(n8002) );
	nor3_1 U7729( .A(n8008), .B(n8009), .C(n8010), .Y(n8000) );
	inv_1 U7730( .A(n7467), .Y(n7981) );
	o22ai_1 U7731( .A1(n7923), .A2(n8011), .B1(n7961), .B2(n8012), .Y(n4675) );
	o22ai_1 U7732( .A1(n7929), .A2(n8011), .B1(n7963), .B2(n5665), .Y(n4674) );
	o22ai_1 U7733( .A1(n7964), .A2(n8013), .B1(n7933), .B2(n8011), .Y(n4673) );
	o21ai_0 U7734( .A1(n8014), .A2(n8015), .B1(n7967), .Y(n8011) );
	nor3_1 U7735( .A(n7956), .B(n8016), .C(n8017), .Y(n8015) );
	inv_1 U7736( .A(n7463), .Y(n8013) );
	o22ai_1 U7737( .A1(n7923), .A2(n8018), .B1(n8019), .B2(n8020), .Y(n4672) );
	o21ai_0 U7738( .A1(n7927), .A2(n8021), .B1(n5763), .Y(n8020) );
	inv_1 U7739( .A(n7583), .Y(n8019) );
	o22ai_1 U7740( .A1(n7929), .A2(n8018), .B1(n8022), .B2(n8023), .Y(n4671) );
	o21ai_0 U7741( .A1(n7932), .A2(n8021), .B1(n5746), .Y(n8023) );
	nand2_1 U7742( .A(n8024), .B(n8025), .Y(n8021) );
	inv_1 U7743( .A(n8026), .Y(n8024) );
	inv_1 U7744( .A(n7584), .Y(n8022) );
	o32ai_1 U7745( .A1(n8027), .A2(RST), .A3(n8028), .B1(n7933), .B2(n8018), .Y(n4670) );
	o211ai_1 U7746( .A1(n7917), .A2(n8029), .B1(n7263), .C1(n8030), .Y(n8018) );
	mux2i_1 U7747( .A0(n7917), .A1(n8029), .S(n8031), .Y(n8030) );
	nor3_1 U7748( .A(n8026), .B(n8032), .C(n8033), .Y(n8028) );
	o22ai_1 U7749( .A1(n7923), .A2(n8034), .B1(n5332), .B2(n7961), .Y(n4669) );
	o22ai_1 U7750( .A1(n7929), .A2(n8034), .B1(n8035), .B2(n7963), .Y(n4668) );
	inv_1 U7751( .A(n7634), .Y(n8035) );
	o22ai_1 U7752( .A1(n5524), .A2(n7964), .B1(n7933), .B2(n8034), .Y(n4667) );
	xnor2_1 U7753( .A(n8036), .B(n7917), .Y(n8034) );
	inv_1 U7754( .A(n8037), .Y(n7917) );
	or2_0 U7755( .A(n8026), .B(n8025), .X(n8036) );
	a21oi_1 U7756( .A1(n8027), .A2(g5472), .B1(n8033), .Y(n8025) );
	o22ai_1 U7757( .A1(n7583), .A2(n7927), .B1(n7584), .B2(n7932), .Y(n8033) );
	inv_1 U7758( .A(n7736), .Y(n8027) );
	nand2_1 U7759( .A(n8038), .B(n7263), .Y(n8026) );
	mux2i_1 U7760( .A0(n8039), .A1(n8040), .S(n8031), .Y(n8038) );
	nand2_1 U7761( .A(n8029), .B(n8037), .Y(n8040) );
	or2_0 U7762( .A(n8037), .B(n8029), .X(n8039) );
	o221ai_1 U7763( .A1(n8032), .A2(n5524), .B1(n7927), .B2(n5332), .C1(n8041), .Y(n8037) );
	nand2_1 U7764( .A(n7634), .B(g6712), .Y(n8041) );
	o22ai_1 U7765( .A1(n7923), .A2(n8042), .B1(n7961), .B2(n5670), .Y(n4666) );
	o22ai_1 U7766( .A1(n7929), .A2(n8042), .B1(n7963), .B2(n8043), .Y(n4665) );
	o22ai_1 U7767( .A1(n7964), .A2(n5633), .B1(n7933), .B2(n8042), .Y(n4664) );
	mux2_1 U7768( .A0(n8031), .A1(n8029), .S(n7263), .X(n8042) );
	o21ai_0 U7769( .A1(n8044), .A2(n8045), .B1(n8046), .Y(n8029) );
	inv_1 U7770( .A(n8047), .Y(n8046) );
	o22ai_1 U7771( .A1(n9973), .A2(n8048), .B1(n7387), .B2(n8049), .Y(n8045) );
	nor2_1 U7772( .A(n7389), .B(n8050), .Y(n8044) );
	a221oi_1 U7773( .A1(g5472), .A2(n9808), .B1(n7775), .B2(n10002), .C1(n8051), .Y(n8031) );
	nor2_1 U7774( .A(n8043), .B(n7932), .Y(n8051) );
	inv_1 U7775( .A(n7630), .Y(n8043) );
	o22ai_1 U7776( .A1(n7923), .A2(n8052), .B1(n8053), .B2(n8054), .Y(n4663) );
	nor2_1 U7777( .A(n8055), .B(n7944), .Y(n8053) );
	o22ai_1 U7778( .A1(n7929), .A2(n8052), .B1(n8056), .B2(n8057), .Y(n4662) );
	nor2_1 U7779( .A(n8055), .B(n7947), .Y(n8056) );
	o22ai_1 U7780( .A1(n7933), .A2(n8052), .B1(n8058), .B2(n8059), .Y(n4661) );
	inv_1 U7781( .A(n7339), .Y(n8059) );
	nor2_1 U7782( .A(n8055), .B(n7936), .Y(n8058) );
	a21oi_1 U7783( .A1(n8060), .A2(n8061), .B1(RST), .Y(n8055) );
	o22ai_1 U7784( .A1(n8062), .A2(n7923), .B1(n5333), .B2(n7961), .Y(n4660) );
	o22ai_1 U7785( .A1(n8062), .A2(n7929), .B1(n8063), .B2(n7963), .Y(n4659) );
	inv_1 U7786( .A(n7620), .Y(n8063) );
	o22ai_1 U7787( .A1(n5525), .A2(n7964), .B1(n8062), .B2(n7933), .Y(n4658) );
	xnor2_1 U7788( .A(n7922), .B(n8064), .Y(n8062) );
	a21oi_1 U7789( .A1(n7978), .A2(n8065), .B1(n8066), .Y(n8064) );
	nor4_1 U7790( .A(n8061), .B(n8067), .C(n7953), .D(n8068), .Y(n8066) );
	inv_1 U7791( .A(n8069), .Y(n8061) );
	o22ai_1 U7792( .A1(n8070), .A2(n7923), .B1(n7961), .B2(n5671), .Y(n4657) );
	inv_1 U7793( .A(n7944), .Y(n7961) );
	nor2_1 U7794( .A(RST), .B(n7775), .Y(n7944) );
	nand2_1 U7795( .A(n7775), .B(n5753), .Y(n7923) );
	o22ai_1 U7796( .A1(n8070), .A2(n7929), .B1(n7963), .B2(n8071), .Y(n4656) );
	inv_1 U7797( .A(n7947), .Y(n7963) );
	nor2_1 U7798( .A(RST), .B(g6712), .Y(n7947) );
	inv_1 U7799( .A(n3961), .Y(n7929) );
	o22ai_1 U7800( .A1(n8070), .A2(n7933), .B1(n7964), .B2(n5672), .Y(n4655) );
	inv_1 U7801( .A(n7936), .Y(n7964) );
	nor2_1 U7802( .A(g5472), .B(RST), .Y(n7936) );
	inv_1 U7803( .A(n138), .Y(n7933) );
	xnor2_1 U7804( .A(n8067), .B(n8072), .Y(n8070) );
	a21oi_1 U7805( .A1(n8073), .A2(n7263), .B1(n8074), .Y(n8072) );
	inv_1 U7806( .A(n8052), .Y(n8074) );
	nand2_1 U7807( .A(n8067), .B(n8060), .Y(n8052) );
	o32ai_1 U7808( .A1(n7953), .A2(n7922), .A3(n8075), .B1(n7978), .B2(n8076), .Y(n8060) );
	inv_1 U7809( .A(n8065), .Y(n8076) );
	nor3_1 U7810( .A(n7953), .B(n7907), .C(n8077), .Y(n8065) );
	inv_1 U7811( .A(n8075), .Y(n8077) );
	inv_1 U7812( .A(n7263), .Y(n7953) );
	a21oi_1 U7813( .A1(n8078), .A2(n8079), .B1(n8067), .Y(n8073) );
	inv_1 U7814( .A(n8068), .Y(n8079) );
	xnor2_1 U7815( .A(n8075), .B(n7907), .Y(n8068) );
	nor3_1 U7816( .A(n8080), .B(n8081), .C(n8047), .Y(n8075) );
	a21oi_1 U7817( .A1(n7978), .A2(n7922), .B1(n8069), .Y(n8078) );
	o21ai_0 U7818( .A1(n7339), .A2(n8032), .B1(n8082), .Y(n8069) );
	a22oi_1 U7819( .A1(g6712), .A2(n8057), .B1(n7775), .B2(n8054), .Y(n8082) );
	inv_1 U7820( .A(n7340), .Y(n8054) );
	inv_1 U7821( .A(n7734), .Y(n8057) );
	inv_1 U7822( .A(n7907), .Y(n7922) );
	o221ai_1 U7823( .A1(n8032), .A2(n5525), .B1(n7927), .B2(n5333), .C1(n8083), .Y(n7907) );
	nand2_1 U7824( .A(n7620), .B(g6712), .Y(n8083) );
	a221oi_1 U7825( .A1(g5472), .A2(n9809), .B1(n7775), .B2(n10003), .C1(n8084), .Y(n8067) );
	nor2_1 U7826( .A(n8071), .B(n7932), .Y(n8084) );
	inv_1 U7827( .A(n7626), .Y(n8071) );
	and2_0 U7828( .A(g5595), .B(n5765), .X(n4654) );
	nor2_1 U7829( .A(n8085), .B(n8086), .Y(n4653) );
	xnor2_1 U7830( .A(n10004), .B(n8087), .Y(n8085) );
	nor2_1 U7831( .A(n8088), .B(n8089), .Y(n8087) );
	nor2_1 U7832( .A(n8090), .B(n8086), .Y(n4652) );
	xnor2_1 U7833( .A(n8088), .B(n8089), .Y(n8090) );
	inv_1 U7834( .A(n7305), .Y(n8089) );
	nand2_1 U7835( .A(n7707), .B(n8091), .Y(n8088) );
	nor2_1 U7836( .A(n8092), .B(n8086), .Y(n4651) );
	xnor2_1 U7837( .A(n7707), .B(n8091), .Y(n8092) );
	a211oi_1 U7838( .A1(n5378), .A2(n8093), .B1(n8086), .C1(n8091), .Y(n4650) );
	nor2_1 U7839( .A(n5378), .B(n8093), .Y(n8091) );
	nor3_1 U7840( .A(n8086), .B(n8094), .C(n8095), .Y(n4649) );
	a21oi_1 U7841( .A1(n10006), .A2(n8096), .B1(n7698), .Y(n8095) );
	inv_1 U7842( .A(n8093), .Y(n8094) );
	nand3_1 U7843( .A(n7698), .B(n8096), .C(n10006), .Y(n8093) );
	nor2_1 U7844( .A(n8097), .B(n8086), .Y(n4648) );
	xnor2_1 U7845( .A(n10006), .B(n8096), .Y(n8097) );
	a211oi_1 U7846( .A1(n8098), .A2(n8099), .B1(n8086), .C1(n8096), .Y(n4647) );
	nor2_1 U7847( .A(n8098), .B(n8099), .Y(n8096) );
	inv_1 U7848( .A(n7711), .Y(n8098) );
	inv_1 U7849( .A(n8100), .Y(n4646) );
	o211ai_1 U7850( .A1(n10007), .A2(n8101), .B1(n8102), .C1(n8099), .Y(n8100) );
	nand2_1 U7851( .A(n10007), .B(n8101), .Y(n8099) );
	inv_1 U7852( .A(n8086), .Y(n8102) );
	nor3_1 U7853( .A(n8086), .B(n8101), .C(n8103), .Y(n4645) );
	a21oi_1 U7854( .A1(n10001), .A2(n8104), .B1(n7701), .Y(n8103) );
	and3_1 U7855( .A(n7701), .B(n8104), .C(n10001), .X(n8101) );
	nor2_1 U7856( .A(n8105), .B(n8086), .Y(n4644) );
	o21ai_0 U7857( .A1(n6131), .A2(n8106), .B1(n5754), .Y(n8086) );
	xnor2_1 U7858( .A(n8104), .B(n10001), .Y(n8105) );
	nor2_1 U7859( .A(n8048), .B(n6337), .Y(n8104) );
	o22ai_1 U7860( .A1(n8107), .A2(n8108), .B1(n8109), .B2(n8110), .Y(n4643) );
	o22ai_1 U7861( .A1(n5728), .A2(n8111), .B1(n8109), .B2(n8112), .Y(n4642) );
	o22ai_1 U7862( .A1(n5685), .A2(n8113), .B1(n8109), .B2(n8114), .Y(n4641) );
	o221ai_1 U7863( .A1(n8115), .A2(n8116), .B1(n8117), .B2(n8118), .C1(n8119), .Y(n8109) );
	xnor2_1 U7864( .A(n8120), .B(n8121), .Y(n8115) );
	nor2_1 U7865( .A(n8122), .B(n8123), .Y(n8121) );
	xnor2_1 U7866( .A(n8124), .B(n8014), .Y(n8122) );
	o22ai_1 U7867( .A1(n8125), .A2(n8108), .B1(n8126), .B2(n8110), .Y(n4640) );
	o22ai_1 U7868( .A1(n5537), .A2(n8111), .B1(n8126), .B2(n8112), .Y(n4639) );
	o22ai_1 U7869( .A1(n5705), .A2(n8113), .B1(n8126), .B2(n8114), .Y(n4638) );
	inv_1 U7870( .A(n8127), .Y(n8126) );
	o221ai_1 U7871( .A1(n8081), .A2(n8118), .B1(n8014), .B2(n8128), .C1(n8129), .Y(n8127) );
	nand2_1 U7872( .A(n8130), .B(n8131), .Y(n8129) );
	inv_1 U7873( .A(n8116), .Y(n8131) );
	xnor2_1 U7874( .A(n8123), .B(n8132), .Y(n8130) );
	o211ai_1 U7875( .A1(n8133), .A2(n8134), .B1(n8135), .C1(n8136), .Y(n8123) );
	mux2i_1 U7876( .A0(n8133), .A1(n8134), .S(n8137), .Y(n8136) );
	o22ai_1 U7877( .A1(n8138), .A2(n8108), .B1(n8139), .B2(n8110), .Y(n4637) );
	o22ai_1 U7878( .A1(n5536), .A2(n8111), .B1(n8139), .B2(n8112), .Y(n4636) );
	o22ai_1 U7879( .A1(n5706), .A2(n8113), .B1(n8139), .B2(n8114), .Y(n4635) );
	inv_1 U7880( .A(n8140), .Y(n8139) );
	o22ai_1 U7881( .A1(n8141), .A2(n8118), .B1(n8116), .B2(n8142), .Y(n8140) );
	xor2_1 U7882( .A(n8134), .B(n8143), .X(n8142) );
	nand2_1 U7883( .A(n8144), .B(n8135), .Y(n8143) );
	inv_1 U7884( .A(n8145), .Y(n8135) );
	xnor2_1 U7885( .A(n8133), .B(n8137), .Y(n8144) );
	o22ai_1 U7886( .A1(n8146), .A2(n8108), .B1(n8147), .B2(n8110), .Y(n4634) );
	o22ai_1 U7887( .A1(n5540), .A2(n8111), .B1(n8147), .B2(n8112), .Y(n4633) );
	o22ai_1 U7888( .A1(n5707), .A2(n8113), .B1(n8147), .B2(n8114), .Y(n4632) );
	inv_1 U7889( .A(n8148), .Y(n8147) );
	o22ai_1 U7890( .A1(n8149), .A2(n8118), .B1(n8116), .B2(n8150), .Y(n8148) );
	xnor2_1 U7891( .A(n8133), .B(n8145), .Y(n8150) );
	mux2i_1 U7892( .A0(n8151), .A1(n8152), .S(n8153), .Y(n8145) );
	o22ai_1 U7893( .A1(n8154), .A2(n8108), .B1(n8155), .B2(n8110), .Y(n4631) );
	o22ai_1 U7894( .A1(n5729), .A2(n8111), .B1(n8155), .B2(n8112), .Y(n4630) );
	o22ai_1 U7895( .A1(n5686), .A2(n8113), .B1(n8155), .B2(n8114), .Y(n4629) );
	inv_1 U7896( .A(n8156), .Y(n8155) );
	o22ai_1 U7897( .A1(n8157), .A2(n8118), .B1(n8158), .B2(n8116), .Y(n8156) );
	xnor2_1 U7898( .A(n8159), .B(n8160), .Y(n8158) );
	nor2_1 U7899( .A(n8152), .B(n8151), .Y(n8160) );
	nor3_1 U7900( .A(n8161), .B(n8014), .C(n8162), .Y(n8151) );
	nor3_1 U7901( .A(n8137), .B(n8163), .C(n8162), .Y(n8152) );
	o22ai_1 U7902( .A1(n8164), .A2(n8108), .B1(n8165), .B2(n8110), .Y(n4628) );
	o22ai_1 U7903( .A1(n5541), .A2(n8111), .B1(n8165), .B2(n8112), .Y(n4627) );
	o22ai_1 U7904( .A1(n5708), .A2(n8113), .B1(n8165), .B2(n8114), .Y(n4626) );
	inv_1 U7905( .A(n8166), .Y(n8165) );
	o22ai_1 U7906( .A1(n8167), .A2(n8118), .B1(n8116), .B2(n8168), .Y(n8166) );
	xnor2_1 U7907( .A(n8162), .B(n8163), .Y(n8168) );
	nand2_1 U7908( .A(n8169), .B(n8170), .Y(n8162) );
	xnor2_1 U7909( .A(n8171), .B(n8137), .Y(n8170) );
	o22ai_1 U7910( .A1(n8172), .A2(n8108), .B1(n8110), .B2(n8173), .Y(n4625) );
	o22ai_1 U7911( .A1(n5535), .A2(n8111), .B1(n8112), .B2(n8173), .Y(n4624) );
	o22ai_1 U7912( .A1(n5709), .A2(n8113), .B1(n8114), .B2(n8173), .Y(n4623) );
	o221ai_1 U7913( .A1(n8174), .A2(n8116), .B1(n7248), .B2(n8118), .C1(n8119), .Y(n8173) );
	xnor2_1 U7914( .A(n8171), .B(n8169), .Y(n8174) );
	nor2_1 U7915( .A(n8175), .B(n8176), .Y(n8169) );
	xnor2_1 U7916( .A(n8177), .B(n8137), .Y(n8176) );
	o22ai_1 U7917( .A1(n8178), .A2(n8108), .B1(n8179), .B2(n8110), .Y(n4622) );
	o22ai_1 U7918( .A1(n5539), .A2(n8111), .B1(n8179), .B2(n8112), .Y(n4621) );
	o22ai_1 U7919( .A1(n5710), .A2(n8113), .B1(n8179), .B2(n8114), .Y(n4620) );
	inv_1 U7920( .A(n8180), .Y(n8179) );
	o221ai_1 U7921( .A1(n8116), .A2(n8181), .B1(n8182), .B2(n8118), .C1(n8183), .Y(n8180) );
	nand2_1 U7922( .A(n8184), .B(n8137), .Y(n8183) );
	xnor2_1 U7923( .A(n8185), .B(n8175), .Y(n8181) );
	o211ai_1 U7924( .A1(n8186), .A2(n8187), .B1(n8188), .C1(n8189), .Y(n8175) );
	mux2i_1 U7925( .A0(n8186), .A1(n8187), .S(n8137), .Y(n8189) );
	o22ai_1 U7926( .A1(n8190), .A2(n8108), .B1(n8110), .B2(n8191), .Y(n4619) );
	o22ai_1 U7927( .A1(n5538), .A2(n8111), .B1(n8112), .B2(n8191), .Y(n4618) );
	o22ai_1 U7928( .A1(n5711), .A2(n8113), .B1(n8114), .B2(n8191), .Y(n4617) );
	o221ai_1 U7929( .A1(n8192), .A2(n8116), .B1(n7251), .B2(n8118), .C1(n8119), .Y(n8191) );
	nand2_1 U7930( .A(n8184), .B(n8014), .Y(n8119) );
	inv_1 U7931( .A(n8128), .Y(n8184) );
	xnor2_1 U7932( .A(n8193), .B(n8194), .Y(n8192) );
	nand2_1 U7933( .A(n8195), .B(n8188), .Y(n8193) );
	xnor2_1 U7934( .A(n8196), .B(n8137), .Y(n8195) );
	o22ai_1 U7935( .A1(n8197), .A2(n8110), .B1(n8198), .B2(n8108), .Y(n4616) );
	nand2_1 U7936( .A(n8048), .B(n5752), .Y(n8108) );
	nand2_1 U7937( .A(n7231), .B(n5751), .Y(n8110) );
	o22ai_1 U7938( .A1(n8197), .A2(n8112), .B1(n5397), .B2(n8111), .Y(n4615) );
	nand2_1 U7939( .A(n8049), .B(n5751), .Y(n8111) );
	inv_1 U7940( .A(n124), .Y(n8112) );
	o22ai_1 U7941( .A1(n5712), .A2(n8113), .B1(n8197), .B2(n8114), .Y(n4614) );
	inv_1 U7942( .A(n123), .Y(n8114) );
	inv_1 U7943( .A(n8199), .Y(n8197) );
	o22ai_1 U7944( .A1(n8200), .A2(n8118), .B1(n8201), .B2(n8116), .Y(n8199) );
	xnor2_1 U7945( .A(n8202), .B(n8196), .Y(n8201) );
	nand2_1 U7946( .A(n8128), .B(n8116), .Y(n8118) );
	o221ai_1 U7947( .A1(n8202), .A2(n8203), .B1(n8016), .B2(n8204), .C1(n8205), .Y(n8116) );
	a21oi_1 U7948( .A1(n8206), .A2(n7937), .B1(n8207), .Y(n8205) );
	inv_1 U7949( .A(n7967), .Y(n8207) );
	a21oi_1 U7950( .A1(n7915), .A2(n8208), .B1(n7992), .Y(n8206) );
	a221oi_1 U7951( .A1(n7949), .A2(g5472), .B1(n7942), .B2(n7775), .C1(n8209), .Y(n7992) );
	nor2_1 U7952( .A(n7932), .B(n7728), .Y(n8209) );
	inv_1 U7953( .A(n7331), .Y(n7942) );
	inv_1 U7954( .A(n7333), .Y(n7949) );
	nand3_1 U7955( .A(n7956), .B(n7958), .C(n7983), .Y(n8208) );
	inv_1 U7956( .A(n7991), .Y(n7956) );
	a21oi_1 U7957( .A1(n7996), .A2(n7997), .B1(n7987), .Y(n7991) );
	inv_1 U7958( .A(n8210), .Y(n7997) );
	o221ai_1 U7959( .A1(n8211), .A2(n8212), .B1(n8213), .B2(n8214), .C1(n8215), .Y(n8210) );
	o221ai_1 U7960( .A1(n8010), .A2(n8216), .B1(n8008), .B2(n8004), .C1(n8009), .Y(n8215) );
	o22ai_1 U7961( .A1(n8009), .A2(n8008), .B1(n8216), .B2(n8004), .Y(n8214) );
	o22ai_1 U7962( .A1(n8010), .A2(n8008), .B1(n8009), .B2(n8216), .Y(n8212) );
	inv_1 U7963( .A(n7999), .Y(n8216) );
	xnor2_1 U7964( .A(n7248), .B(n8217), .Y(n7999) );
	xnor2_1 U7965( .A(n7251), .B(n8186), .Y(n8009) );
	xnor2_1 U7966( .A(n8141), .B(n8134), .Y(n8008) );
	inv_1 U7967( .A(n8213), .Y(n8010) );
	xnor2_1 U7968( .A(n8159), .B(n8157), .Y(n8213) );
	inv_1 U7969( .A(n8153), .Y(n8159) );
	inv_1 U7970( .A(n8004), .Y(n8211) );
	xnor2_1 U7971( .A(n8080), .B(n8218), .Y(n8004) );
	inv_1 U7972( .A(n8219), .Y(n7996) );
	o221ai_1 U7973( .A1(n8007), .A2(n8220), .B1(n8006), .B2(n8221), .C1(n8222), .Y(n8219) );
	o221ai_1 U7974( .A1(n8223), .A2(n8224), .B1(n8225), .B2(n8226), .C1(n8003), .Y(n8222) );
	o22ai_1 U7975( .A1(n8226), .A2(n8224), .B1(n8223), .B2(n8003), .Y(n8221) );
	inv_1 U7976( .A(n8007), .Y(n8224) );
	o22ai_1 U7977( .A1(n8223), .A2(n8225), .B1(n8226), .B2(n8003), .Y(n8220) );
	xnor2_1 U7978( .A(n8227), .B(n8124), .Y(n8003) );
	inv_1 U7979( .A(n8005), .Y(n8226) );
	xnor2_1 U7980( .A(n7240), .B(n8228), .Y(n8005) );
	inv_1 U7981( .A(n8006), .Y(n8225) );
	xnor2_1 U7982( .A(n7245), .B(n8161), .Y(n8006) );
	inv_1 U7983( .A(n7998), .Y(n8223) );
	xnor2_1 U7984( .A(n7592), .B(n8177), .Y(n7998) );
	xnor2_1 U7985( .A(n7593), .B(n8187), .Y(n8007) );
	inv_1 U7986( .A(n8017), .Y(n7915) );
	nor3_1 U7987( .A(n8016), .B(n7955), .C(n7975), .Y(n8017) );
	inv_1 U7988( .A(n7970), .Y(n7955) );
	inv_1 U7989( .A(n7978), .Y(n8204) );
	nor2_1 U7990( .A(n8229), .B(n8230), .Y(n7978) );
	inv_1 U7991( .A(n7718), .Y(n8230) );
	a21oi_1 U7992( .A1(n8231), .A2(n8137), .B1(n8232), .Y(n8203) );
	inv_1 U7993( .A(n8014), .Y(n8137) );
	o211ai_1 U7994( .A1(n8231), .A2(n8232), .B1(n8188), .C1(n7967), .Y(n8128) );
	nand2_1 U7995( .A(n7937), .B(n7939), .Y(n7967) );
	o221ai_1 U7996( .A1(n7377), .A2(n8032), .B1(n7378), .B2(n7927), .C1(n8233), .Y(n7939) );
	nand2_1 U7997( .A(g6712), .B(n7930), .Y(n8233) );
	inv_1 U7998( .A(n7739), .Y(n7930) );
	and2_0 U7999( .A(n8234), .B(n8235), .X(n7937) );
	nor4_1 U8000( .A(n8236), .B(n8237), .C(n8238), .D(n8239), .Y(n8235) );
	xnor2_1 U8001( .A(n8240), .B(n8117), .Y(n8239) );
	a222oi_1 U8002( .A1(g6518), .A2(n8241), .B1(n7231), .B2(n5432), .C1(g6368), .C2(n8242), .Y(n8240) );
	xnor2_1 U8003( .A(n8243), .B(n8227), .Y(n8238) );
	a222oi_1 U8004( .A1(g6518), .A2(n8244), .B1(n7231), .B2(n5433), .C1(g6368), .C2(n8245), .Y(n8243) );
	mux2i_1 U8005( .A0(n8246), .A1(n8247), .S(n8157), .Y(n8237) );
	nand2_1 U8006( .A(n10008), .B(n8247), .Y(n8246) );
	nand3_1 U8007( .A(n8248), .B(n8249), .C(n7976), .Y(n8236) );
	inv_1 U8008( .A(n7987), .Y(n7976) );
	nand2_1 U8009( .A(n7718), .B(n8229), .Y(n7987) );
	o21ai_0 U8010( .A1(n10009), .A2(n8048), .B1(n8250), .Y(n8229) );
	a22oi_1 U8011( .A1(g6368), .A2(n8251), .B1(g6518), .B2(n8252), .Y(n8250) );
	xnor2_1 U8012( .A(n8253), .B(n8254), .Y(n8249) );
	a222oi_1 U8013( .A1(g6518), .A2(n8255), .B1(n7231), .B2(n5440), .C1(g6368), .C2(n8256), .Y(n8254) );
	xnor2_1 U8014( .A(n8200), .B(n8257), .Y(n8248) );
	a222oi_1 U8015( .A1(g6518), .A2(n8258), .B1(n7231), .B2(n5441), .C1(g6368), .C2(n8259), .Y(n8257) );
	nor4_1 U8016( .A(n8260), .B(n8261), .C(n8262), .D(n8263), .Y(n8234) );
	mux2i_1 U8017( .A0(n8264), .A1(n8265), .S(n8266), .Y(n8263) );
	nand2_1 U8018( .A(n7615), .B(n8265), .Y(n8264) );
	mux2i_1 U8019( .A0(n8267), .A1(n8268), .S(n8149), .Y(n8262) );
	nand2_1 U8020( .A(n7612), .B(n8268), .Y(n8267) );
	mux2i_1 U8021( .A0(n8269), .A1(n8270), .S(n8141), .Y(n8261) );
	nand2_1 U8022( .A(n7285), .B(n8270), .Y(n8269) );
	nand3_1 U8023( .A(n8271), .B(n8272), .C(n8273), .Y(n8260) );
	mux2i_1 U8024( .A0(n8274), .A1(n8275), .S(n8182), .Y(n8273) );
	nor2_1 U8025( .A(n8275), .B(n5306), .Y(n8274) );
	mux2i_1 U8026( .A0(n8276), .A1(n8277), .S(n8048), .Y(n8272) );
	nand2_1 U8027( .A(n8278), .B(n8279), .Y(n8277) );
	a222oi_1 U8028( .A1(n7222), .A2(n8270), .B1(n7270), .B2(n8247), .C1(n7248), .C2(n8265), .Y(n8279) );
	a22oi_1 U8029( .A1(n5495), .A2(g6518), .B1(n5326), .B2(g6368), .Y(n8265) );
	a22oi_1 U8030( .A1(n5494), .A2(g6518), .B1(n5325), .B2(g6368), .Y(n8247) );
	a22oi_1 U8031( .A1(n5492), .A2(g6518), .B1(n5323), .B2(g6368), .Y(n8270) );
	a222oi_1 U8032( .A1(n7592), .A2(n8280), .B1(n7240), .B2(n8268), .C1(n7245), .C2(n8281), .Y(n8278) );
	inv_1 U8033( .A(n8282), .Y(n8281) );
	a22oi_1 U8034( .A1(n5493), .A2(g6518), .B1(n5324), .B2(g6368), .Y(n8268) );
	inv_1 U8035( .A(n8275), .Y(n8280) );
	o22ai_1 U8036( .A1(n9827), .A2(n8049), .B1(n9828), .B2(n8050), .Y(n8275) );
	nand2_1 U8037( .A(n8283), .B(n8284), .Y(n8276) );
	a222oi_1 U8038( .A1(n8167), .A2(n8285), .B1(n8141), .B2(n8286), .C1(n8149), .C2(n8287), .Y(n8284) );
	a222oi_1 U8039( .A1(n8182), .A2(n5306), .B1(n8266), .B2(n8288), .C1(n8157), .C2(n5375), .Y(n8283) );
	mux2i_1 U8040( .A0(n8289), .A1(n8282), .S(n8167), .Y(n8271) );
	nor2_1 U8041( .A(n8282), .B(n8285), .Y(n8289) );
	o22ai_1 U8042( .A1(n9825), .A2(n8049), .B1(n9826), .B2(n8050), .Y(n8282) );
	inv_1 U8043( .A(n8202), .Y(n8188) );
	nor2_1 U8044( .A(n7986), .B(n8014), .Y(n8202) );
	and4_1 U8045( .A(n8290), .B(n8132), .C(n8014), .D(n8291), .X(n8232) );
	nor4_1 U8046( .A(n8186), .B(n8120), .C(n8171), .D(n8185), .Y(n8291) );
	inv_1 U8047( .A(n8218), .Y(n8120) );
	nor3_1 U8048( .A(n7970), .B(n7983), .C(n7958), .Y(n8014) );
	inv_1 U8049( .A(n7975), .Y(n7983) );
	nand2_1 U8050( .A(n8050), .B(n5751), .Y(n8113) );
	o22ai_1 U8051( .A1(n8292), .A2(n5603), .B1(n8293), .B2(n8294), .Y(n4613) );
	o22ai_1 U8052( .A1(n8295), .A2(n8296), .B1(n8294), .B2(n8297), .Y(n4612) );
	inv_1 U8053( .A(n7387), .Y(n8296) );
	o22ai_1 U8054( .A1(n8298), .A2(n8299), .B1(n8294), .B2(n8300), .Y(n4611) );
	nand2_1 U8055( .A(n8047), .B(n5750), .Y(n8294) );
	nand2_1 U8056( .A(n8301), .B(n8302), .Y(n8047) );
	nor4_1 U8057( .A(n8253), .B(n8200), .C(n8157), .D(n8149), .Y(n8302) );
	inv_1 U8058( .A(n7240), .Y(n8149) );
	inv_1 U8059( .A(n7593), .Y(n8200) );
	inv_1 U8060( .A(n7251), .Y(n8253) );
	nor4_1 U8061( .A(n8266), .B(n8141), .C(n8167), .D(n8182), .Y(n8301) );
	inv_1 U8062( .A(n7592), .Y(n8182) );
	inv_1 U8063( .A(n7245), .Y(n8167) );
	inv_1 U8064( .A(n7222), .Y(n8141) );
	inv_1 U8065( .A(n7248), .Y(n8266) );
	inv_1 U8066( .A(n7389), .Y(n8299) );
	o22ai_1 U8067( .A1(n8293), .A2(n8303), .B1(n8292), .B2(n8304), .Y(n4610) );
	inv_1 U8068( .A(n7437), .Y(n8304) );
	o22ai_1 U8069( .A1(n8297), .A2(n8303), .B1(n8295), .B2(n5412), .Y(n4609) );
	o22ai_1 U8070( .A1(n8300), .A2(n8303), .B1(n8298), .B2(n8305), .Y(n4608) );
	o22ai_1 U8071( .A1(n8293), .A2(n8306), .B1(n8292), .B2(n8307), .Y(n4607) );
	inv_1 U8072( .A(n7430), .Y(n8307) );
	o22ai_1 U8073( .A1(n8297), .A2(n8306), .B1(n8295), .B2(n8308), .Y(n4606) );
	o22ai_1 U8074( .A1(n8300), .A2(n8306), .B1(n8298), .B2(n5400), .Y(n4605) );
	o22ai_1 U8075( .A1(n8293), .A2(n8309), .B1(n8292), .B2(n5677), .Y(n4604) );
	nand2_1 U8076( .A(n8293), .B(n5750), .Y(n8292) );
	nand2_1 U8077( .A(n7231), .B(n6529), .Y(n8293) );
	o22ai_1 U8078( .A1(n8297), .A2(n8309), .B1(n8295), .B2(n8252), .Y(n4603) );
	inv_1 U8079( .A(n7395), .Y(n8252) );
	nand2_1 U8080( .A(n8297), .B(n5750), .Y(n8295) );
	nand2_1 U8081( .A(g6518), .B(n6529), .Y(n8297) );
	o22ai_1 U8082( .A1(n8300), .A2(n8309), .B1(n8298), .B2(n8251), .Y(n4602) );
	inv_1 U8083( .A(n7396), .Y(n8251) );
	nand2_1 U8084( .A(n8300), .B(n5750), .Y(n8298) );
	nand4_1 U8085( .A(n132), .B(n7245), .C(n7222), .D(n8157), .Y(n8309) );
	inv_1 U8086( .A(n7270), .Y(n8157) );
	nand2_1 U8087( .A(g6368), .B(n6529), .Y(n8300) );
	o22ai_1 U8088( .A1(n8310), .A2(n5432), .B1(n8106), .B2(n8311), .Y(n4601) );
	o22ai_1 U8089( .A1(n8312), .A2(n8241), .B1(n8311), .B2(n8313), .Y(n4600) );
	inv_1 U8090( .A(n7421), .Y(n8241) );
	nor2_1 U8091( .A(RST), .B(n7267), .Y(n46) );
	o22ai_1 U8092( .A1(n8314), .A2(n8242), .B1(n8311), .B2(n8315), .Y(n4599) );
	nand2_1 U8093( .A(n8080), .B(n5749), .Y(n8311) );
	inv_1 U8094( .A(n8117), .Y(n8080) );
	o21ai_0 U8095( .A1(n7430), .A2(n8048), .B1(n8316), .Y(n8117) );
	a22oi_1 U8096( .A1(g6368), .A2(n5400), .B1(g6518), .B2(n8308), .Y(n8316) );
	inv_1 U8097( .A(n7429), .Y(n8308) );
	inv_1 U8098( .A(n7428), .Y(n8242) );
	o22ai_1 U8099( .A1(n8310), .A2(n5433), .B1(n8106), .B2(n8317), .Y(n4598) );
	o22ai_1 U8100( .A1(n8312), .A2(n8244), .B1(n8313), .B2(n8317), .Y(n4597) );
	inv_1 U8101( .A(n7431), .Y(n8244) );
	o22ai_1 U8102( .A1(n8314), .A2(n8245), .B1(n8315), .B2(n8317), .Y(n4596) );
	nand2_1 U8103( .A(n8081), .B(n5749), .Y(n8317) );
	inv_1 U8104( .A(n8227), .Y(n8081) );
	o21ai_0 U8105( .A1(n7437), .A2(n8048), .B1(n8318), .Y(n8227) );
	a22oi_1 U8106( .A1(g6368), .A2(n8305), .B1(g6518), .B2(n5412), .Y(n8318) );
	inv_1 U8107( .A(n7438), .Y(n8305) );
	inv_1 U8108( .A(n7436), .Y(n8245) );
	o22ai_1 U8109( .A1(n8106), .A2(n8319), .B1(n8286), .B2(n8310), .Y(n4595) );
	inv_1 U8110( .A(n7285), .Y(n8286) );
	o22ai_1 U8111( .A1(n8313), .A2(n8319), .B1(n8312), .B2(n5492), .Y(n4594) );
	o22ai_1 U8112( .A1(n8315), .A2(n8319), .B1(n8314), .B2(n5323), .Y(n4593) );
	inv_1 U8113( .A(n133), .Y(n8319) );
	o22ai_1 U8114( .A1(n8106), .A2(n8320), .B1(n8287), .B2(n8310), .Y(n4592) );
	inv_1 U8115( .A(n7612), .Y(n8287) );
	o22ai_1 U8116( .A1(n8320), .A2(n8313), .B1(n8312), .B2(n5493), .Y(n4591) );
	o22ai_1 U8117( .A1(n8320), .A2(n8315), .B1(n8314), .B2(n5324), .Y(n4590) );
	inv_1 U8118( .A(n132), .Y(n8320) );
	o22ai_1 U8119( .A1(n8106), .A2(n8321), .B1(n5375), .B2(n8310), .Y(n4589) );
	o22ai_1 U8120( .A1(n8313), .A2(n8321), .B1(n8312), .B2(n5494), .Y(n4588) );
	o22ai_1 U8121( .A1(n8315), .A2(n8321), .B1(n8314), .B2(n5325), .Y(n4587) );
	inv_1 U8122( .A(n131), .Y(n8321) );
	o22ai_1 U8123( .A1(n8106), .A2(n8322), .B1(n8285), .B2(n8310), .Y(n4586) );
	inv_1 U8124( .A(n7323), .Y(n8285) );
	o22ai_1 U8125( .A1(n8313), .A2(n8322), .B1(n8312), .B2(n5656), .Y(n4585) );
	o22ai_1 U8126( .A1(n8315), .A2(n8322), .B1(n8314), .B2(n5639), .Y(n4584) );
	inv_1 U8127( .A(n130), .Y(n8322) );
	o22ai_1 U8128( .A1(n8106), .A2(n8323), .B1(n8288), .B2(n8310), .Y(n4583) );
	inv_1 U8129( .A(n7615), .Y(n8288) );
	o22ai_1 U8130( .A1(n8313), .A2(n8323), .B1(n8312), .B2(n5495), .Y(n4582) );
	o22ai_1 U8131( .A1(n8315), .A2(n8323), .B1(n8314), .B2(n5326), .Y(n4581) );
	inv_1 U8132( .A(n129), .Y(n8323) );
	o22ai_1 U8133( .A1(n8106), .A2(n8324), .B1(n5306), .B2(n8310), .Y(n4580) );
	o22ai_1 U8134( .A1(n8313), .A2(n8324), .B1(n8312), .B2(n5657), .Y(n4579) );
	o22ai_1 U8135( .A1(n8315), .A2(n8324), .B1(n8314), .B2(n5640), .Y(n4578) );
	inv_1 U8136( .A(n128), .Y(n8324) );
	o22ai_1 U8137( .A1(n8106), .A2(n8306), .B1(n8310), .B2(n5440), .Y(n4577) );
	o22ai_1 U8138( .A1(n8306), .A2(n8313), .B1(n8312), .B2(n8255), .Y(n4576) );
	inv_1 U8139( .A(n7412), .Y(n8255) );
	o22ai_1 U8140( .A1(n8306), .A2(n8315), .B1(n8314), .B2(n8256), .Y(n4575) );
	inv_1 U8141( .A(n7422), .Y(n8256) );
	inv_1 U8142( .A(n126), .Y(n8306) );
	o22ai_1 U8143( .A1(n8106), .A2(n8303), .B1(n8310), .B2(n5441), .Y(n4574) );
	nand2_1 U8144( .A(n5755), .B(n8106), .Y(n8310) );
	nand2_1 U8145( .A(n7718), .B(n7231), .Y(n8106) );
	o22ai_1 U8146( .A1(n8303), .A2(n8313), .B1(n8312), .B2(n8258), .Y(n4573) );
	inv_1 U8147( .A(n7423), .Y(n8258) );
	nand2_1 U8148( .A(n5755), .B(n8313), .Y(n8312) );
	nand2_1 U8149( .A(n7718), .B(g6518), .Y(n8313) );
	o22ai_1 U8150( .A1(n8303), .A2(n8315), .B1(n8314), .B2(n8259), .Y(n4572) );
	inv_1 U8151( .A(n7432), .Y(n8259) );
	nand2_1 U8152( .A(n5755), .B(n8315), .Y(n8314) );
	nand2_1 U8153( .A(n7718), .B(g6368), .Y(n8315) );
	inv_1 U8154( .A(n125), .Y(n8303) );
	a21oi_1 U8155( .A1(n8325), .A2(n8326), .B1(n8327), .Y(n4571) );
	a21oi_1 U8156( .A1(n5336), .A2(n8328), .B1(n8329), .Y(n4570) );
	a21oi_1 U8157( .A1(n5545), .A2(n8330), .B1(n8331), .Y(n4569) );
	o22ai_1 U8158( .A1(n8332), .A2(n8333), .B1(n8334), .B2(n8335), .Y(n4568) );
	inv_1 U8159( .A(n7547), .Y(n8333) );
	o22ai_1 U8160( .A1(n8336), .A2(n8337), .B1(n8334), .B2(n8338), .Y(n4567) );
	inv_1 U8161( .A(n7570), .Y(n8337) );
	o22ai_1 U8162( .A1(n8339), .A2(n8340), .B1(n8334), .B2(n8341), .Y(n4566) );
	nand4_1 U8163( .A(n8342), .B(n8343), .C(n8344), .D(n8345), .Y(n8334) );
	a222oi_1 U8164( .A1(g6911), .A2(n8346), .B1(n7239), .B2(n8347), .C1(g6677), .C2(n5393), .Y(n8345) );
	nand2_1 U8165( .A(n9870), .B(n10010), .Y(n8347) );
	nand4_1 U8166( .A(n8348), .B(n8349), .C(n8350), .D(n8351), .Y(n8344) );
	nor3_1 U8167( .A(n8352), .B(n8353), .C(n8354), .Y(n8351) );
	xor2_1 U8168( .A(n8355), .B(n10012), .X(n8354) );
	xor2_1 U8169( .A(n8356), .B(n7688), .X(n8353) );
	nand3_1 U8170( .A(n8357), .B(n8358), .C(n8359), .Y(n8352) );
	xor2_1 U8171( .A(n9954), .B(n8360), .X(n8359) );
	xnor2_1 U8172( .A(n10013), .B(n8361), .Y(n8358) );
	xnor2_1 U8173( .A(n10014), .B(n8362), .Y(n8357) );
	nor3_1 U8174( .A(n8363), .B(n8364), .C(n8365), .Y(n8350) );
	xor2_1 U8175( .A(n8366), .B(n9974), .X(n8365) );
	xor2_1 U8176( .A(n8367), .B(n10011), .X(n8364) );
	xnor2_1 U8177( .A(n8368), .B(n8369), .Y(n8363) );
	xnor2_1 U8178( .A(n7298), .B(n8370), .Y(n8349) );
	xnor2_1 U8179( .A(n7694), .B(n8371), .Y(n8348) );
	o22ai_1 U8180( .A1(n8327), .A2(n5573), .B1(n8372), .B2(n8373), .Y(n4565) );
	o22ai_1 U8181( .A1(n8329), .A2(n8374), .B1(n8372), .B2(n8375), .Y(n4564) );
	o22ai_1 U8182( .A1(n8331), .A2(n5468), .B1(n8372), .B2(n5819), .Y(n4563) );
	nand2_1 U8183( .A(n8376), .B(n9975), .Y(n8372) );
	o22ai_1 U8184( .A1(n8327), .A2(n5625), .B1(n8373), .B2(n8377), .Y(n4562) );
	o21ai_0 U8185( .A1(n5364), .A2(n8378), .B1(n5756), .Y(n8327) );
	o22ai_1 U8186( .A1(n8329), .A2(n8346), .B1(n8375), .B2(n8377), .Y(n4561) );
	inv_1 U8187( .A(n5292), .Y(n8375) );
	nor2_1 U8188( .A(n8379), .B(RST), .Y(n5292) );
	inv_1 U8189( .A(n7450), .Y(n8346) );
	o22ai_1 U8190( .A1(n8331), .A2(n5393), .B1(n5819), .B2(n8377), .Y(n4560) );
	nand2_1 U8191( .A(n8380), .B(n9975), .Y(n8377) );
	nand2_1 U8192( .A(g6677), .B(n5749), .Y(n5819) );
	o21ai_0 U8193( .A1(n5364), .A2(n8381), .B1(n5755), .Y(n8331) );
	o22ai_1 U8194( .A1(n8332), .A2(n8382), .B1(n10013), .B2(n8335), .Y(n4559) );
	inv_1 U8195( .A(n7549), .Y(n8382) );
	o22ai_1 U8196( .A1(n8336), .A2(n8383), .B1(n10013), .B2(n8338), .Y(n4558) );
	inv_1 U8197( .A(n7548), .Y(n8383) );
	o22ai_1 U8198( .A1(n8339), .A2(n5463), .B1(n10013), .B2(n8341), .Y(n4557) );
	o22ai_1 U8199( .A1(n8332), .A2(n8384), .B1(n10014), .B2(n8335), .Y(n4556) );
	inv_1 U8200( .A(n7551), .Y(n8384) );
	o22ai_1 U8201( .A1(n8336), .A2(n8385), .B1(n10014), .B2(n8338), .Y(n4555) );
	inv_1 U8202( .A(n7550), .Y(n8385) );
	o22ai_1 U8203( .A1(n8339), .A2(n5466), .B1(n10014), .B2(n8341), .Y(n4554) );
	o22ai_1 U8204( .A1(n8332), .A2(n8386), .B1(n7694), .B2(n8335), .Y(n4553) );
	inv_1 U8205( .A(n7560), .Y(n8386) );
	o22ai_1 U8206( .A1(n8336), .A2(n8387), .B1(n7694), .B2(n8338), .Y(n4552) );
	inv_1 U8207( .A(n7559), .Y(n8387) );
	o22ai_1 U8208( .A1(n8339), .A2(n5472), .B1(n7694), .B2(n8341), .Y(n4551) );
	o22ai_1 U8209( .A1(n8332), .A2(n8388), .B1(n10011), .B2(n8335), .Y(n4550) );
	inv_1 U8210( .A(n7562), .Y(n8388) );
	o22ai_1 U8211( .A1(n8336), .A2(n8389), .B1(n10011), .B2(n8338), .Y(n4549) );
	inv_1 U8212( .A(n7561), .Y(n8389) );
	o22ai_1 U8213( .A1(n8339), .A2(n5469), .B1(n10011), .B2(n8341), .Y(n4548) );
	o22ai_1 U8214( .A1(n8332), .A2(n8390), .B1(n7298), .B2(n8335), .Y(n4547) );
	inv_1 U8215( .A(n7564), .Y(n8390) );
	o22ai_1 U8216( .A1(n8336), .A2(n8391), .B1(n7298), .B2(n8338), .Y(n4546) );
	inv_1 U8217( .A(n7563), .Y(n8391) );
	o22ai_1 U8218( .A1(n8339), .A2(n5470), .B1(n7298), .B2(n8341), .Y(n4545) );
	o22ai_1 U8219( .A1(n8332), .A2(n8392), .B1(n10012), .B2(n8335), .Y(n4544) );
	inv_1 U8220( .A(n7566), .Y(n8392) );
	o22ai_1 U8221( .A1(n8336), .A2(n8393), .B1(n10012), .B2(n8338), .Y(n4543) );
	inv_1 U8222( .A(n7565), .Y(n8393) );
	o22ai_1 U8223( .A1(n8339), .A2(n5467), .B1(n10012), .B2(n8341), .Y(n4542) );
	o22ai_1 U8224( .A1(n8332), .A2(n8394), .B1(n7302), .B2(n8335), .Y(n4541) );
	inv_1 U8225( .A(n7557), .Y(n8394) );
	o22ai_1 U8226( .A1(n8336), .A2(n8395), .B1(n7302), .B2(n8338), .Y(n4540) );
	inv_1 U8227( .A(n7556), .Y(n8395) );
	o22ai_1 U8228( .A1(n8339), .A2(n5465), .B1(n7302), .B2(n8341), .Y(n4539) );
	o22ai_1 U8229( .A1(n8332), .A2(n8396), .B1(n9954), .B2(n8335), .Y(n4538) );
	o22ai_1 U8230( .A1(n8336), .A2(n8397), .B1(n9954), .B2(n8338), .Y(n4537) );
	o22ai_1 U8231( .A1(n8339), .A2(n5626), .B1(n9954), .B2(n8341), .Y(n4536) );
	o22ai_1 U8232( .A1(n8332), .A2(n8398), .B1(n7688), .B2(n8335), .Y(n4535) );
	inv_1 U8233( .A(n7555), .Y(n8398) );
	o22ai_1 U8234( .A1(n8336), .A2(n8399), .B1(n7688), .B2(n8338), .Y(n4534) );
	inv_1 U8235( .A(n7554), .Y(n8399) );
	o22ai_1 U8236( .A1(n8339), .A2(n5464), .B1(n7688), .B2(n8341), .Y(n4533) );
	o22ai_1 U8237( .A1(n8332), .A2(n8400), .B1(n9974), .B2(n8335), .Y(n4532) );
	or2_0 U8238( .A(n8326), .B(RST), .X(n8335) );
	inv_1 U8239( .A(n7568), .Y(n8400) );
	nand2_1 U8240( .A(n5756), .B(n8326), .Y(n8332) );
	nand3_1 U8241( .A(n9976), .B(n8401), .C(n9869), .Y(n8326) );
	o22ai_1 U8242( .A1(n8336), .A2(n8402), .B1(n9974), .B2(n8338), .Y(n4531) );
	or2_0 U8243( .A(n8328), .B(RST), .X(n8338) );
	inv_1 U8244( .A(n7567), .Y(n8402) );
	nand2_1 U8245( .A(n5756), .B(n8328), .Y(n8336) );
	nand2_1 U8246( .A(n8403), .B(g6911), .Y(n8328) );
	o22ai_1 U8247( .A1(n8339), .A2(n5471), .B1(n9974), .B2(n8341), .Y(n4530) );
	or2_0 U8248( .A(n8330), .B(RST), .X(n8341) );
	nand2_1 U8249( .A(n5756), .B(n8330), .Y(n8339) );
	nand2_1 U8250( .A(n8403), .B(g6677), .Y(n8330) );
	and3_1 U8251( .A(n9976), .B(n8404), .C(n9869), .X(n8403) );
	nor2_1 U8252( .A(n8405), .B(n8329), .Y(n4529) );
	xnor2_1 U8253( .A(n8406), .B(n10013), .Y(n8405) );
	a211oi_1 U8254( .A1(n5368), .A2(n8407), .B1(n8329), .C1(n8406), .Y(n4528) );
	nor2_1 U8255( .A(n8407), .B(n5368), .Y(n8406) );
	nor3_1 U8256( .A(n8329), .B(n8408), .C(n8409), .Y(n4527) );
	a21oi_1 U8257( .A1(n8410), .A2(n10011), .B1(n7694), .Y(n8409) );
	inv_1 U8258( .A(n8407), .Y(n8408) );
	nand3_1 U8259( .A(n7694), .B(n10011), .C(n8410), .Y(n8407) );
	nor2_1 U8260( .A(n8411), .B(n8329), .Y(n4526) );
	xnor2_1 U8261( .A(n8410), .B(n10011), .Y(n8411) );
	nor3_1 U8262( .A(n8329), .B(n8410), .C(n8412), .Y(n4525) );
	a21oi_1 U8263( .A1(n8413), .A2(n10012), .B1(n7298), .Y(n8412) );
	and3_1 U8264( .A(n7298), .B(n10012), .C(n8413), .X(n8410) );
	nor2_1 U8265( .A(n8414), .B(n8329), .Y(n4524) );
	xnor2_1 U8266( .A(n10012), .B(n8413), .Y(n8414) );
	a211oi_1 U8267( .A1(n8369), .A2(n5818), .B1(n8329), .C1(n8413), .Y(n4523) );
	nor2_1 U8268( .A(n5818), .B(n8369), .Y(n8413) );
	nand2_1 U8269( .A(n9954), .B(n5816), .Y(n5818) );
	inv_1 U8270( .A(n7302), .Y(n8369) );
	nor3_1 U8271( .A(n8329), .B(n5816), .C(n8415), .Y(n4522) );
	a21oi_1 U8272( .A1(n9974), .A2(n8401), .B1(n7688), .Y(n8415) );
	and3_1 U8273( .A(n7688), .B(n8401), .C(n9974), .X(n5816) );
	nor2_1 U8274( .A(n8416), .B(n8329), .Y(n4521) );
	inv_1 U8275( .A(n5817), .Y(n8329) );
	a21oi_1 U8276( .A1(g6911), .A2(n9975), .B1(RST), .Y(n5817) );
	xnor2_1 U8277( .A(n8401), .B(n9974), .Y(n8416) );
	nor2_1 U8278( .A(n8378), .B(n7278), .Y(n8401) );
	o32ai_1 U8279( .A1(n8404), .A2(n7239), .A3(RST), .B1(n5981), .B2(n8373), .Y(n4520) );
	inv_1 U8280( .A(n7278), .Y(n8404) );
	o32ai_1 U8281( .A1(n5364), .A2(n7239), .A3(RST), .B1(n8373), .B2(n8417), .Y(n4519) );
	nand2_1 U8282( .A(n7239), .B(n5748), .Y(n8373) );
	o22ai_1 U8283( .A1(n5983), .A2(n8418), .B1(n5984), .B2(n5394), .Y(n4518) );
	and2_0 U8284( .A(n5762), .B(g16297), .X(n4517) );
	and2_0 U8285( .A(n5747), .B(n8419), .X(n4516) );
	o22ai_1 U8286( .A1(n5565), .A2(n8420), .B1(n8421), .B2(n8422), .Y(n4515) );
	o22ai_1 U8287( .A1(n5730), .A2(n8423), .B1(n8422), .B2(n8424), .Y(n4514) );
	o22ai_1 U8288( .A1(n8425), .A2(n8426), .B1(n8422), .B2(n8427), .Y(n4513) );
	nand3_1 U8289( .A(n7591), .B(n8380), .C(n8428), .Y(n8422) );
	inv_1 U8290( .A(n7639), .Y(n8425) );
	o22ai_1 U8291( .A1(n5558), .A2(n8420), .B1(n8429), .B2(n8421), .Y(n4512) );
	o22ai_1 U8292( .A1(n5348), .A2(n8423), .B1(n8429), .B2(n8424), .Y(n4511) );
	o22ai_1 U8293( .A1(n8429), .A2(n8427), .B1(n8430), .B2(n8426), .Y(n4510) );
	inv_1 U8294( .A(n7665), .Y(n8430) );
	mux2i_1 U8295( .A0(n8431), .A1(n8432), .S(n5999), .Y(n8429) );
	nor2_1 U8296( .A(n8433), .B(n8434), .Y(n8431) );
	mux2_1 U8297( .A0(n8435), .A1(n8436), .S(n8437), .X(n8433) );
	o22ai_1 U8298( .A1(n5557), .A2(n8420), .B1(n8438), .B2(n8421), .Y(n4509) );
	o22ai_1 U8299( .A1(n5347), .A2(n8423), .B1(n8438), .B2(n8424), .Y(n4508) );
	o22ai_1 U8300( .A1(n8438), .A2(n8427), .B1(n8439), .B2(n8426), .Y(n4507) );
	inv_1 U8301( .A(n7664), .Y(n8439) );
	mux2i_1 U8302( .A0(n8440), .A1(n8441), .S(n5999), .Y(n8438) );
	nor2_1 U8303( .A(n8442), .B(n8443), .Y(n8440) );
	inv_1 U8304( .A(n8436), .Y(n8443) );
	a222oi_1 U8305( .A1(n8444), .A2(n8445), .B1(n8446), .B2(n8447), .C1(n8448), .C2(n8449), .Y(n8436) );
	o22ai_1 U8306( .A1(n8444), .A2(n8450), .B1(n8451), .B2(n8452), .Y(n8449) );
	o22ai_1 U8307( .A1(n8453), .A2(n8454), .B1(n8455), .B2(n8444), .Y(n8447) );
	a21oi_1 U8308( .A1(n8456), .A2(n8457), .B1(n8458), .Y(n8455) );
	o22ai_1 U8309( .A1(n8459), .A2(n8460), .B1(n8461), .B2(n8462), .Y(n8456) );
	o32ai_1 U8310( .A1(n8448), .A2(n8463), .A3(n8461), .B1(n8464), .B2(n8446), .Y(n8445) );
	a21oi_1 U8311( .A1(n8465), .A2(n8461), .B1(n8466), .Y(n8464) );
	mux2i_1 U8312( .A0(n8459), .A1(n8467), .S(n8457), .Y(n8466) );
	or2_0 U8313( .A(n8454), .B(n8460), .X(n8467) );
	mux2i_1 U8314( .A0(n8434), .A1(n8437), .S(n8435), .Y(n8442) );
	inv_1 U8315( .A(n8468), .Y(n8437) );
	nand2_1 U8316( .A(n8469), .B(n8470), .Y(n8434) );
	nand3_1 U8317( .A(n8460), .B(n8471), .C(n8472), .Y(n8470) );
	inv_1 U8318( .A(n8453), .Y(n8460) );
	mux2i_1 U8319( .A0(n8473), .A1(n8474), .S(n8444), .Y(n8469) );
	o221ai_1 U8320( .A1(n8475), .A2(n15067), .B1(n5356), .B2(n15066), .C1(n8476), .Y(n8444) );
	nand2_1 U8321( .A(g349), .B(g5629), .Y(n8476) );
	o221ai_1 U8322( .A1(n8477), .A2(n8450), .B1(n8448), .B2(n8478), .C1(n8479), .Y(n8474) );
	mux2i_1 U8323( .A0(n8480), .A1(n8481), .S(n8446), .Y(n8479) );
	nor2_1 U8324( .A(n8482), .B(n8457), .Y(n8481) );
	a21oi_1 U8325( .A1(n8463), .A2(n8477), .B1(n8471), .Y(n8482) );
	nor2_1 U8326( .A(n8453), .B(n8483), .Y(n8480) );
	a221oi_1 U8327( .A1(n8484), .A2(n8453), .B1(n8485), .B2(n8471), .C1(n8458), .Y(n8478) );
	inv_1 U8328( .A(n8457), .Y(n8448) );
	o21ai_0 U8329( .A1(n8463), .A2(n8486), .B1(n8487), .Y(n8473) );
	mux2i_1 U8330( .A0(n8488), .A1(n8489), .S(n8457), .Y(n8487) );
	o221ai_1 U8331( .A1(n8475), .A2(n15073), .B1(n5356), .B2(n15071), .C1(n8490), .Y(n8457) );
	nand2_1 U8332( .A(g364), .B(g5629), .Y(n8490) );
	o22ai_1 U8333( .A1(n8477), .A2(n8454), .B1(n8491), .B2(n8452), .Y(n8489) );
	inv_1 U8334( .A(n8485), .Y(n8452) );
	nor2_1 U8335( .A(n8446), .B(n8461), .Y(n8485) );
	nor3_1 U8336( .A(n8484), .B(n8458), .C(n8472), .Y(n8488) );
	nor2_1 U8337( .A(n8477), .B(n8451), .Y(n8458) );
	a21oi_1 U8338( .A1(n8453), .A2(n8446), .B1(n8461), .Y(n8486) );
	inv_1 U8339( .A(n8477), .Y(n8461) );
	o221ai_1 U8340( .A1(n8475), .A2(n15069), .B1(n5356), .B2(n15068), .C1(n8492), .Y(n8477) );
	nand2_1 U8341( .A(g379), .B(g5629), .Y(n8492) );
	o221ai_1 U8342( .A1(n8475), .A2(n15065), .B1(n5356), .B2(n15064), .C1(n8493), .Y(n8453) );
	nand2_1 U8343( .A(g5629), .B(g394), .Y(n8493) );
	o22ai_1 U8344( .A1(n8420), .A2(n5627), .B1(n8421), .B2(n8494), .Y(n4506) );
	o22ai_1 U8345( .A1(n8423), .A2(n5599), .B1(n8424), .B2(n8494), .Y(n4505) );
	o22ai_1 U8346( .A1(n8426), .A2(n5408), .B1(n8427), .B2(n8494), .Y(n4504) );
	nand2_1 U8347( .A(n8435), .B(n5999), .Y(n8494) );
	o211ai_1 U8348( .A1(n8495), .A2(n5408), .B1(n8496), .C1(n8497), .Y(n8435) );
	a22oi_1 U8349( .A1(n9830), .A2(g6642), .B1(n9829), .B2(n7227), .Y(n8497) );
	nand3_1 U8350( .A(n7256), .B(n8498), .C(g542), .Y(n8496) );
	o22ai_1 U8351( .A1(n8420), .A2(n5628), .B1(n8421), .B2(n8499), .Y(n4503) );
	o22ai_1 U8352( .A1(n8423), .A2(n5600), .B1(n8424), .B2(n8499), .Y(n4502) );
	inv_1 U8353( .A(n110), .Y(n8424) );
	nand2_1 U8354( .A(n8500), .B(n5748), .Y(n8423) );
	o22ai_1 U8355( .A1(n8426), .A2(n5409), .B1(n8427), .B2(n8499), .Y(n4501) );
	nand2_1 U8356( .A(n8468), .B(n5999), .Y(n8499) );
	o211ai_1 U8357( .A1(n8495), .A2(n5409), .B1(n8501), .C1(n8502), .Y(n8468) );
	a22oi_1 U8358( .A1(n9832), .A2(g6642), .B1(n9831), .B2(n7227), .Y(n8502) );
	nand3_1 U8359( .A(n7256), .B(n8503), .C(g524), .Y(n8501) );
	inv_1 U8360( .A(n109), .Y(n8427) );
	nand2_1 U8361( .A(n5756), .B(n8495), .Y(n8426) );
	o22ai_1 U8362( .A1(n8504), .A2(n8505), .B1(n8506), .B2(n8507), .Y(n4500) );
	inv_1 U8363( .A(n7373), .Y(n8507) );
	nor2_1 U8364( .A(RST), .B(n7232), .Y(n45) );
	o22ai_1 U8365( .A1(n8504), .A2(n8508), .B1(n8509), .B2(n8510), .Y(n4499) );
	inv_1 U8366( .A(n7374), .Y(n8510) );
	o22ai_1 U8367( .A1(n8504), .A2(n8511), .B1(n8512), .B2(n5516), .Y(n4498) );
	o21ai_0 U8368( .A1(n8454), .A2(n8513), .B1(n5748), .Y(n8504) );
	nand2_1 U8369( .A(n8451), .B(n8459), .Y(n8454) );
	o22ai_1 U8370( .A1(n8505), .A2(n8514), .B1(n8506), .B2(n8515), .Y(n4497) );
	inv_1 U8371( .A(n7367), .Y(n8515) );
	o22ai_1 U8372( .A1(n8508), .A2(n8514), .B1(n8509), .B2(n8516), .Y(n4496) );
	inv_1 U8373( .A(n7368), .Y(n8516) );
	o22ai_1 U8374( .A1(n8511), .A2(n8514), .B1(n8512), .B2(n5515), .Y(n4495) );
	o221ai_1 U8375( .A1(n8451), .A2(n8517), .B1(n8518), .B2(n8462), .C1(n5744), .Y(n8514) );
	inv_1 U8376( .A(n8465), .Y(n8462) );
	nor2_1 U8377( .A(n8483), .B(n8491), .Y(n8465) );
	mux2i_1 U8378( .A0(n5984), .A1(n5983), .S(n8446), .Y(n8517) );
	inv_1 U8379( .A(n6098), .Y(n5984) );
	o22ai_1 U8380( .A1(n8505), .A2(n8519), .B1(n8506), .B2(n8520), .Y(n4494) );
	inv_1 U8381( .A(n7369), .Y(n8520) );
	o22ai_1 U8382( .A1(n8508), .A2(n8519), .B1(n8509), .B2(n8521), .Y(n4493) );
	inv_1 U8383( .A(n7370), .Y(n8521) );
	o22ai_1 U8384( .A1(n8511), .A2(n8519), .B1(n8512), .B2(n5514), .Y(n4492) );
	o211ai_1 U8385( .A1(n8459), .A2(n8518), .B1(n8450), .C1(n5740), .Y(n8519) );
	inv_1 U8386( .A(n8513), .Y(n8518) );
	xnor2_1 U8387( .A(n8472), .B(n5983), .Y(n8513) );
	inv_1 U8388( .A(n8446), .Y(n8472) );
	o22ai_1 U8389( .A1(n8505), .A2(n8522), .B1(n8506), .B2(n8523), .Y(n4491) );
	inv_1 U8390( .A(n7371), .Y(n8523) );
	nand2_1 U8391( .A(n8505), .B(n5748), .Y(n8506) );
	nand2_1 U8392( .A(n7227), .B(n8419), .Y(n8505) );
	o22ai_1 U8393( .A1(n8508), .A2(n8522), .B1(n8509), .B2(n8524), .Y(n4490) );
	inv_1 U8394( .A(n7372), .Y(n8524) );
	nand2_1 U8395( .A(n8508), .B(n5748), .Y(n8509) );
	nand2_1 U8396( .A(g6642), .B(n8419), .Y(n8508) );
	o22ai_1 U8397( .A1(n8511), .A2(n8522), .B1(n8512), .B2(n5513), .Y(n4489) );
	nand2_1 U8398( .A(n8511), .B(n5748), .Y(n8512) );
	o221ai_1 U8399( .A1(n6098), .A2(n8463), .B1(g3229), .B2(n8450), .C1(n8525), .Y(n8522) );
	a21oi_1 U8400( .A1(n8526), .A2(n8446), .B1(RST), .Y(n8525) );
	o221ai_1 U8401( .A1(n7372), .A2(n8500), .B1(n7371), .B2(n8527), .C1(n8528), .Y(n8446) );
	nand2_1 U8402( .A(g6485), .B(n5513), .Y(n8528) );
	o22ai_1 U8403( .A1(n8459), .A2(n5983), .B1(n8529), .B2(n8483), .Y(n8526) );
	nor2_1 U8404( .A(n8451), .B(n5983), .Y(n8529) );
	inv_1 U8405( .A(n8471), .Y(n8459) );
	inv_1 U8406( .A(n8484), .Y(n8450) );
	nor2_1 U8407( .A(n8471), .B(n8451), .Y(n8484) );
	inv_1 U8408( .A(n8491), .Y(n8451) );
	o221ai_1 U8409( .A1(n7370), .A2(n8500), .B1(n7369), .B2(n8527), .C1(n8530), .Y(n8491) );
	nand2_1 U8410( .A(g6485), .B(n5514), .Y(n8530) );
	o221ai_1 U8411( .A1(n7368), .A2(n8500), .B1(n7367), .B2(n8527), .C1(n8531), .Y(n8471) );
	nand2_1 U8412( .A(g6485), .B(n5515), .Y(n8531) );
	inv_1 U8413( .A(n8483), .Y(n8463) );
	o221ai_1 U8414( .A1(n7374), .A2(n8500), .B1(n7373), .B2(n8527), .C1(n8532), .Y(n8483) );
	nand2_1 U8415( .A(g6485), .B(n5516), .Y(n8532) );
	nand2_1 U8416( .A(g6485), .B(n8419), .Y(n8511) );
	o32ai_1 U8417( .A1(n8533), .A2(n8380), .A3(n8417), .B1(n6755), .B2(n8534), .Y(n8419) );
	nor2_1 U8418( .A(n8428), .B(n8376), .Y(n8534) );
	inv_1 U8419( .A(n8432), .Y(n8376) );
	inv_1 U8420( .A(n8533), .Y(n8428) );
	inv_1 U8421( .A(n8441), .Y(n8380) );
	o21ai_0 U8422( .A1(n8527), .A2(n5565), .B1(n8535), .Y(n8533) );
	a22oi_1 U8423( .A1(n7639), .A2(g6485), .B1(n9833), .B2(g6642), .Y(n8535) );
	and2_0 U8424( .A(g558), .B(n5764), .X(n4488) );
	o22ai_1 U8425( .A1(n8536), .A2(n8537), .B1(n8538), .B2(n5658), .Y(n4486) );
	o22ai_1 U8426( .A1(n8536), .A2(n8539), .B1(n8540), .B2(n8541), .Y(n4485) );
	inv_1 U8427( .A(n7462), .Y(n8541) );
	o22ai_1 U8428( .A1(n8536), .A2(n8542), .B1(n8543), .B2(n5425), .Y(n4484) );
	o22ai_1 U8429( .A1(n8537), .A2(n8544), .B1(n8538), .B2(n5659), .Y(n4483) );
	o22ai_1 U8430( .A1(n8539), .A2(n8544), .B1(n8540), .B2(n8545), .Y(n4482) );
	inv_1 U8431( .A(n7458), .Y(n8545) );
	o22ai_1 U8432( .A1(n8542), .A2(n8544), .B1(n8543), .B2(n5426), .Y(n4481) );
	o22ai_1 U8433( .A1(n8546), .A2(n8537), .B1(n8538), .B2(n5660), .Y(n4480) );
	or2_0 U8434( .A(RST), .B(n7259), .X(n8538) );
	o22ai_1 U8435( .A1(n8546), .A2(n8539), .B1(n8540), .B2(n8547), .Y(n4479) );
	inv_1 U8436( .A(n7456), .Y(n8547) );
	or2_0 U8437( .A(RST), .B(g7956), .X(n8540) );
	o22ai_1 U8438( .A1(n8546), .A2(n8542), .B1(n8543), .B2(n5424), .Y(n4478) );
	or2_0 U8439( .A(RST), .B(g7909), .X(n8543) );
	and2_0 U8440( .A(g568), .B(n5765), .X(n4477) );
	and2_0 U8441( .A(g574), .B(n5765), .X(n4476) );
	and2_0 U8442( .A(g572), .B(n5765), .X(n4475) );
	and2_0 U8443( .A(g564), .B(n5765), .X(n4474) );
	o22ai_1 U8444( .A1(n8417), .A2(n8420), .B1(n8421), .B2(n8548), .Y(n4473) );
	o22ai_1 U8445( .A1(n8420), .A2(n8548), .B1(n9977), .B2(n8421), .Y(n4472) );
	o22ai_1 U8446( .A1(n8420), .A2(n5592), .B1(n6118), .B2(n8421), .Y(n4471) );
	nand2_1 U8447( .A(n7227), .B(n5748), .Y(n8421) );
	inv_1 U8448( .A(n5999), .Y(n6118) );
	nand3_1 U8449( .A(n9955), .B(n9956), .C(n8549), .Y(n5999) );
	nor3_1 U8450( .A(n5874), .B(n10034), .C(n7704), .Y(n8549) );
	nand4_1 U8451( .A(n7283), .B(n7254), .C(n7326), .D(n8550), .Y(n5874) );
	nor4_1 U8452( .A(n10082), .B(n10083), .C(n7716), .D(n8551), .Y(n8550) );
	inv_1 U8453( .A(n7249), .Y(n8551) );
	nand2_1 U8454( .A(n8527), .B(n5748), .Y(n8420) );
	nor2_1 U8455( .A(RST), .B(n8475), .Y(n4470) );
	inv_1 U8456( .A(g5648), .Y(n8475) );
	and2_0 U8457( .A(g397), .B(n5765), .X(n4469) );
	and2_0 U8458( .A(g395), .B(n5764), .X(n4468) );
	and2_0 U8459( .A(g382), .B(n5765), .X(n4467) );
	and2_0 U8460( .A(g380), .B(n5765), .X(n4466) );
	and2_0 U8461( .A(g367), .B(n5764), .X(n4465) );
	and2_0 U8462( .A(g365), .B(n5765), .X(n4464) );
	and2_0 U8463( .A(g352), .B(n5765), .X(n4463) );
	and2_0 U8464( .A(g350), .B(n5764), .X(n4462) );
	a221oi_1 U8465( .A1(n8552), .A2(n8553), .B1(n8554), .B2(n8555), .C1(RST), .Y(n4461) );
	nor4_1 U8466( .A(n8556), .B(n8557), .C(n8558), .D(n8559), .Y(n8553) );
	xnor2_1 U8467( .A(n7712), .B(n8560), .Y(n8559) );
	xor2_1 U8468( .A(n8561), .B(n10029), .X(n8558) );
	xor2_1 U8469( .A(n8562), .B(n7708), .X(n8557) );
	nand3_1 U8470( .A(n8563), .B(n6131), .C(n8564), .Y(n8556) );
	xnor2_1 U8471( .A(n10025), .B(n8565), .Y(n8564) );
	nor4_1 U8472( .A(n8566), .B(n8567), .C(n8568), .D(n8569), .Y(n8552) );
	xnor2_1 U8473( .A(n7306), .B(n8570), .Y(n8569) );
	xnor2_1 U8474( .A(n7702), .B(n8571), .Y(n8568) );
	xnor2_1 U8475( .A(n10028), .B(n8572), .Y(n8567) );
	nand3_1 U8476( .A(n8573), .B(n8574), .C(n8575), .Y(n8566) );
	xnor2_1 U8477( .A(n10026), .B(n8576), .Y(n8575) );
	xnor2_1 U8478( .A(n10027), .B(n8577), .Y(n8574) );
	xnor2_1 U8479( .A(n7304), .B(n8578), .Y(n8573) );
	nor2_1 U8480( .A(RST), .B(n7921), .Y(n4460) );
	mux2i_1 U8481( .A0(n15426), .A1(n8579), .S(n7745), .Y(n7921) );
	nor2_1 U8482( .A(g6447), .B(n5394), .Y(n8579) );
	nor2_1 U8483( .A(RST), .B(n8580), .Y(n4459) );
	and2_0 U8484( .A(g290), .B(n5765), .X(n4458) );
	o22ai_1 U8485( .A1(n8581), .A2(n8582), .B1(n8583), .B2(n8584), .Y(n4457) );
	inv_1 U8486( .A(n7379), .Y(n8584) );
	nor2_1 U8487( .A(n8585), .B(n8586), .Y(n8583) );
	o22ai_1 U8488( .A1(n8582), .A2(n8587), .B1(n8588), .B2(n8589), .Y(n4456) );
	inv_1 U8489( .A(n7380), .Y(n8589) );
	nor2_1 U8490( .A(n8585), .B(n8590), .Y(n8588) );
	o22ai_1 U8491( .A1(n8582), .A2(n8591), .B1(n8592), .B2(n8593), .Y(n4455) );
	nor2_1 U8492( .A(n8585), .B(n8594), .Y(n8592) );
	and2_0 U8493( .A(n8595), .B(n5765), .X(n8585) );
	nand2_1 U8494( .A(n7266), .B(n8595), .Y(n8582) );
	or3_1 U8495( .A(n8596), .B(n8597), .C(n8598), .X(n8595) );
	o22ai_1 U8496( .A1(n8581), .A2(n8599), .B1(n8600), .B2(n8601), .Y(n4454) );
	nor2_1 U8497( .A(n8602), .B(n8586), .Y(n8600) );
	o22ai_1 U8498( .A1(n8587), .A2(n8599), .B1(n8603), .B2(n8604), .Y(n4453) );
	nor2_1 U8499( .A(n8602), .B(n8590), .Y(n8603) );
	o22ai_1 U8500( .A1(n8591), .A2(n8599), .B1(n8605), .B2(n8606), .Y(n4452) );
	inv_1 U8501( .A(n7729), .Y(n8606) );
	nor2_1 U8502( .A(n8602), .B(n8594), .Y(n8605) );
	a21oi_1 U8503( .A1(n8607), .A2(n8608), .B1(RST), .Y(n8602) );
	inv_1 U8504( .A(n8609), .Y(n8607) );
	o21ai_0 U8505( .A1(n8609), .A2(n8596), .B1(n8610), .Y(n8599) );
	mux2i_1 U8506( .A0(n8598), .A1(n8611), .S(n8544), .Y(n8610) );
	a21oi_1 U8507( .A1(n8612), .A2(n7266), .B1(n8613), .Y(n8609) );
	and4_1 U8508( .A(n8614), .B(n8615), .C(n8616), .D(n8617), .X(n8613) );
	o22ai_1 U8509( .A1(n8618), .A2(n8619), .B1(n8581), .B2(n8620), .Y(n4451) );
	o22ai_1 U8510( .A1(n8621), .A2(n8622), .B1(n8587), .B2(n8620), .Y(n4450) );
	inv_1 U8511( .A(n7472), .Y(n8622) );
	o22ai_1 U8512( .A1(n8623), .A2(n5629), .B1(n8591), .B2(n8620), .Y(n4449) );
	nand2_1 U8513( .A(n8624), .B(n8625), .Y(n8620) );
	mux2i_1 U8514( .A0(n8626), .A1(n8627), .S(n8628), .Y(n8624) );
	nand2_1 U8515( .A(n8617), .B(n8627), .Y(n8626) );
	o211ai_1 U8516( .A1(n8614), .A2(n8629), .B1(n8617), .C1(n8630), .Y(n8627) );
	mux2i_1 U8517( .A0(n8631), .A1(n8632), .S(n8633), .Y(n8630) );
	a21oi_1 U8518( .A1(n8634), .A2(n8635), .B1(n8636), .Y(n8632) );
	nand2_1 U8519( .A(n8614), .B(n8616), .Y(n8635) );
	nand3_1 U8520( .A(n8614), .B(n8615), .C(n7266), .Y(n8631) );
	inv_1 U8521( .A(n8611), .Y(n8629) );
	nand2_1 U8522( .A(n8634), .B(n8616), .Y(n8611) );
	o22ai_1 U8523( .A1(n8618), .A2(n8637), .B1(n8581), .B2(n8638), .Y(n4448) );
	o22ai_1 U8524( .A1(n8621), .A2(n8639), .B1(n8587), .B2(n8638), .Y(n4447) );
	inv_1 U8525( .A(n7474), .Y(n8639) );
	o22ai_1 U8526( .A1(n8623), .A2(n5630), .B1(n8591), .B2(n8638), .Y(n4446) );
	nand2_1 U8527( .A(n8640), .B(n8625), .Y(n8638) );
	xnor2_1 U8528( .A(n8641), .B(n8642), .Y(n8640) );
	a21oi_1 U8529( .A1(n8643), .A2(n8617), .B1(n8554), .Y(n8642) );
	o22ai_1 U8530( .A1(n8644), .A2(n8645), .B1(n8646), .B2(n8633), .Y(n8643) );
	a21oi_1 U8531( .A1(n8647), .A2(n8608), .B1(n8636), .Y(n8646) );
	a21oi_1 U8532( .A1(n8648), .A2(n8614), .B1(n8649), .Y(n8647) );
	mux2i_1 U8533( .A0(n8650), .A1(n8651), .S(n8633), .Y(n8645) );
	o21ai_0 U8534( .A1(n8628), .A2(n8652), .B1(n8653), .Y(n8651) );
	and2_0 U8535( .A(n8652), .B(n8614), .X(n8650) );
	nand2_1 U8536( .A(n8654), .B(n8616), .Y(n8652) );
	nand4_1 U8537( .A(n8655), .B(n8656), .C(n8657), .D(n8658), .Y(n8616) );
	nor3_1 U8538( .A(n8659), .B(n8660), .C(n8661), .Y(n8658) );
	or3_1 U8539( .A(n8662), .B(n8663), .C(n8664), .X(n8659) );
	nor3_1 U8540( .A(n8665), .B(n8666), .C(n8667), .Y(n8657) );
	o22ai_1 U8541( .A1(n8618), .A2(n8668), .B1(n8581), .B2(n8669), .Y(n4445) );
	o22ai_1 U8542( .A1(n8621), .A2(n8670), .B1(n8587), .B2(n8669), .Y(n4444) );
	inv_1 U8543( .A(n7470), .Y(n8670) );
	o22ai_1 U8544( .A1(n8623), .A2(n5631), .B1(n8591), .B2(n8669), .Y(n4443) );
	o21ai_0 U8545( .A1(n8671), .A2(n8672), .B1(n8625), .Y(n8669) );
	nor3_1 U8546( .A(n8615), .B(n8673), .C(n8612), .Y(n8672) );
	o22ai_1 U8547( .A1(n8581), .A2(n8674), .B1(n8675), .B2(n8676), .Y(n4442) );
	inv_1 U8548( .A(n7313), .Y(n8676) );
	nor2_1 U8549( .A(n8677), .B(n8586), .Y(n8675) );
	o22ai_1 U8550( .A1(n8587), .A2(n8674), .B1(n8678), .B2(n8679), .Y(n4441) );
	inv_1 U8551( .A(n7314), .Y(n8679) );
	nor2_1 U8552( .A(n8677), .B(n8590), .Y(n8678) );
	o22ai_1 U8553( .A1(n8591), .A2(n8674), .B1(n8680), .B2(n8681), .Y(n4440) );
	nor2_1 U8554( .A(n8677), .B(n8594), .Y(n8680) );
	a21oi_1 U8555( .A1(n8682), .A2(n8683), .B1(RST), .Y(n8677) );
	inv_1 U8556( .A(n8684), .Y(n8683) );
	o211ai_1 U8557( .A1(n8546), .A2(n8685), .B1(n7266), .C1(n8686), .Y(n8674) );
	mux2i_1 U8558( .A0(n8546), .A1(n8685), .S(n8687), .Y(n8686) );
	o22ai_1 U8559( .A1(n5552), .A2(n8618), .B1(n8581), .B2(n8688), .Y(n4439) );
	o22ai_1 U8560( .A1(n5342), .A2(n8621), .B1(n8587), .B2(n8688), .Y(n4438) );
	o22ai_1 U8561( .A1(n8689), .A2(n8623), .B1(n8591), .B2(n8688), .Y(n4437) );
	xnor2_1 U8562( .A(n8690), .B(n8546), .Y(n8688) );
	inv_1 U8563( .A(n8691), .Y(n8546) );
	nand2_1 U8564( .A(n8682), .B(n8684), .Y(n8690) );
	o221ai_1 U8565( .A1(n7314), .A2(n8692), .B1(n7313), .B2(n8693), .C1(n8694), .Y(n8684) );
	nand2_1 U8566( .A(g5437), .B(n8681), .Y(n8694) );
	inv_1 U8567( .A(n7715), .Y(n8681) );
	and2_0 U8568( .A(n8695), .B(n7266), .X(n8682) );
	mux2i_1 U8569( .A0(n8696), .A1(n8697), .S(n8687), .Y(n8695) );
	nand2_1 U8570( .A(n8685), .B(n8691), .Y(n8697) );
	or2_0 U8571( .A(n8691), .B(n8685), .X(n8696) );
	o221ai_1 U8572( .A1(n8692), .A2(n5342), .B1(n8693), .B2(n5552), .C1(n8698), .Y(n8691) );
	nand2_1 U8573( .A(n7635), .B(g5437), .Y(n8698) );
	inv_1 U8574( .A(n7635), .Y(n8689) );
	o22ai_1 U8575( .A1(n8618), .A2(n5632), .B1(n8581), .B2(n8699), .Y(n4436) );
	o22ai_1 U8576( .A1(n8621), .A2(n5381), .B1(n8587), .B2(n8699), .Y(n4435) );
	o22ai_1 U8577( .A1(n8623), .A2(n8700), .B1(n8591), .B2(n8699), .Y(n4434) );
	mux2_1 U8578( .A0(n8687), .A1(n8685), .S(n7266), .X(n8699) );
	o21ai_0 U8579( .A1(n8701), .A2(n8702), .B1(n8703), .Y(n8685) );
	inv_1 U8580( .A(n8704), .Y(n8703) );
	o22ai_1 U8581( .A1(n9978), .A2(n8705), .B1(n7390), .B2(n8706), .Y(n8702) );
	nor2_1 U8582( .A(n7393), .B(n8707), .Y(n8701) );
	a21oi_1 U8583( .A1(n7784), .A2(n10023), .B1(n8708), .Y(n8687) );
	o22ai_1 U8584( .A1(n8700), .A2(n8709), .B1(n5381), .B2(n8692), .Y(n8708) );
	inv_1 U8585( .A(n7631), .Y(n8700) );
	o22ai_1 U8586( .A1(n8581), .A2(n8710), .B1(n8711), .B2(n8712), .Y(n4433) );
	inv_1 U8587( .A(n7341), .Y(n8712) );
	nor2_1 U8588( .A(n8713), .B(n8586), .Y(n8711) );
	o22ai_1 U8589( .A1(n8587), .A2(n8710), .B1(n8714), .B2(n8715), .Y(n4432) );
	inv_1 U8590( .A(n7342), .Y(n8715) );
	nor2_1 U8591( .A(n8713), .B(n8590), .Y(n8714) );
	o22ai_1 U8592( .A1(n8591), .A2(n8710), .B1(n8716), .B2(n8717), .Y(n4431) );
	nor2_1 U8593( .A(n8713), .B(n8594), .Y(n8716) );
	a21oi_1 U8594( .A1(n8718), .A2(n8719), .B1(RST), .Y(n8713) );
	o22ai_1 U8595( .A1(n5553), .A2(n8618), .B1(n8720), .B2(n8581), .Y(n4430) );
	o22ai_1 U8596( .A1(n5343), .A2(n8621), .B1(n8720), .B2(n8587), .Y(n4429) );
	o22ai_1 U8597( .A1(n8721), .A2(n8623), .B1(n8720), .B2(n8591), .Y(n4428) );
	xnor2_1 U8598( .A(n8580), .B(n8722), .Y(n8720) );
	a21oi_1 U8599( .A1(n8636), .A2(n8723), .B1(n8724), .Y(n8722) );
	nor4_1 U8600( .A(n8725), .B(n8719), .C(n8598), .D(n8726), .Y(n8724) );
	inv_1 U8601( .A(n8727), .Y(n8719) );
	inv_1 U8602( .A(n7622), .Y(n8721) );
	o22ai_1 U8603( .A1(n8728), .A2(n8581), .B1(n8618), .B2(n5673), .Y(n4427) );
	inv_1 U8604( .A(n8586), .Y(n8618) );
	nor2_1 U8605( .A(n7784), .B(RST), .Y(n8586) );
	nand2_1 U8606( .A(n7784), .B(n5747), .Y(n8581) );
	o22ai_1 U8607( .A1(n8621), .A2(n5634), .B1(n8728), .B2(n8587), .Y(n4426) );
	inv_1 U8608( .A(n100), .Y(n8587) );
	inv_1 U8609( .A(n8590), .Y(n8621) );
	nor2_1 U8610( .A(g6447), .B(RST), .Y(n8590) );
	o22ai_1 U8611( .A1(n8728), .A2(n8591), .B1(n8623), .B2(n8729), .Y(n4425) );
	inv_1 U8612( .A(n8594), .Y(n8623) );
	nor2_1 U8613( .A(g5437), .B(RST), .Y(n8594) );
	inv_1 U8614( .A(n3958), .Y(n8591) );
	xnor2_1 U8615( .A(n8725), .B(n8730), .Y(n8728) );
	a21oi_1 U8616( .A1(n8731), .A2(n7266), .B1(n8732), .Y(n8730) );
	inv_1 U8617( .A(n8710), .Y(n8732) );
	nand2_1 U8618( .A(n8725), .B(n8718), .Y(n8710) );
	o32ai_1 U8619( .A1(n8598), .A2(n8580), .A3(n8733), .B1(n8636), .B2(n8734), .Y(n8718) );
	inv_1 U8620( .A(n8723), .Y(n8734) );
	nor3_1 U8621( .A(n8598), .B(n8536), .C(n8735), .Y(n8723) );
	inv_1 U8622( .A(n8733), .Y(n8735) );
	inv_1 U8623( .A(n7266), .Y(n8598) );
	a21oi_1 U8624( .A1(n8736), .A2(n8737), .B1(n8725), .Y(n8731) );
	inv_1 U8625( .A(n8726), .Y(n8737) );
	xnor2_1 U8626( .A(n8733), .B(n8536), .Y(n8726) );
	nor3_1 U8627( .A(n8738), .B(n8739), .C(n8704), .Y(n8733) );
	a21oi_1 U8628( .A1(n8636), .A2(n8580), .B1(n8727), .Y(n8736) );
	o221ai_1 U8629( .A1(n7342), .A2(n8692), .B1(n7341), .B2(n8693), .C1(n8740), .Y(n8727) );
	nand2_1 U8630( .A(g5437), .B(n8717), .Y(n8740) );
	inv_1 U8631( .A(n7735), .Y(n8717) );
	inv_1 U8632( .A(n8536), .Y(n8580) );
	o221ai_1 U8633( .A1(n8692), .A2(n5343), .B1(n8693), .B2(n5553), .C1(n8741), .Y(n8536) );
	nand2_1 U8634( .A(n7622), .B(g5437), .Y(n8741) );
	a221oi_1 U8635( .A1(g6447), .A2(n9839), .B1(n7784), .B2(n10024), .C1(n8742), .Y(n8725) );
	nor2_1 U8636( .A(n8729), .B(n8709), .Y(n8742) );
	inv_1 U8637( .A(n7627), .Y(n8729) );
	and2_0 U8638( .A(g5549), .B(n5765), .X(n4424) );
	nor2_1 U8639( .A(n8743), .B(n8744), .Y(n4423) );
	xnor2_1 U8640( .A(n10025), .B(n8745), .Y(n8743) );
	nor2_1 U8641( .A(n8746), .B(n8747), .Y(n8745) );
	nor2_1 U8642( .A(n8748), .B(n8744), .Y(n4422) );
	xnor2_1 U8643( .A(n8747), .B(n8746), .Y(n8748) );
	inv_1 U8644( .A(n7306), .Y(n8746) );
	nand2_1 U8645( .A(n8749), .B(n7708), .Y(n8747) );
	nor2_1 U8646( .A(n8750), .B(n8744), .Y(n4421) );
	xnor2_1 U8647( .A(n7708), .B(n8749), .Y(n8750) );
	a211oi_1 U8648( .A1(n5373), .A2(n8751), .B1(n8744), .C1(n8749), .Y(n4420) );
	nor2_1 U8649( .A(n8751), .B(n5373), .Y(n8749) );
	nor3_1 U8650( .A(n8744), .B(n8752), .C(n8753), .Y(n4419) );
	a21oi_1 U8651( .A1(n8754), .A2(n10027), .B1(n7304), .Y(n8753) );
	inv_1 U8652( .A(n8751), .Y(n8752) );
	nand3_1 U8653( .A(n7304), .B(n10027), .C(n8754), .Y(n8751) );
	nor2_1 U8654( .A(n8755), .B(n8744), .Y(n4418) );
	xnor2_1 U8655( .A(n10027), .B(n8754), .Y(n8755) );
	a211oi_1 U8656( .A1(n8756), .A2(n8757), .B1(n8744), .C1(n8754), .Y(n4417) );
	nor2_1 U8657( .A(n8757), .B(n8756), .Y(n8754) );
	inv_1 U8658( .A(n8758), .Y(n8757) );
	inv_1 U8659( .A(n7712), .Y(n8756) );
	a211oi_1 U8660( .A1(n5374), .A2(n8759), .B1(n8744), .C1(n8758), .Y(n4416) );
	nor2_1 U8661( .A(n8759), .B(n5374), .Y(n8758) );
	nor3_1 U8662( .A(n8744), .B(n8760), .C(n8761), .Y(n4415) );
	a21oi_1 U8663( .A1(n8762), .A2(n10029), .B1(n7702), .Y(n8761) );
	inv_1 U8664( .A(n8759), .Y(n8760) );
	nand3_1 U8665( .A(n7702), .B(n10029), .C(n8762), .Y(n8759) );
	nor2_1 U8666( .A(n8763), .B(n8744), .Y(n4414) );
	o21ai_0 U8667( .A1(n6131), .A2(n8764), .B1(n5742), .Y(n8744) );
	xnor2_1 U8668( .A(n8762), .B(n10029), .Y(n8763) );
	nor2_1 U8669( .A(n8705), .B(n6337), .Y(n8762) );
	o22ai_1 U8670( .A1(n8765), .A2(n8766), .B1(n8767), .B2(n8768), .Y(n4413) );
	o22ai_1 U8671( .A1(n5731), .A2(n8769), .B1(n8767), .B2(n8770), .Y(n4412) );
	o22ai_1 U8672( .A1(n5687), .A2(n8771), .B1(n8767), .B2(n8772), .Y(n4411) );
	o221ai_1 U8673( .A1(n8773), .A2(n8774), .B1(n8775), .B2(n8776), .C1(n8777), .Y(n8767) );
	xnor2_1 U8674( .A(n8778), .B(n8565), .Y(n8773) );
	nand2_1 U8675( .A(n8779), .B(n8780), .Y(n8778) );
	xnor2_1 U8676( .A(n8570), .B(n8781), .Y(n8780) );
	o22ai_1 U8677( .A1(n8782), .A2(n8766), .B1(n8783), .B2(n8768), .Y(n4410) );
	o22ai_1 U8678( .A1(n5527), .A2(n8769), .B1(n8783), .B2(n8770), .Y(n4409) );
	o22ai_1 U8679( .A1(n5713), .A2(n8771), .B1(n8783), .B2(n8772), .Y(n4408) );
	inv_1 U8680( .A(n8784), .Y(n8783) );
	o221ai_1 U8681( .A1(n8774), .A2(n8785), .B1(n8671), .B2(n8786), .C1(n8787), .Y(n8784) );
	nand2_1 U8682( .A(n8788), .B(n8789), .Y(n8787) );
	xnor2_1 U8683( .A(n8790), .B(n8779), .Y(n8785) );
	nor2_1 U8684( .A(n8791), .B(n8792), .Y(n8779) );
	xnor2_1 U8685( .A(n8562), .B(n8781), .Y(n8792) );
	o22ai_1 U8686( .A1(n8793), .A2(n8766), .B1(n8768), .B2(n8794), .Y(n4407) );
	o22ai_1 U8687( .A1(n5732), .A2(n8769), .B1(n8770), .B2(n8794), .Y(n4406) );
	o22ai_1 U8688( .A1(n5688), .A2(n8771), .B1(n8772), .B2(n8794), .Y(n4405) );
	nand2_1 U8689( .A(n8795), .B(n8786), .Y(n8794) );
	mux2i_1 U8690( .A0(n8796), .A1(n8797), .S(n8774), .Y(n8795) );
	xor2_1 U8691( .A(n8791), .B(n8562), .X(n8796) );
	nand2_1 U8692( .A(n8798), .B(n8799), .Y(n8791) );
	xnor2_1 U8693( .A(n8576), .B(n8671), .Y(n8799) );
	o22ai_1 U8694( .A1(n8800), .A2(n8766), .B1(n8801), .B2(n8768), .Y(n4404) );
	o22ai_1 U8695( .A1(n5733), .A2(n8769), .B1(n8801), .B2(n8770), .Y(n4403) );
	o22ai_1 U8696( .A1(n5689), .A2(n8771), .B1(n8801), .B2(n8772), .Y(tempn4402) );
	inv_1 U8697( .A(n8802), .Y(n8801) );
	o22ai_1 U8698( .A1(n8803), .A2(n8776), .B1(n8774), .B2(n8804), .Y(n8802) );
	xnor2_1 U8699( .A(n8576), .B(n8798), .Y(n8804) );
	nor2_1 U8700( .A(n8805), .B(n8806), .Y(n8798) );
	xnor2_1 U8701( .A(n8578), .B(n8781), .Y(n8806) );
	o22ai_1 U8702( .A1(n8807), .A2(n8766), .B1(n8768), .B2(n8808), .Y(n4401) );
	o22ai_1 U8703( .A1(n5734), .A2(n8769), .B1(n8770), .B2(n8808), .Y(n4400) );
	o22ai_1 U8704( .A1(n5690), .A2(n8771), .B1(n8772), .B2(n8808), .Y(n4399) );
	nand2_1 U8705( .A(n8809), .B(n8786), .Y(n8808) );
	mux2i_1 U8706( .A0(n8810), .A1(n8811), .S(n8774), .Y(n8809) );
	xor2_1 U8707( .A(n8805), .B(n8578), .X(n8810) );
	nand2_1 U8708( .A(n8812), .B(n8813), .Y(n8805) );
	xnor2_1 U8709( .A(n8814), .B(n8781), .Y(n8813) );
	o22ai_1 U8710( .A1(n8815), .A2(n8766), .B1(n8816), .B2(n8768), .Y(n4398) );
	o22ai_1 U8711( .A1(n5735), .A2(n8769), .B1(n8816), .B2(n8770), .Y(n4397) );
	o22ai_1 U8712( .A1(n5691), .A2(n8771), .B1(n8816), .B2(n8772), .Y(n4396) );
	inv_1 U8713( .A(n8817), .Y(n8816) );
	o22ai_1 U8714( .A1(n8818), .A2(n8776), .B1(n8774), .B2(n8819), .Y(n8817) );
	xnor2_1 U8715( .A(n8577), .B(n8812), .Y(n8819) );
	nor2_1 U8716( .A(n8820), .B(n8821), .Y(n8812) );
	xnor2_1 U8717( .A(n8822), .B(n8781), .Y(n8821) );
	o22ai_1 U8718( .A1(n8823), .A2(n8766), .B1(n8768), .B2(n8824), .Y(n4395) );
	o22ai_1 U8719( .A1(n5526), .A2(n8769), .B1(n8770), .B2(n8824), .Y(n4394) );
	o22ai_1 U8720( .A1(n5714), .A2(n8771), .B1(n8772), .B2(n8824), .Y(n4393) );
	o221ai_1 U8721( .A1(n8825), .A2(n8774), .B1(n7282), .B2(n8776), .C1(n8777), .Y(n8824) );
	xnor2_1 U8722( .A(n8820), .B(n8822), .Y(n8825) );
	nand2_1 U8723( .A(n8826), .B(n8827), .Y(n8820) );
	xnor2_1 U8724( .A(n8572), .B(n8781), .Y(n8827) );
	o22ai_1 U8725( .A1(n8828), .A2(n8766), .B1(n8829), .B2(n8768), .Y(n4392) );
	o22ai_1 U8726( .A1(n5528), .A2(n8769), .B1(n8829), .B2(n8770), .Y(n4391) );
	o22ai_1 U8727( .A1(n5715), .A2(n8771), .B1(n8829), .B2(n8772), .Y(n4390) );
	inv_1 U8728( .A(n8830), .Y(n8829) );
	o221ai_1 U8729( .A1(n8774), .A2(n8831), .B1(n8671), .B2(n8786), .C1(n8832), .Y(n8830) );
	nand2_1 U8730( .A(n8788), .B(n7233), .Y(n8832) );
	inv_1 U8731( .A(n8776), .Y(n8788) );
	xnor2_1 U8732( .A(n8833), .B(n8826), .Y(n8831) );
	nor2_1 U8733( .A(n8834), .B(n8835), .Y(n8826) );
	xnor2_1 U8734( .A(n8836), .B(n8781), .Y(n8835) );
	o22ai_1 U8735( .A1(n8837), .A2(n8766), .B1(n8768), .B2(n8838), .Y(n4389) );
	o22ai_1 U8736( .A1(n5529), .A2(n8769), .B1(n8770), .B2(n8838), .Y(n4388) );
	o22ai_1 U8737( .A1(n5716), .A2(n8771), .B1(n8772), .B2(n8838), .Y(n4387) );
	o221ai_1 U8738( .A1(n8839), .A2(n8774), .B1(n7252), .B2(n8776), .C1(n8777), .Y(n8838) );
	or2_0 U8739( .A(n8786), .B(n8781), .X(n8777) );
	xnor2_1 U8740( .A(n8834), .B(n8836), .Y(n8839) );
	nand2_1 U8741( .A(n8840), .B(n8841), .Y(n8834) );
	xnor2_1 U8742( .A(n8561), .B(n8671), .Y(n8840) );
	o22ai_1 U8743( .A1(n8842), .A2(n8768), .B1(n8843), .B2(n8766), .Y(n4386) );
	nand2_1 U8744( .A(n8705), .B(n5747), .Y(n8766) );
	nand2_1 U8745( .A(n7230), .B(n5747), .Y(n8768) );
	o22ai_1 U8746( .A1(n5736), .A2(n8769), .B1(n8842), .B2(n8770), .Y(n4385) );
	inv_1 U8747( .A(n91), .Y(n8770) );
	nor2_1 U8748( .A(n8706), .B(RST), .Y(n91) );
	nand2_1 U8749( .A(n8706), .B(n5747), .Y(n8769) );
	o22ai_1 U8750( .A1(n5692), .A2(n8771), .B1(n8842), .B2(n8772), .Y(n4384) );
	inv_1 U8751( .A(n90), .Y(n8772) );
	nor2_1 U8752( .A(n8707), .B(RST), .Y(n90) );
	inv_1 U8753( .A(n8844), .Y(n8842) );
	o22ai_1 U8754( .A1(n8845), .A2(n8776), .B1(n8846), .B2(n8774), .Y(n8844) );
	xnor2_1 U8755( .A(n8841), .B(n8561), .Y(n8846) );
	nand2_1 U8756( .A(n8786), .B(n8774), .Y(n8776) );
	o221ai_1 U8757( .A1(n8847), .A2(n8848), .B1(n8673), .B2(n8849), .C1(n8850), .Y(n8774) );
	a21oi_1 U8758( .A1(n8851), .A2(n8608), .B1(n8852), .Y(n8850) );
	inv_1 U8759( .A(n8625), .Y(n8852) );
	a21oi_1 U8760( .A1(n8544), .A2(n8853), .B1(n8649), .Y(n8851) );
	a221oi_1 U8761( .A1(n8604), .A2(g6447), .B1(n8601), .B2(n7784), .C1(n8854), .Y(n8649) );
	nor2_1 U8762( .A(n8709), .B(n7729), .Y(n8854) );
	inv_1 U8763( .A(n7332), .Y(n8601) );
	inv_1 U8764( .A(n7334), .Y(n8604) );
	nand3_1 U8765( .A(n8615), .B(n8617), .C(n8641), .Y(n8853) );
	inv_1 U8766( .A(n8648), .Y(n8615) );
	a21oi_1 U8767( .A1(n8653), .A2(n8654), .B1(n8644), .Y(n8648) );
	inv_1 U8768( .A(n8855), .Y(n8654) );
	o221ai_1 U8769( .A1(n8856), .A2(n8857), .B1(n8858), .B2(n8859), .C1(n8860), .Y(n8855) );
	o221ai_1 U8770( .A1(n8666), .A2(n8861), .B1(n8667), .B2(n8665), .C1(n8661), .Y(n8860) );
	o22ai_1 U8771( .A1(n8666), .A2(n8665), .B1(n8861), .B2(n8661), .Y(n8859) );
	inv_1 U8772( .A(n8856), .Y(n8666) );
	o22ai_1 U8773( .A1(n8667), .A2(n8861), .B1(n8665), .B2(n8661), .Y(n8857) );
	xnor2_1 U8774( .A(n8775), .B(n8862), .Y(n8661) );
	inv_1 U8775( .A(n8565), .Y(n8862) );
	xnor2_1 U8776( .A(n8562), .B(n8797), .Y(n8665) );
	inv_1 U8777( .A(n8656), .Y(n8861) );
	xnor2_1 U8778( .A(n7282), .B(n8822), .Y(n8656) );
	inv_1 U8779( .A(n8858), .Y(n8667) );
	xor2_1 U8780( .A(n8578), .B(n8811), .X(n8858) );
	xnor2_1 U8781( .A(n7252), .B(n8836), .Y(n8856) );
	inv_1 U8782( .A(n8863), .Y(n8653) );
	o221ai_1 U8783( .A1(n8864), .A2(n8865), .B1(n8866), .B2(n8867), .C1(n8868), .Y(n8863) );
	o221ai_1 U8784( .A1(n8869), .A2(n8660), .B1(n8663), .B2(n8662), .C1(n8664), .Y(n8868) );
	o22ai_1 U8785( .A1(n8869), .A2(n8664), .B1(n8663), .B2(n8660), .Y(n8867) );
	o22ai_1 U8786( .A1(n8869), .A2(n8662), .B1(n8663), .B2(n8664), .Y(n8865) );
	xnor2_1 U8787( .A(n8561), .B(n8845), .Y(n8664) );
	xor2_1 U8788( .A(n8870), .B(n8572), .X(n8663) );
	inv_1 U8789( .A(n8866), .Y(n8662) );
	xnor2_1 U8790( .A(n8814), .B(n8818), .Y(n8866) );
	inv_1 U8791( .A(n8577), .Y(n8814) );
	inv_1 U8792( .A(n8655), .Y(n8869) );
	xor2_1 U8793( .A(n8576), .B(n8803), .X(n8655) );
	inv_1 U8794( .A(n8660), .Y(n8864) );
	xnor2_1 U8795( .A(n8739), .B(n8790), .Y(n8660) );
	inv_1 U8796( .A(n8612), .Y(n8544) );
	nor3_1 U8797( .A(n8673), .B(n8614), .C(n8633), .Y(n8612) );
	inv_1 U8798( .A(n8628), .Y(n8614) );
	inv_1 U8799( .A(n8636), .Y(n8849) );
	nor2_1 U8800( .A(n8871), .B(n8872), .Y(n8636) );
	inv_1 U8801( .A(n7719), .Y(n8872) );
	a21oi_1 U8802( .A1(n8555), .A2(n8781), .B1(n8873), .Y(n8848) );
	inv_1 U8803( .A(n8671), .Y(n8781) );
	o211ai_1 U8804( .A1(n8555), .A2(n8873), .B1(n8841), .C1(n8625), .Y(n8786) );
	nand2_1 U8805( .A(n8608), .B(n8597), .Y(n8625) );
	o221ai_1 U8806( .A1(n7380), .A2(n8692), .B1(n7379), .B2(n8693), .C1(n8874), .Y(n8597) );
	nand2_1 U8807( .A(g5437), .B(n8593), .Y(n8874) );
	inv_1 U8808( .A(n7740), .Y(n8593) );
	inv_1 U8809( .A(n8596), .Y(n8608) );
	nand2_1 U8810( .A(n8875), .B(n8876), .Y(n8596) );
	nor4_1 U8811( .A(n8877), .B(n8878), .C(n8879), .D(n8880), .Y(n8876) );
	xnor2_1 U8812( .A(n8881), .B(n8775), .Y(n8880) );
	a222oi_1 U8813( .A1(g6313), .A2(n8882), .B1(n7230), .B2(n5434), .C1(g6231), .C2(n8883), .Y(n8881) );
	xnor2_1 U8814( .A(n8884), .B(n8789), .Y(n8879) );
	a222oi_1 U8815( .A1(g6313), .A2(n8885), .B1(n7230), .B2(n5435), .C1(g6231), .C2(n8886), .Y(n8884) );
	mux2i_1 U8816( .A0(n8887), .A1(n8888), .S(n8811), .Y(n8878) );
	nand2_1 U8817( .A(n10030), .B(n8888), .Y(n8887) );
	nand3_1 U8818( .A(n8889), .B(n8890), .C(n8634), .Y(n8877) );
	inv_1 U8819( .A(n8644), .Y(n8634) );
	nand2_1 U8820( .A(n7719), .B(n8871), .Y(n8644) );
	o21ai_0 U8821( .A1(n10031), .A2(n8705), .B1(n8891), .Y(n8871) );
	a22oi_1 U8822( .A1(g6231), .A2(n8892), .B1(g6313), .B2(n8893), .Y(n8891) );
	xnor2_1 U8823( .A(n8894), .B(n8895), .Y(n8890) );
	a222oi_1 U8824( .A1(g6313), .A2(n8896), .B1(n7230), .B2(n5436), .C1(g6231), .C2(n8897), .Y(n8895) );
	xnor2_1 U8825( .A(n8845), .B(n8898), .Y(n8889) );
	a222oi_1 U8826( .A1(g6313), .A2(n8899), .B1(n7230), .B2(n5442), .C1(g6231), .C2(n8900), .Y(n8898) );
	nor4_1 U8827( .A(n8901), .B(n8902), .C(n8903), .D(n8904), .Y(n8875) );
	mux2i_1 U8828( .A0(n8905), .A1(n8906), .S(n8907), .Y(n8904) );
	nand2_1 U8829( .A(n7616), .B(n8906), .Y(n8905) );
	mux2i_1 U8830( .A0(n8908), .A1(n8909), .S(n8803), .Y(n8903) );
	nand2_1 U8831( .A(n7613), .B(n8909), .Y(n8908) );
	mux2i_1 U8832( .A0(n8910), .A1(n8911), .S(n8797), .Y(n8902) );
	nand2_1 U8833( .A(n7286), .B(n8911), .Y(n8910) );
	nand3_1 U8834( .A(n8912), .B(n8913), .C(n8914), .Y(n8901) );
	mux2i_1 U8835( .A0(n8915), .A1(n8916), .S(n8870), .Y(n8914) );
	nor2_1 U8836( .A(n8916), .B(n5358), .Y(n8915) );
	mux2i_1 U8837( .A0(n8917), .A1(n8918), .S(n8705), .Y(n8913) );
	nand2_1 U8838( .A(n8919), .B(n8920), .Y(n8918) );
	a222oi_1 U8839( .A1(n7223), .A2(n8911), .B1(n7269), .B2(n8888), .C1(n7282), .C2(n8906), .Y(n8920) );
	a22oi_1 U8840( .A1(n5499), .A2(g6313), .B1(n5330), .B2(g6231), .Y(n8906) );
	a22oi_1 U8841( .A1(n5498), .A2(g6313), .B1(n5329), .B2(g6231), .Y(n8888) );
	a22oi_1 U8842( .A1(n5496), .A2(g6313), .B1(n5327), .B2(g6231), .Y(n8911) );
	a222oi_1 U8843( .A1(n7233), .A2(n8921), .B1(n7241), .B2(n8909), .C1(n7244), .C2(n8922), .Y(n8919) );
	inv_1 U8844( .A(n8923), .Y(n8922) );
	a22oi_1 U8845( .A1(n5497), .A2(g6313), .B1(n5328), .B2(g6231), .Y(n8909) );
	inv_1 U8846( .A(n8916), .Y(n8921) );
	o22ai_1 U8847( .A1(n9861), .A2(n8706), .B1(n9862), .B2(n8707), .Y(n8916) );
	nand2_1 U8848( .A(n8924), .B(n8925), .Y(n8917) );
	a222oi_1 U8849( .A1(n8803), .A2(n8926), .B1(n8797), .B2(n8927), .C1(n8870), .C2(n5358), .Y(n8925) );
	a222oi_1 U8850( .A1(n8907), .A2(n8928), .B1(n8818), .B2(n8929), .C1(n8811), .C2(n5376), .Y(n8924) );
	mux2i_1 U8851( .A0(n8930), .A1(n8923), .S(n8818), .Y(n8912) );
	nor2_1 U8852( .A(n8923), .B(n8929), .Y(n8930) );
	o22ai_1 U8853( .A1(n9859), .A2(n8706), .B1(n9860), .B2(n8707), .Y(n8923) );
	inv_1 U8854( .A(n8847), .Y(n8841) );
	nor2_1 U8855( .A(n8554), .B(n8671), .Y(n8847) );
	and4_1 U8856( .A(n8931), .B(n8565), .C(n8671), .D(n8932), .X(n8873) );
	nor4_1 U8857( .A(n8571), .B(n8572), .C(n8570), .D(n8560), .Y(n8932) );
	inv_1 U8858( .A(n8822), .Y(n8560) );
	inv_1 U8859( .A(n8790), .Y(n8570) );
	nor3_1 U8860( .A(n8617), .B(n8641), .C(n8628), .Y(n8671) );
	inv_1 U8861( .A(n8633), .Y(n8641) );
	and4_1 U8862( .A(n8571), .B(n8572), .C(n8931), .D(n8933), .X(n8555) );
	nor3_1 U8863( .A(n8790), .B(n8565), .C(n8822), .Y(n8933) );
	o221ai_1 U8864( .A1(n8706), .A2(n5526), .B1(n8705), .B2(n8823), .C1(n8934), .Y(n8822) );
	nand2_1 U8865( .A(n9845), .B(g6231), .Y(n8934) );
	inv_1 U8866( .A(n7621), .Y(n8823) );
	o21ai_0 U8867( .A1(n8705), .A2(n8765), .B1(n8935), .Y(n8565) );
	a22oi_1 U8868( .A1(n9844), .A2(g6231), .B1(n9843), .B2(g6313), .Y(n8935) );
	inv_1 U8869( .A(n7654), .Y(n8765) );
	o221ai_1 U8870( .A1(n8706), .A2(n5527), .B1(n8705), .B2(n8782), .C1(n8936), .Y(n8790) );
	nand2_1 U8871( .A(n9856), .B(g6231), .Y(n8936) );
	inv_1 U8872( .A(n7657), .Y(n8782) );
	nor4_1 U8873( .A(n8577), .B(n8576), .C(n8937), .D(n8578), .Y(n8931) );
	o21ai_0 U8874( .A1(n8705), .A2(n8807), .B1(n8938), .Y(n8578) );
	a22oi_1 U8875( .A1(n9851), .A2(g6231), .B1(n9850), .B2(g6313), .Y(n8938) );
	inv_1 U8876( .A(n7649), .Y(n8807) );
	or2_0 U8877( .A(n8562), .B(n8561), .X(n8937) );
	o21ai_0 U8878( .A1(n8705), .A2(n8843), .B1(n8939), .Y(n8561) );
	a22oi_1 U8879( .A1(n9849), .A2(g6231), .B1(n9848), .B2(g6313), .Y(n8939) );
	inv_1 U8880( .A(n7651), .Y(n8843) );
	o21ai_0 U8881( .A1(n8705), .A2(n8793), .B1(n8940), .Y(n8562) );
	a22oi_1 U8882( .A1(n9847), .A2(g6231), .B1(n9846), .B2(g6313), .Y(n8940) );
	inv_1 U8883( .A(n7655), .Y(n8793) );
	o21ai_0 U8884( .A1(n8705), .A2(n8800), .B1(n8941), .Y(n8576) );
	a22oi_1 U8885( .A1(n9853), .A2(g6231), .B1(n9852), .B2(g6313), .Y(n8941) );
	inv_1 U8886( .A(n7650), .Y(n8800) );
	o21ai_0 U8887( .A1(n8705), .A2(n8815), .B1(n8942), .Y(n8577) );
	a22oi_1 U8888( .A1(n9855), .A2(g6231), .B1(n9854), .B2(g6313), .Y(n8942) );
	inv_1 U8889( .A(n7653), .Y(n8815) );
	inv_1 U8890( .A(n8833), .Y(n8572) );
	o221ai_1 U8891( .A1(n8706), .A2(n5528), .B1(n8705), .B2(n8828), .C1(n8943), .Y(n8833) );
	nand2_1 U8892( .A(n9857), .B(g6231), .Y(n8943) );
	inv_1 U8893( .A(n7656), .Y(n8828) );
	inv_1 U8894( .A(n8836), .Y(n8571) );
	o221ai_1 U8895( .A1(n8706), .A2(n5529), .B1(n8705), .B2(n8837), .C1(n8944), .Y(n8836) );
	nand2_1 U8896( .A(n9858), .B(g6231), .Y(n8944) );
	inv_1 U8897( .A(n7652), .Y(n8837) );
	inv_1 U8898( .A(g6313), .Y(n8706) );
	nand2_1 U8899( .A(n8707), .B(n5747), .Y(n8771) );
	inv_1 U8900( .A(g6231), .Y(n8707) );
	o22ai_1 U8901( .A1(n8945), .A2(n5604), .B1(n8946), .B2(n8947), .Y(n4383) );
	o22ai_1 U8902( .A1(n8948), .A2(n8949), .B1(n8947), .B2(n8950), .Y(n4382) );
	inv_1 U8903( .A(n7390), .Y(n8949) );
	o22ai_1 U8904( .A1(n8951), .A2(n8952), .B1(n8947), .B2(n8953), .Y(n4381) );
	nand2_1 U8905( .A(n8704), .B(n5747), .Y(n8947) );
	nand2_1 U8906( .A(n8954), .B(n8955), .Y(n8704) );
	nor4_1 U8907( .A(n8894), .B(n8845), .C(n8811), .D(n8803), .Y(n8955) );
	inv_1 U8908( .A(n7241), .Y(n8803) );
	inv_1 U8909( .A(n7594), .Y(n8845) );
	inv_1 U8910( .A(n7252), .Y(n8894) );
	nor4_1 U8911( .A(n8907), .B(n8797), .C(n8818), .D(n8870), .Y(n8954) );
	inv_1 U8912( .A(n7233), .Y(n8870) );
	inv_1 U8913( .A(n7244), .Y(n8818) );
	inv_1 U8914( .A(n7223), .Y(n8797) );
	inv_1 U8915( .A(n7282), .Y(n8907) );
	inv_1 U8916( .A(n7393), .Y(n8952) );
	o22ai_1 U8917( .A1(n8946), .A2(n8956), .B1(n8945), .B2(n8957), .Y(n4380) );
	inv_1 U8918( .A(n7445), .Y(n8957) );
	o22ai_1 U8919( .A1(n8950), .A2(n8956), .B1(n8948), .B2(n5413), .Y(n4379) );
	o22ai_1 U8920( .A1(n8953), .A2(n8956), .B1(n8951), .B2(n8958), .Y(n4378) );
	o22ai_1 U8921( .A1(n8946), .A2(n8959), .B1(n8945), .B2(n8960), .Y(n4377) );
	inv_1 U8922( .A(n7441), .Y(n8960) );
	o22ai_1 U8923( .A1(n8950), .A2(n8959), .B1(n8948), .B2(n8961), .Y(n4376) );
	o22ai_1 U8924( .A1(n8953), .A2(n8959), .B1(n8951), .B2(n5401), .Y(n4375) );
	o22ai_1 U8925( .A1(n8946), .A2(n8962), .B1(n8945), .B2(n5678), .Y(n4374) );
	nand2_1 U8926( .A(n8946), .B(n5747), .Y(n8945) );
	nand2_1 U8927( .A(n7230), .B(n6529), .Y(n8946) );
	o22ai_1 U8928( .A1(n8950), .A2(n8962), .B1(n8948), .B2(n8893), .Y(n4373) );
	inv_1 U8929( .A(n7397), .Y(n8893) );
	nand2_1 U8930( .A(n8950), .B(n5747), .Y(n8948) );
	nand2_1 U8931( .A(n6529), .B(g6313), .Y(n8950) );
	o22ai_1 U8932( .A1(n8953), .A2(n8962), .B1(n8951), .B2(n8892), .Y(n4372) );
	inv_1 U8933( .A(n7398), .Y(n8892) );
	nand2_1 U8934( .A(n8953), .B(n5747), .Y(n8951) );
	nand4_1 U8935( .A(n98), .B(n7244), .C(n7223), .D(n8811), .Y(n8962) );
	inv_1 U8936( .A(n7269), .Y(n8811) );
	nand2_1 U8937( .A(n6529), .B(g6231), .Y(n8953) );
	inv_1 U8938( .A(n8963), .Y(n6529) );
	o22ai_1 U8939( .A1(n8964), .A2(n5434), .B1(n8764), .B2(n8965), .Y(n4371) );
	o22ai_1 U8940( .A1(n8966), .A2(n8882), .B1(n8965), .B2(n8967), .Y(n4370) );
	inv_1 U8941( .A(n7433), .Y(n8882) );
	o22ai_1 U8942( .A1(n8968), .A2(n8883), .B1(n8965), .B2(n8969), .Y(n4369) );
	nand2_1 U8943( .A(n8738), .B(n5746), .Y(n8965) );
	inv_1 U8944( .A(n8775), .Y(n8738) );
	o21ai_0 U8945( .A1(n7441), .A2(n8705), .B1(n8970), .Y(n8775) );
	a22oi_1 U8946( .A1(g6231), .A2(n5401), .B1(g6313), .B2(n8961), .Y(n8970) );
	inv_1 U8947( .A(n7440), .Y(n8961) );
	inv_1 U8948( .A(n7439), .Y(n8883) );
	o22ai_1 U8949( .A1(n8964), .A2(n5435), .B1(n8764), .B2(n8971), .Y(n4368) );
	o22ai_1 U8950( .A1(n8966), .A2(n8885), .B1(n8967), .B2(n8971), .Y(n4367) );
	inv_1 U8951( .A(n7442), .Y(n8885) );
	o22ai_1 U8952( .A1(n8968), .A2(n8886), .B1(n8969), .B2(n8971), .Y(n4366) );
	nand2_1 U8953( .A(n8739), .B(n5744), .Y(n8971) );
	inv_1 U8954( .A(n8789), .Y(n8739) );
	o21ai_0 U8955( .A1(n7445), .A2(n8705), .B1(n8972), .Y(n8789) );
	a22oi_1 U8956( .A1(g6231), .A2(n8958), .B1(g6313), .B2(n5413), .Y(n8972) );
	inv_1 U8957( .A(n7446), .Y(n8958) );
	inv_1 U8958( .A(n7230), .Y(n8705) );
	inv_1 U8959( .A(n7444), .Y(n8886) );
	o22ai_1 U8960( .A1(n8764), .A2(n8973), .B1(n8927), .B2(n8964), .Y(n4365) );
	inv_1 U8961( .A(n7286), .Y(n8927) );
	o22ai_1 U8962( .A1(n8967), .A2(n8973), .B1(n8966), .B2(n5496), .Y(n4364) );
	o22ai_1 U8963( .A1(n8969), .A2(n8973), .B1(n8968), .B2(n5327), .Y(n4363) );
	inv_1 U8964( .A(n99), .Y(n8973) );
	nor2_1 U8965( .A(RST), .B(n7223), .Y(n99) );
	o22ai_1 U8966( .A1(n8764), .A2(n8974), .B1(n8926), .B2(n8964), .Y(n4362) );
	inv_1 U8967( .A(n7613), .Y(n8926) );
	o22ai_1 U8968( .A1(n8974), .A2(n8967), .B1(n8966), .B2(n5497), .Y(n4361) );
	o22ai_1 U8969( .A1(n8974), .A2(n8969), .B1(n8968), .B2(n5328), .Y(n4360) );
	inv_1 U8970( .A(n98), .Y(n8974) );
	nor2_1 U8971( .A(RST), .B(n7241), .Y(n98) );
	o22ai_1 U8972( .A1(n8764), .A2(n8975), .B1(n5376), .B2(n8964), .Y(n4359) );
	o22ai_1 U8973( .A1(n8967), .A2(n8975), .B1(n8966), .B2(n5498), .Y(n4358) );
	o22ai_1 U8974( .A1(n8969), .A2(n8975), .B1(n8968), .B2(n5329), .Y(n4357) );
	inv_1 U8975( .A(n97), .Y(n8975) );
	nor2_1 U8976( .A(RST), .B(n7269), .Y(n97) );
	o22ai_1 U8977( .A1(n8764), .A2(n8976), .B1(n8929), .B2(n8964), .Y(n4356) );
	inv_1 U8978( .A(n7325), .Y(n8929) );
	o22ai_1 U8979( .A1(n8967), .A2(n8976), .B1(n8966), .B2(n5661), .Y(n4355) );
	o22ai_1 U8980( .A1(n8969), .A2(n8976), .B1(n8968), .B2(n5641), .Y(n4354) );
	inv_1 U8981( .A(n96), .Y(n8976) );
	nor2_1 U8982( .A(RST), .B(n7244), .Y(n96) );
	o22ai_1 U8983( .A1(n8764), .A2(n8977), .B1(n8928), .B2(n8964), .Y(n4353) );
	inv_1 U8984( .A(n7616), .Y(n8928) );
	o22ai_1 U8985( .A1(n8967), .A2(n8977), .B1(n8966), .B2(n5499), .Y(n4352) );
	o22ai_1 U8986( .A1(n8969), .A2(n8977), .B1(n8968), .B2(n5330), .Y(n4351) );
	inv_1 U8987( .A(n95), .Y(n8977) );
	nor2_1 U8988( .A(RST), .B(n7282), .Y(n95) );
	o22ai_1 U8989( .A1(n8764), .A2(n8978), .B1(n5358), .B2(n8964), .Y(n4350) );
	o22ai_1 U8990( .A1(n8967), .A2(n8978), .B1(n8966), .B2(n5662), .Y(n4349) );
	o22ai_1 U8991( .A1(n8969), .A2(n8978), .B1(n8968), .B2(n5642), .Y(n4348) );
	inv_1 U8992( .A(n94), .Y(n8978) );
	nor2_1 U8993( .A(RST), .B(n7233), .Y(n94) );
	o22ai_1 U8994( .A1(n8964), .A2(n5436), .B1(n8764), .B2(n8959), .Y(n4347) );
	o22ai_1 U8995( .A1(n8966), .A2(n8896), .B1(n8959), .B2(n8967), .Y(n4346) );
	inv_1 U8996( .A(n7424), .Y(n8896) );
	o22ai_1 U8997( .A1(n8968), .A2(n8897), .B1(n8959), .B2(n8969), .Y(n4345) );
	inv_1 U8998( .A(n93), .Y(n8959) );
	nor2_1 U8999( .A(n7252), .B(RST), .Y(n93) );
	inv_1 U9000( .A(n7434), .Y(n8897) );
	o22ai_1 U9001( .A1(n8764), .A2(n8956), .B1(n8964), .B2(n5442), .Y(n4344) );
	nand2_1 U9002( .A(n5756), .B(n8764), .Y(n8964) );
	nand2_1 U9003( .A(n7719), .B(n7230), .Y(n8764) );
	o22ai_1 U9004( .A1(n8956), .A2(n8967), .B1(n8966), .B2(n8899), .Y(n4343) );
	inv_1 U9005( .A(n7435), .Y(n8899) );
	nand2_1 U9006( .A(n5756), .B(n8967), .Y(n8966) );
	nand2_1 U9007( .A(n7719), .B(g6313), .Y(n8967) );
	o22ai_1 U9008( .A1(n8956), .A2(n8969), .B1(n8968), .B2(n8900), .Y(n4342) );
	inv_1 U9009( .A(n7443), .Y(n8900) );
	nand2_1 U9010( .A(n5756), .B(n8969), .Y(n8968) );
	nand2_1 U9011( .A(n7719), .B(g6231), .Y(n8969) );
	inv_1 U9012( .A(n92), .Y(n8956) );
	nor2_1 U9013( .A(n7594), .B(RST), .Y(n92) );
	nor2_1 U9014( .A(RST), .B(g27380), .Y(n4341) );
	and2_0 U9015( .A(n5741), .B(g26135), .X(n4340) );
	and2_0 U9016( .A(n5761), .B(g26104), .X(n4339) );
	nor2_1 U9017( .A(RST), .B(n8979), .Y(n4338) );
	and2_0 U9018( .A(n5759), .B(g26149), .X(n4337) );
	and2_0 U9019( .A(n5764), .B(g25442), .X(n4336) );
	and2_0 U9020( .A(n5740), .B(g25435), .X(n4335) );
	and2_0 U9021( .A(n5765), .B(g25420), .X(n4334) );
	nor2_1 U9022( .A(RST), .B(g24734), .Y(n4333) );
	and2_0 U9023( .A(n5745), .B(g24734), .X(n4332) );
	o22ai_1 U9024( .A1(n8980), .A2(n5304), .B1(n5575), .B2(n8981), .Y(n4331) );
	o22ai_1 U9025( .A1(n8980), .A2(n8982), .B1(n5386), .B2(n8983), .Y(n4330) );
	o22ai_1 U9026( .A1(n8980), .A2(n8984), .B1(n5576), .B2(n8985), .Y(n4329) );
	o22ai_1 U9027( .A1(n5304), .A2(n8986), .B1(n5385), .B2(n8981), .Y(n4328) );
	o22ai_1 U9028( .A1(n8982), .A2(n8986), .B1(n5310), .B2(n8983), .Y(n4327) );
	o22ai_1 U9029( .A1(n8984), .A2(n8986), .B1(n5581), .B2(n8985), .Y(n4326) );
	o22ai_1 U9030( .A1(n5304), .A2(n8987), .B1(n5582), .B2(n8981), .Y(n4325) );
	o22ai_1 U9031( .A1(n8982), .A2(n8987), .B1(n5308), .B2(n8983), .Y(n4324) );
	o22ai_1 U9032( .A1(n8984), .A2(n8987), .B1(n5309), .B2(n8985), .Y(n4323) );
	o22ai_1 U9033( .A1(n5304), .A2(n8988), .B1(n5383), .B2(n8981), .Y(n4322) );
	o22ai_1 U9034( .A1(n8982), .A2(n8988), .B1(n5307), .B2(n8983), .Y(n4321) );
	o22ai_1 U9035( .A1(n8984), .A2(n8988), .B1(n5384), .B2(n8985), .Y(n4320) );
	o22ai_1 U9036( .A1(n5304), .A2(n8989), .B1(n5583), .B2(n8981), .Y(n4319) );
	inv_1 U9037( .A(n34), .Y(n8989) );
	o22ai_1 U9038( .A1(n8990), .A2(n8991), .B1(n5584), .B2(n8983), .Y(n4318) );
	o22ai_1 U9039( .A1(n8990), .A2(n8992), .B1(n5312), .B2(n8985), .Y(n4317) );
	o22ai_1 U9040( .A1(n5304), .A2(n6758), .B1(n5387), .B2(n8981), .Y(n4316) );
	o22ai_1 U9041( .A1(n8982), .A2(n6758), .B1(n5577), .B2(n8983), .Y(n4315) );
	o22ai_1 U9042( .A1(n8984), .A2(n6758), .B1(n5388), .B2(n8985), .Y(n4314) );
	nand2_1 U9043( .A(n8993), .B(n5744), .Y(n6758) );
	o22ai_1 U9044( .A1(n5304), .A2(n8994), .B1(n5578), .B2(n8981), .Y(n4313) );
	inv_1 U9045( .A(n31), .Y(n8994) );
	o22ai_1 U9046( .A1(n8991), .A2(n8995), .B1(n8996), .B2(n8983), .Y(n4312) );
	inv_1 U9047( .A(n7666), .Y(n8996) );
	o22ai_1 U9048( .A1(n8992), .A2(n8995), .B1(n5311), .B2(n8985), .Y(n4311) );
	o22ai_1 U9049( .A1(n5304), .A2(n8997), .B1(n5579), .B2(n8981), .Y(n4310) );
	o22ai_1 U9050( .A1(n8982), .A2(n8997), .B1(n5585), .B2(n8983), .Y(n4309) );
	o22ai_1 U9051( .A1(n8984), .A2(n8997), .B1(n5569), .B2(n8985), .Y(n4308) );
	inv_1 U9052( .A(n4487), .Y(n8997) );
	nor2_1 U9053( .A(n8998), .B(RST), .Y(n4487) );
	o22ai_1 U9054( .A1(n5737), .A2(n8981), .B1(n8999), .B2(n9000), .Y(n4307) );
	o22ai_1 U9055( .A1(n8991), .A2(n9000), .B1(n5586), .B2(n8983), .Y(n4306) );
	o22ai_1 U9056( .A1(n8992), .A2(n9000), .B1(n5314), .B2(n8985), .Y(n4305) );
	inv_1 U9057( .A(n7294), .Y(n9000) );
	o22ai_1 U9058( .A1(n5500), .A2(n8981), .B1(n8999), .B2(n9001), .Y(n4304) );
	o22ai_1 U9059( .A1(n8991), .A2(n9001), .B1(n5580), .B2(n8983), .Y(n4303) );
	o22ai_1 U9060( .A1(n8992), .A2(n9001), .B1(n5389), .B2(n8985), .Y(n4302) );
	inv_1 U9061( .A(n7289), .Y(n9001) );
	o22ai_1 U9062( .A1(n5717), .A2(n8981), .B1(n8999), .B2(n9002), .Y(n4301) );
	o22ai_1 U9063( .A1(n8991), .A2(n9002), .B1(n9003), .B2(n8983), .Y(n4300) );
	inv_1 U9064( .A(n7640), .Y(n9003) );
	nor2_1 U9065( .A(RST), .B(n7261), .Y(n43) );
	o22ai_1 U9066( .A1(n8992), .A2(n9002), .B1(n5313), .B2(n8985), .Y(n4299) );
	inv_1 U9067( .A(n7288), .Y(n9002) );
	o22ai_1 U9068( .A1(n5718), .A2(n8981), .B1(n8999), .B2(n9004), .Y(n4298) );
	nand2_1 U9069( .A(n10089), .B(n5744), .Y(n8999) );
	nand2_1 U9070( .A(n5304), .B(n5744), .Y(n8981) );
	o22ai_1 U9071( .A1(n8991), .A2(n9004), .B1(n5587), .B2(n8983), .Y(n4297) );
	nand2_1 U9072( .A(n8982), .B(n5744), .Y(n8983) );
	inv_1 U9073( .A(n4295), .Y(n8991) );
	o22ai_1 U9074( .A1(n8992), .A2(n9004), .B1(n5588), .B2(n8985), .Y(n4296) );
	nand2_1 U9075( .A(n8984), .B(n5744), .Y(n8985) );
	inv_1 U9076( .A(n7272), .Y(n9004) );
	inv_1 U9077( .A(n4209), .Y(n8992) );
	nor2_1 U9078( .A(n8982), .B(RST), .Y(n4295) );
	inv_1 U9079( .A(g8030), .Y(n8982) );
	and2_0 U9080( .A(g3213), .B(n5765), .X(n4294) );
	and2_0 U9081( .A(g3214), .B(n5764), .X(n4293) );
	and2_0 U9082( .A(g3215), .B(n5765), .X(n4292) );
	and2_0 U9083( .A(g3216), .B(n5764), .X(n4291) );
	and2_0 U9084( .A(g3217), .B(n5765), .X(n4290) );
	and2_0 U9085( .A(g3218), .B(n5764), .X(n4289) );
	and2_0 U9086( .A(g3219), .B(n5765), .X(n4288) );
	and2_0 U9087( .A(g3220), .B(n5764), .X(n4287) );
	and2_0 U9088( .A(g3221), .B(n5764), .X(n4286) );
	and2_0 U9089( .A(g3222), .B(n5764), .X(n4285) );
	and2_0 U9090( .A(g3223), .B(n5764), .X(n4284) );
	and2_0 U9091( .A(g3224), .B(n5763), .X(n4283) );
	and2_0 U9092( .A(g3225), .B(n5764), .X(n4282) );
	and2_0 U9093( .A(g3226), .B(n5764), .X(n4281) );
	and2_0 U9094( .A(g3227), .B(n5764), .X(n4280) );
	and2_0 U9095( .A(g3228), .B(n5764), .X(n4279) );
	inv_1 U9096( .A(n9005), .Y(n4278) );
	nor2_1 U9097( .A(RST), .B(n9006), .Y(n4277) );
	xnor2_1 U9098( .A(n9007), .B(g2962), .Y(n9006) );
	nor2_1 U9099( .A(RST), .B(n9008), .Y(n4276) );
	xnor2_1 U9100( .A(n9009), .B(g2934), .Y(n9008) );
	nor2_1 U9101( .A(n9010), .B(n9011), .Y(n4275) );
	xnor2_1 U9102( .A(n10066), .B(n9012), .Y(n9010) );
	nor3_1 U9103( .A(n9011), .B(n9012), .C(n9013), .Y(n4274) );
	a21oi_1 U9104( .A1(n10065), .A2(n9014), .B1(n7703), .Y(n9013) );
	and3_1 U9105( .A(n9014), .B(n7703), .C(n10065), .X(n9012) );
	nor2_1 U9106( .A(n9015), .B(n9011), .Y(n4273) );
	nand3_1 U9107( .A(n5751), .B(n5361), .C(n9016), .Y(n9011) );
	nand4_1 U9108( .A(n10066), .B(n9014), .C(n9017), .D(n5369), .Y(n9016) );
	xnor2_1 U9109( .A(n9014), .B(n10065), .Y(n9015) );
	nor2_1 U9110( .A(n9018), .B(n9019), .Y(n9014) );
	inv_1 U9111( .A(n7303), .Y(n9018) );
	a21oi_1 U9112( .A1(n9020), .A2(n5361), .B1(RST), .Y(n4272) );
	mux2i_1 U9113( .A0(n9021), .A1(n7303), .S(n9019), .Y(n9020) );
	nand2_1 U9114( .A(n7303), .B(n9022), .Y(n9021) );
	nand3_1 U9115( .A(n9017), .B(n5369), .C(n10066), .Y(n9022) );
	inv_1 U9116( .A(n7703), .Y(n9017) );
	nor2_1 U9117( .A(n9023), .B(n9024), .Y(n4271) );
	xnor2_1 U9118( .A(n7247), .B(n9025), .Y(n9023) );
	and2_0 U9119( .A(n9026), .B(n7320), .X(n9025) );
	nor2_1 U9120( .A(n9027), .B(n9024), .Y(n4270) );
	xnor2_1 U9121( .A(n9026), .B(n7320), .Y(n9027) );
	nor3_1 U9122( .A(n9024), .B(n9026), .C(n9028), .Y(n4269) );
	a21oi_1 U9123( .A1(n9029), .A2(n7279), .B1(n7321), .Y(n9028) );
	and3_1 U9124( .A(n7321), .B(n7279), .C(n9029), .X(n9026) );
	nor2_1 U9125( .A(n9030), .B(n9024), .Y(n4268) );
	xnor2_1 U9126( .A(n7279), .B(n9029), .Y(n9030) );
	nor3_1 U9127( .A(n9024), .B(n9029), .C(n9031), .Y(n4267) );
	a21oi_1 U9128( .A1(n9032), .A2(n7721), .B1(n10084), .Y(n9031) );
	and3_1 U9129( .A(n9032), .B(n7721), .C(n10084), .X(n9029) );
	nor2_1 U9130( .A(n9033), .B(n9024), .Y(n4266) );
	or2_0 U9131( .A(n9034), .B(RST), .X(n9024) );
	xnor2_1 U9132( .A(n9032), .B(n7721), .Y(n9033) );
	nor3_1 U9133( .A(n14868), .B(g51), .C(RST), .Y(n4265) );
	nor2_1 U9134( .A(g51), .B(n9035), .Y(n4264) );
	mux2i_1 U9135( .A0(n5796), .A1(n9036), .S(n9037), .Y(n4263) );
	nand2_1 U9136( .A(g2466), .B(n5742), .Y(n5796) );
	mux2i_1 U9137( .A0(n5797), .A1(n9036), .S(n9038), .Y(n4262) );
	nand2_1 U9138( .A(g2463), .B(n5742), .Y(n5797) );
	mux2i_1 U9139( .A0(n5798), .A1(n9039), .S(n9037), .Y(n4261) );
	nand2_1 U9140( .A(g2451), .B(n5742), .Y(n5798) );
	mux2i_1 U9141( .A0(n5804), .A1(n9039), .S(n9038), .Y(n4260) );
	nand2_1 U9142( .A(g2448), .B(n5742), .Y(n5804) );
	mux2i_1 U9143( .A0(n5996), .A1(n9040), .S(n9037), .Y(n4259) );
	nand2_1 U9144( .A(g2436), .B(n5742), .Y(n5996) );
	mux2i_1 U9145( .A0(n6355), .A1(n9040), .S(n9038), .Y(n4258) );
	nand2_1 U9146( .A(g2433), .B(n5742), .Y(n6355) );
	mux2i_1 U9147( .A0(n6614), .A1(n9041), .S(n9037), .Y(n4257) );
	nor2_1 U9148( .A(n9042), .B(n6265), .Y(n9037) );
	nand2_1 U9149( .A(g2421), .B(n5742), .Y(n6614) );
	mux2i_1 U9150( .A0(n6876), .A1(n9041), .S(n9038), .Y(n4256) );
	nor2_1 U9151( .A(n9042), .B(n6264), .Y(n9038) );
	nand2_1 U9152( .A(g2418), .B(n5742), .Y(n6876) );
	mux2i_1 U9153( .A0(n9043), .A1(n9044), .S(n9045), .Y(n4255) );
	mux2i_1 U9154( .A0(n9046), .A1(n9044), .S(n9047), .Y(n4254) );
	mux2i_1 U9155( .A0(n9048), .A1(n9049), .S(n9045), .Y(n4253) );
	mux2i_1 U9156( .A0(n9050), .A1(n9049), .S(n9047), .Y(n4252) );
	mux2i_1 U9157( .A0(n9051), .A1(n9052), .S(n9045), .Y(n4251) );
	mux2i_1 U9158( .A0(n9053), .A1(n9052), .S(n9047), .Y(n4250) );
	mux2i_1 U9159( .A0(n9054), .A1(n9055), .S(n9045), .Y(n4249) );
	and2_0 U9160( .A(n9056), .B(n7782), .X(n9045) );
	mux2i_1 U9161( .A0(n9057), .A1(n9055), .S(n9047), .Y(n4248) );
	and2_0 U9162( .A(n9056), .B(g7014), .X(n9047) );
	mux2i_1 U9163( .A0(n9058), .A1(n9059), .S(n9060), .Y(n4247) );
	mux2i_1 U9164( .A0(n9061), .A1(n9059), .S(n9062), .Y(n4246) );
	mux2i_1 U9165( .A0(n9063), .A1(n9064), .S(n9060), .Y(n4245) );
	mux2i_1 U9166( .A0(n9065), .A1(n9064), .S(n9062), .Y(n4244) );
	inv_1 U9167( .A(n143), .Y(n9065) );
	mux2i_1 U9168( .A0(n9066), .A1(n9067), .S(n9060), .Y(n4243) );
	mux2i_1 U9169( .A0(n9068), .A1(n9067), .S(n9062), .Y(n4242) );
	inv_1 U9170( .A(n141), .Y(n9068) );
	mux2i_1 U9171( .A0(n9069), .A1(n9070), .S(n9060), .Y(n4241) );
	nor2_1 U9172( .A(n9071), .B(n7927), .Y(n9060) );
	mux2i_1 U9173( .A0(n9072), .A1(n9070), .S(n9062), .Y(n4240) );
	nor2_1 U9174( .A(n9071), .B(n8032), .Y(n9062) );
	inv_1 U9175( .A(n139), .Y(n9072) );
	mux2i_1 U9176( .A0(n9073), .A1(n9074), .S(n9075), .Y(n4239) );
	mux2i_1 U9177( .A0(n9076), .A1(n9074), .S(n9077), .Y(n4238) );
	mux2i_1 U9178( .A0(n9078), .A1(n9079), .S(n9075), .Y(n4237) );
	mux2i_1 U9179( .A0(n9080), .A1(n9079), .S(n9077), .Y(n4236) );
	mux2i_1 U9180( .A0(n9081), .A1(n9082), .S(n9075), .Y(n4235) );
	mux2i_1 U9181( .A0(n9083), .A1(n9082), .S(n9077), .Y(n4234) );
	mux2i_1 U9182( .A0(n9084), .A1(n9085), .S(n9075), .Y(n4233) );
	nor2_1 U9183( .A(n9086), .B(n8693), .Y(n9075) );
	mux2i_1 U9184( .A0(n9087), .A1(n9085), .S(n9077), .Y(n4232) );
	nor2_1 U9185( .A(n9086), .B(n8692), .Y(n9077) );
	nor2_1 U9186( .A(n5888), .B(RST), .Y(n4231) );
	inv_1 U9187( .A(g3080), .Y(n5888) );
	and2_0 U9188( .A(n5752), .B(n9088), .X(n4230) );
	and2_0 U9189( .A(n5756), .B(n9089), .X(n4229) );
	mux2i_1 U9190( .A0(n9090), .A1(n9036), .S(n9091), .Y(n4228) );
	nand2_1 U9191( .A(n5757), .B(n9092), .Y(n9036) );
	nand3_1 U9192( .A(n9093), .B(n9094), .C(n9095), .Y(n9092) );
	inv_1 U9193( .A(n9096), .Y(n9094) );
	mux2i_1 U9194( .A0(n9097), .A1(n9039), .S(n9091), .Y(n4227) );
	nand2_1 U9195( .A(n9098), .B(n5741), .Y(n9039) );
	mux2i_1 U9196( .A0(n9099), .A1(n9100), .S(n9096), .Y(n9098) );
	mux2i_1 U9197( .A0(n6098), .A1(g3229), .S(n9101), .Y(n9100) );
	nor2_1 U9198( .A(n9093), .B(n9102), .Y(n9099) );
	mux2i_1 U9199( .A0(n9103), .A1(n9040), .S(n9091), .Y(n4226) );
	o211ai_1 U9200( .A1(n9095), .A2(n9093), .B1(n9104), .C1(n5740), .Y(n9040) );
	xnor2_1 U9201( .A(n9105), .B(g3229), .Y(n9093) );
	mux2i_1 U9202( .A0(n9106), .A1(n9041), .S(n9091), .Y(n4225) );
	nor2_1 U9203( .A(n9042), .B(n6281), .Y(n9091) );
	o21ai_0 U9204( .A1(n6121), .A2(n6131), .B1(n6130), .Y(n9042) );
	o211ai_1 U9205( .A1(n6098), .A2(n9107), .B1(n5740), .C1(n9108), .Y(n9041) );
	mux2i_1 U9206( .A0(n5983), .A1(n9109), .S(n9104), .Y(n9108) );
	nand2_1 U9207( .A(n9095), .B(n9096), .Y(n9104) );
	o221ai_1 U9208( .A1(g2436), .A2(n6265), .B1(g2444), .B2(n6281), .C1(n9110), .Y(n9096) );
	or2_0 U9209( .A(n6264), .B(g2433), .X(n9110) );
	inv_1 U9210( .A(n9111), .Y(n9095) );
	o221ai_1 U9211( .A1(g2451), .A2(n6265), .B1(g2459), .B2(n6281), .C1(n9112), .Y(n9111) );
	or2_0 U9212( .A(n6264), .B(g2448), .X(n9112) );
	nor2_1 U9213( .A(n9105), .B(n9102), .Y(n9109) );
	inv_1 U9214( .A(n9101), .Y(n9105) );
	o221ai_1 U9215( .A1(g2421), .A2(n6265), .B1(g2429), .B2(n6281), .C1(n9113), .Y(n9101) );
	or2_0 U9216( .A(n6264), .B(g2418), .X(n9113) );
	inv_1 U9217( .A(n9102), .Y(n9107) );
	o221ai_1 U9218( .A1(g2466), .A2(n6265), .B1(g2473), .B2(n6281), .C1(n9114), .Y(n9102) );
	or2_0 U9219( .A(n6264), .B(g2463), .X(n9114) );
	inv_1 U9220( .A(n7780), .Y(n6265) );
	mux2i_1 U9221( .A0(n9115), .A1(n9044), .S(n9116), .Y(n4224) );
	nand2_1 U9222( .A(n5755), .B(n9117), .Y(n9044) );
	nand3_1 U9223( .A(n9118), .B(n9119), .C(n9120), .Y(n9117) );
	inv_1 U9224( .A(n9121), .Y(n9119) );
	mux2i_1 U9225( .A0(n9122), .A1(n9049), .S(n9116), .Y(n4223) );
	nand2_1 U9226( .A(n9123), .B(n5747), .Y(n9049) );
	mux2i_1 U9227( .A0(n9124), .A1(n9125), .S(n9121), .Y(n9123) );
	mux2i_1 U9228( .A0(n6098), .A1(g3229), .S(n9126), .Y(n9125) );
	nor2_1 U9229( .A(n9118), .B(n9127), .Y(n9124) );
	mux2i_1 U9230( .A0(n9128), .A1(n9052), .S(n9116), .Y(n4222) );
	o211ai_1 U9231( .A1(n9120), .A2(n9118), .B1(n9129), .C1(n5740), .Y(n9052) );
	xnor2_1 U9232( .A(n9130), .B(g3229), .Y(n9118) );
	mux2i_1 U9233( .A0(n9131), .A1(n9055), .S(n9116), .Y(n4221) );
	and2_0 U9234( .A(n9056), .B(g5511), .X(n9116) );
	a21oi_1 U9235( .A1(n9132), .A2(n6337), .B1(n9133), .Y(n9056) );
	o211ai_1 U9236( .A1(n6098), .A2(n9134), .B1(n5740), .C1(n9135), .Y(n9055) );
	mux2i_1 U9237( .A0(n5983), .A1(n9136), .S(n9129), .Y(n9135) );
	nand2_1 U9238( .A(n9120), .B(n9121), .Y(n9129) );
	o221ai_1 U9239( .A1(g1742), .A2(n6888), .B1(g1750), .B2(n6939), .C1(n9137), .Y(n9121) );
	or2_0 U9240( .A(n6774), .B(g1739), .X(n9137) );
	inv_1 U9241( .A(n9138), .Y(n9120) );
	o221ai_1 U9242( .A1(g1757), .A2(n6888), .B1(g1765), .B2(n6939), .C1(n9139), .Y(n9138) );
	or2_0 U9243( .A(n6774), .B(g1754), .X(n9139) );
	nor2_1 U9244( .A(n9130), .B(n9127), .Y(n9136) );
	inv_1 U9245( .A(n9126), .Y(n9130) );
	o221ai_1 U9246( .A1(g1727), .A2(n6888), .B1(g1735), .B2(n6939), .C1(n9140), .Y(n9126) );
	or2_0 U9247( .A(n6774), .B(g1724), .X(n9140) );
	inv_1 U9248( .A(n9127), .Y(n9134) );
	o221ai_1 U9249( .A1(g1772), .A2(n6888), .B1(g1779), .B2(n6939), .C1(n9141), .Y(n9127) );
	or2_0 U9250( .A(n6774), .B(g1769), .X(n9141) );
	inv_1 U9251( .A(n7782), .Y(n6888) );
	mux2i_1 U9252( .A0(n9142), .A1(n9059), .S(n9143), .Y(n4220) );
	nand2_1 U9253( .A(n5757), .B(n9144), .Y(n9059) );
	nand3_1 U9254( .A(n9145), .B(n9146), .C(n9147), .Y(n9144) );
	mux2i_1 U9255( .A0(n9148), .A1(n9064), .S(n9143), .Y(n4219) );
	nand2_1 U9256( .A(n9149), .B(n5741), .Y(n9064) );
	mux2i_1 U9257( .A0(n9150), .A1(n9151), .S(n9152), .Y(n9149) );
	mux2i_1 U9258( .A0(g3229), .A1(n6098), .S(n9153), .Y(n9151) );
	nor2_1 U9259( .A(n9145), .B(n9154), .Y(n9150) );
	mux2i_1 U9260( .A0(n9155), .A1(n9067), .S(n9143), .Y(n4218) );
	o211ai_1 U9261( .A1(n9147), .A2(n9145), .B1(n9156), .C1(n5740), .Y(n9067) );
	xnor2_1 U9262( .A(n9153), .B(g3229), .Y(n9145) );
	mux2i_1 U9263( .A0(n9157), .A1(n9070), .S(n9143), .Y(n4217) );
	nor2_1 U9264( .A(n9071), .B(n7932), .Y(n9143) );
	o21ai_0 U9265( .A1(n7986), .A2(n6131), .B1(n9158), .Y(n9071) );
	o211ai_1 U9266( .A1(n6098), .A2(n9159), .B1(n5741), .C1(n9160), .Y(n9070) );
	mux2i_1 U9267( .A0(n5983), .A1(n9161), .S(n9156), .Y(n9160) );
	nand2_1 U9268( .A(n9147), .B(n9152), .Y(n9156) );
	inv_1 U9269( .A(n9146), .Y(n9152) );
	a21oi_1 U9270( .A1(n9162), .A2(g5472), .B1(n9163), .Y(n9146) );
	o22ai_1 U9271( .A1(n7932), .A2(g1045), .B1(n7927), .B2(g1048), .Y(n9163) );
	a21oi_1 U9272( .A1(n9164), .A2(g5472), .B1(n9165), .Y(n9147) );
	o22ai_1 U9273( .A1(n7932), .A2(g1060), .B1(n7927), .B2(g1063), .Y(n9165) );
	nor2_1 U9274( .A(n9153), .B(n9154), .Y(n9161) );
	inv_1 U9275( .A(n9159), .Y(n9154) );
	a21oi_1 U9276( .A1(n9166), .A2(g5472), .B1(n9167), .Y(n9153) );
	o22ai_1 U9277( .A1(n7932), .A2(g1030), .B1(n7927), .B2(g1033), .Y(n9167) );
	a21oi_1 U9278( .A1(n9168), .A2(g5472), .B1(n9169), .Y(n9159) );
	o22ai_1 U9279( .A1(n7932), .A2(g1075), .B1(n7927), .B2(g1078), .Y(n9169) );
	inv_1 U9280( .A(n7775), .Y(n7927) );
	inv_1 U9281( .A(g1085), .Y(n9168) );
	mux2i_1 U9282( .A0(n9170), .A1(n9074), .S(n9171), .Y(n4216) );
	nand2_1 U9283( .A(n5757), .B(n9172), .Y(n9074) );
	nand3_1 U9284( .A(n9173), .B(n9174), .C(n9175), .Y(n9172) );
	inv_1 U9285( .A(n9176), .Y(n9174) );
	mux2i_1 U9286( .A0(n9177), .A1(n9079), .S(n9171), .Y(n4215) );
	nand2_1 U9287( .A(n9178), .B(n5741), .Y(n9079) );
	mux2i_1 U9288( .A0(n9179), .A1(n9180), .S(n9176), .Y(n9178) );
	mux2i_1 U9289( .A0(n6098), .A1(g3229), .S(n9181), .Y(n9180) );
	nor2_1 U9290( .A(n9173), .B(n9182), .Y(n9179) );
	mux2i_1 U9291( .A0(n9183), .A1(n9082), .S(n9171), .Y(n4214) );
	o211ai_1 U9292( .A1(n9175), .A2(n9173), .B1(n9184), .C1(n5740), .Y(n9082) );
	xnor2_1 U9293( .A(n9185), .B(g3229), .Y(n9173) );
	mux2i_1 U9294( .A0(n9186), .A1(n9085), .S(n9171), .Y(n4213) );
	nor2_1 U9295( .A(n9086), .B(n8709), .Y(n9171) );
	o21ai_0 U9296( .A1(n8554), .A2(n6131), .B1(n8563), .Y(n9086) );
	o211ai_1 U9297( .A1(n6098), .A2(n9187), .B1(n5741), .C1(n9188), .Y(n9085) );
	mux2i_1 U9298( .A0(n5983), .A1(n9189), .S(n9184), .Y(n9188) );
	nand2_1 U9299( .A(n9175), .B(n9176), .Y(n9184) );
	o221ai_1 U9300( .A1(g361), .A2(n8693), .B1(g369), .B2(n8709), .C1(n9190), .Y(n9176) );
	or2_0 U9301( .A(n8692), .B(g358), .X(n9190) );
	inv_1 U9302( .A(n9191), .Y(n9175) );
	o221ai_1 U9303( .A1(g376), .A2(n8693), .B1(g384), .B2(n8709), .C1(n9192), .Y(n9191) );
	or2_0 U9304( .A(n8692), .B(g373), .X(n9192) );
	nor2_1 U9305( .A(n9185), .B(n9182), .Y(n9189) );
	inv_1 U9306( .A(n9181), .Y(n9185) );
	o221ai_1 U9307( .A1(g346), .A2(n8693), .B1(g354), .B2(n8709), .C1(n9193), .Y(n9181) );
	or2_0 U9308( .A(n8692), .B(g343), .X(n9193) );
	inv_1 U9309( .A(g3229), .Y(n5983) );
	inv_1 U9310( .A(n9182), .Y(n9187) );
	o221ai_1 U9311( .A1(g391), .A2(n8693), .B1(g398), .B2(n8709), .C1(n9194), .Y(n9182) );
	or2_0 U9312( .A(n8692), .B(g388), .X(n9194) );
	inv_1 U9313( .A(n7784), .Y(n8693) );
	and2_0 U9314( .A(g2623), .B(n5764), .X(n4212) );
	and2_0 U9315( .A(g1235), .B(n5764), .X(n4211) );
	and2_0 U9316( .A(g549), .B(n5763), .X(n4210) );
	nor2_1 U9317( .A(n8984), .B(RST), .Y(n4209) );
	inv_1 U9318( .A(g8106), .Y(n8984) );
	and2_0 U9319( .A(g1929), .B(n5764), .X(n4208) );
	and2_0 U9320( .A(n5751), .B(g5747), .X(n4207) );
	and2_0 U9321( .A(n5755), .B(g5695), .X(n4206) );
	and2_0 U9322( .A(n5745), .B(g5657), .X(n4205) );
	and2_0 U9323( .A(n5759), .B(g5629), .X(n4204) );
	o21ai_0 U9324( .A1(RST), .A2(n9195), .B1(n9196), .Y(n4203) );
	nand4_1 U9325( .A(n9863), .B(n9197), .C(n9198), .D(n6098), .Y(n9196) );
	a221oi_1 U9326( .A1(n7588), .A2(n9199), .B1(n7290), .B2(n9200), .C1(n9201), .Y(n9195) );
	and4_1 U9327( .A(n9872), .B(g3229), .C(n9198), .D(n9197), .X(n9201) );
	inv_1 U9328( .A(n9202), .Y(n9198) );
	xor2_1 U9329( .A(n9203), .B(n9204), .X(n9200) );
	xor2_1 U9330( .A(n9205), .B(n9206), .X(n9199) );
	xor2_1 U9331( .A(n9207), .B(n9208), .X(n9206) );
	xor2_1 U9332( .A(n9209), .B(n9210), .X(n9208) );
	xor2_1 U9333( .A(n9211), .B(n9212), .X(n9207) );
	xor2_1 U9334( .A(n9213), .B(n9214), .X(n9205) );
	xor2_1 U9335( .A(n9215), .B(n9216), .X(n9214) );
	xor2_1 U9336( .A(n9217), .B(n9218), .X(n9213) );
	a21oi_1 U9337( .A1(n9219), .A2(n9220), .B1(RST), .Y(n4202) );
	nand2_1 U9338( .A(n9221), .B(n9204), .Y(n9220) );
	nand2_1 U9339( .A(n9222), .B(n9223), .Y(n9204) );
	mux2i_1 U9340( .A0(n5944), .A1(n9224), .S(n5926), .Y(n9222) );
	o221ai_1 U9341( .A1(n9225), .A2(n9210), .B1(g2611), .B2(n9202), .C1(n9197), .Y(n9219) );
	mux2i_1 U9342( .A0(n9226), .A1(n9227), .S(n5930), .Y(n9210) );
	a21oi_1 U9343( .A1(n9228), .A2(n9229), .B1(RST), .Y(n4201) );
	nand2_1 U9344( .A(n9221), .B(n9203), .Y(n9229) );
	nand2_1 U9345( .A(n9230), .B(n9231), .Y(n9203) );
	mux2i_1 U9346( .A0(n5940), .A1(n9232), .S(n5925), .Y(n9230) );
	o221ai_1 U9347( .A1(n9225), .A2(n9211), .B1(g2610), .B2(n9202), .C1(n9197), .Y(n9228) );
	nand2_1 U9348( .A(n9233), .B(n9231), .Y(n9211) );
	mux2i_1 U9349( .A0(n5940), .A1(n9232), .S(n5920), .Y(n9233) );
	o21ai_0 U9350( .A1(n9234), .A2(n9235), .B1(n9236), .Y(n4200) );
	o22ai_1 U9351( .A1(n9225), .A2(n9216), .B1(g2608), .B2(n9202), .Y(n9235) );
	nand2_1 U9352( .A(n9237), .B(n9223), .Y(n9216) );
	a21oi_1 U9353( .A1(n5944), .A2(n9238), .B1(n9239), .Y(n9223) );
	mux2i_1 U9354( .A0(n9224), .A1(n5944), .S(n5924), .Y(n9237) );
	nor2_1 U9355( .A(RST), .B(n7273), .Y(n42) );
	o21ai_0 U9356( .A1(n9234), .A2(n9240), .B1(n9236), .Y(n4199) );
	o22ai_1 U9357( .A1(n9225), .A2(n9215), .B1(g2607), .B2(n9202), .Y(n9240) );
	nand2_1 U9358( .A(n9241), .B(n9231), .Y(n9215) );
	a21oi_1 U9359( .A1(n5940), .A2(n9238), .B1(n9239), .Y(n9231) );
	mux2i_1 U9360( .A0(n5940), .A1(n9232), .S(n5932), .Y(n9241) );
	a21oi_1 U9361( .A1(n9242), .A2(n9243), .B1(RST), .Y(n4198) );
	o221ai_1 U9362( .A1(n9225), .A2(n9209), .B1(g2606), .B2(n9202), .C1(n9197), .Y(n9243) );
	mux2i_1 U9363( .A0(n9226), .A1(n9227), .S(n5919), .Y(n9209) );
	o21ai_0 U9364( .A1(n9234), .A2(n9244), .B1(n9245), .Y(n4197) );
	o22ai_1 U9365( .A1(n9225), .A2(n9218), .B1(g2605), .B2(n9202), .Y(n9244) );
	nand2_1 U9366( .A(n9246), .B(n9247), .Y(n9218) );
	mux2i_1 U9367( .A0(n5940), .A1(n9232), .S(n5931), .Y(n9246) );
	o21ai_0 U9368( .A1(n9234), .A2(n9248), .B1(n9245), .Y(n4196) );
	and2_0 U9369( .A(n9236), .B(n9249), .X(n9245) );
	nand3_1 U9370( .A(n47), .B(n9250), .C(n9221), .Y(n9249) );
	inv_1 U9371( .A(n8980), .Y(n47) );
	nand2_1 U9372( .A(g2574), .B(n5741), .Y(n8980) );
	nand2_1 U9373( .A(n9251), .B(n5742), .Y(n9236) );
	o22ai_1 U9374( .A1(n9225), .A2(n9212), .B1(g2604), .B2(n9202), .Y(n9248) );
	mux2i_1 U9375( .A0(n9226), .A1(n9227), .S(n5934), .Y(n9212) );
	nor2_1 U9376( .A(n9239), .B(n9224), .Y(n9227) );
	nor2_1 U9377( .A(n5944), .B(n9238), .Y(n9224) );
	nor2_1 U9378( .A(n9239), .B(n5944), .Y(n9226) );
	nand2_1 U9379( .A(n9197), .B(n5742), .Y(n9234) );
	a21oi_1 U9380( .A1(n9242), .A2(n9252), .B1(RST), .Y(n4195) );
	o221ai_1 U9381( .A1(n9225), .A2(n9217), .B1(g2603), .B2(n9202), .C1(n9197), .Y(n9252) );
	nand2_1 U9382( .A(n9225), .B(n9253), .Y(n9202) );
	nand2_1 U9383( .A(n9254), .B(n9247), .Y(n9217) );
	inv_1 U9384( .A(n9239), .Y(n9247) );
	nand2_1 U9385( .A(n9253), .B(g2574), .Y(n9239) );
	mux2i_1 U9386( .A0(n5940), .A1(n9232), .S(n5935), .Y(n9254) );
	nor2_1 U9387( .A(n5940), .B(n9238), .Y(n9232) );
	inv_1 U9388( .A(n9255), .Y(n9225) );
	nor2_1 U9389( .A(n9256), .B(n9251), .Y(n9242) );
	nor2_1 U9390( .A(n9257), .B(n9253), .Y(n9251) );
	nor3_1 U9391( .A(n7294), .B(g2637), .C(n9258), .Y(n9253) );
	a21oi_1 U9392( .A1(n9250), .A2(g2574), .B1(n9257), .Y(n9256) );
	inv_1 U9393( .A(n9221), .Y(n9257) );
	nor2_1 U9394( .A(n9255), .B(n9197), .Y(n9221) );
	a21oi_1 U9395( .A1(n5574), .A2(n5982), .B1(n7290), .Y(n9197) );
	o21ai_0 U9396( .A1(n7290), .A2(n9959), .B1(n5982), .Y(n9255) );
	inv_1 U9397( .A(n7588), .Y(n5982) );
	o221ai_1 U9398( .A1(n7498), .A2(n5943), .B1(n7475), .B2(n5942), .C1(n9259), .Y(n9250) );
	a21oi_1 U9399( .A1(g7425), .A2(n5904), .B1(n9238), .Y(n9259) );
	and4_1 U9400( .A(n9260), .B(n9261), .C(n9262), .D(n9263), .X(n9238) );
	and3_1 U9401( .A(n5932), .B(n5920), .C(n5925), .X(n9263) );
	o221ai_1 U9402( .A1(n7476), .A2(n5943), .B1(n7477), .B2(n5942), .C1(n9264), .Y(n5925) );
	nand2_1 U9403( .A(g7425), .B(n5443), .Y(n9264) );
	o221ai_1 U9404( .A1(n7482), .A2(n5943), .B1(n7483), .B2(n5942), .C1(n9265), .Y(n5920) );
	nand2_1 U9405( .A(g7425), .B(n5444), .Y(n9265) );
	o221ai_1 U9406( .A1(n7484), .A2(n5943), .B1(n7485), .B2(n5942), .C1(n9266), .Y(n5932) );
	nand2_1 U9407( .A(g7425), .B(n5445), .Y(n9266) );
	nor3_1 U9408( .A(n9267), .B(n9268), .C(n5924), .Y(n9262) );
	a221oi_1 U9409( .A1(n5961), .A2(g7487), .B1(n5960), .B2(n7236), .C1(n9269), .Y(n5924) );
	nor2_1 U9410( .A(n5945), .B(n10039), .Y(n9269) );
	inv_1 U9411( .A(g7425), .Y(n5945) );
	inv_1 U9412( .A(n7481), .Y(n5960) );
	inv_1 U9413( .A(n7480), .Y(n5961) );
	inv_1 U9414( .A(n5926), .Y(n9268) );
	o221ai_1 U9415( .A1(n7478), .A2(n5943), .B1(n7479), .B2(n5942), .C1(n9270), .Y(n5926) );
	nand2_1 U9416( .A(g7425), .B(n5446), .Y(n9270) );
	a222oi_1 U9417( .A1(n7236), .A2(n5889), .B1(g7425), .B2(n5543), .C1(g7487), .C2(n5334), .Y(n9267) );
	inv_1 U9418( .A(n7315), .Y(n5889) );
	nor3_1 U9419( .A(n5931), .B(n9271), .C(n5919), .Y(n9261) );
	o221ai_1 U9420( .A1(n7493), .A2(n5943), .B1(n7494), .B2(n5942), .C1(n9272), .Y(n5919) );
	nand2_1 U9421( .A(g7425), .B(n5447), .Y(n9272) );
	inv_1 U9422( .A(n9273), .Y(n9271) );
	o211ai_1 U9423( .A1(n5942), .A2(n9871), .B1(n5907), .C1(n5906), .Y(n9273) );
	nand2_1 U9424( .A(g7487), .B(n5938), .Y(n5906) );
	inv_1 U9425( .A(n7486), .Y(n5938) );
	nand2_1 U9426( .A(g7425), .B(n5448), .Y(n5907) );
	o221ai_1 U9427( .A1(n7491), .A2(n5943), .B1(n7492), .B2(n5942), .C1(n9274), .Y(n5931) );
	nand2_1 U9428( .A(g7425), .B(n5449), .Y(n9274) );
	nor3_1 U9429( .A(n5935), .B(n5930), .C(n5934), .Y(n9260) );
	o221ai_1 U9430( .A1(n7489), .A2(n5943), .B1(n7490), .B2(n5942), .C1(n9275), .Y(n5934) );
	nand2_1 U9431( .A(g7425), .B(n5450), .Y(n9275) );
	o221ai_1 U9432( .A1(n7495), .A2(n5943), .B1(n7496), .B2(n5942), .C1(n9276), .Y(n5930) );
	nand2_1 U9433( .A(g7425), .B(n5451), .Y(n9276) );
	o221ai_1 U9434( .A1(n7487), .A2(n5943), .B1(n7488), .B2(n5942), .C1(n9277), .Y(n5935) );
	nand2_1 U9435( .A(g7425), .B(n5452), .Y(n9277) );
	inv_1 U9436( .A(n7497), .Y(n5904) );
	inv_1 U9437( .A(n7236), .Y(n5942) );
	inv_1 U9438( .A(g7487), .Y(n5943) );
	o21ai_0 U9439( .A1(RST), .A2(n9278), .B1(n9279), .Y(n4194) );
	nand4_1 U9440( .A(n9864), .B(n9280), .C(n9281), .D(n6098), .Y(n9279) );
	a221oi_1 U9441( .A1(n7589), .A2(n9282), .B1(n7291), .B2(n9283), .C1(n9284), .Y(n9278) );
	and4_1 U9442( .A(g3229), .B(n9914), .C(n9281), .D(n9280), .X(n9284) );
	xor2_1 U9443( .A(n9285), .B(n9286), .X(n9283) );
	xor2_1 U9444( .A(n9287), .B(n9288), .X(n9282) );
	xor2_1 U9445( .A(n9289), .B(n9290), .X(n9288) );
	xor2_1 U9446( .A(n9291), .B(n9292), .X(n9290) );
	xor2_1 U9447( .A(n9293), .B(n9294), .X(n9289) );
	xor2_1 U9448( .A(n9295), .B(n9296), .X(n9287) );
	xor2_1 U9449( .A(n9297), .B(n9298), .X(n9296) );
	xor2_1 U9450( .A(n9299), .B(n9300), .X(n9295) );
	a21oi_1 U9451( .A1(n9301), .A2(n9302), .B1(RST), .Y(n4193) );
	nand2_1 U9452( .A(n9303), .B(n9286), .Y(n9302) );
	nand2_1 U9453( .A(n9304), .B(n9305), .Y(n9286) );
	mux2i_1 U9454( .A0(n6662), .A1(n9306), .S(n6582), .Y(n9304) );
	o221ai_1 U9455( .A1(n9307), .A2(n9291), .B1(g1917), .B2(n9308), .C1(n9281), .Y(n9301) );
	mux2i_1 U9456( .A0(n9309), .A1(n9310), .S(n6586), .Y(n9291) );
	a21oi_1 U9457( .A1(n9311), .A2(n9312), .B1(RST), .Y(n4192) );
	nand2_1 U9458( .A(n9303), .B(n9285), .Y(n9312) );
	nand2_1 U9459( .A(n9313), .B(n9314), .Y(n9285) );
	mux2i_1 U9460( .A0(n6653), .A1(n9315), .S(n6581), .Y(n9313) );
	o221ai_1 U9461( .A1(n9307), .A2(n9298), .B1(g1916), .B2(n9308), .C1(n9281), .Y(n9311) );
	nand2_1 U9462( .A(n9316), .B(n9314), .Y(n9298) );
	mux2i_1 U9463( .A0(n6653), .A1(n9315), .S(n6576), .Y(n9316) );
	o21ai_0 U9464( .A1(n9317), .A2(n9318), .B1(n9319), .Y(n4191) );
	o22ai_1 U9465( .A1(n9307), .A2(n9300), .B1(g1914), .B2(n9308), .Y(n9318) );
	nand2_1 U9466( .A(n9320), .B(n9305), .Y(n9300) );
	a21oi_1 U9467( .A1(n6662), .A2(n9321), .B1(n9322), .Y(n9305) );
	mux2i_1 U9468( .A0(n9306), .A1(n6662), .S(n6580), .Y(n9320) );
	a21oi_1 U9469( .A1(n9323), .A2(n9324), .B1(RST), .Y(n4190) );
	o221ai_1 U9470( .A1(n9307), .A2(n9294), .B1(g1912), .B2(n9308), .C1(n9281), .Y(n9324) );
	mux2i_1 U9471( .A0(n9309), .A1(n9310), .S(n6575), .Y(n9294) );
	o21ai_0 U9472( .A1(n9317), .A2(n9325), .B1(n9326), .Y(n4189) );
	o22ai_1 U9473( .A1(n9307), .A2(n9299), .B1(g1911), .B2(n9308), .Y(n9325) );
	nand2_1 U9474( .A(n9327), .B(n9328), .Y(n9299) );
	mux2i_1 U9475( .A0(n6653), .A1(n9315), .S(n6588), .Y(n9327) );
	o21ai_0 U9476( .A1(n9317), .A2(n9329), .B1(n9326), .Y(n4188) );
	and2_0 U9477( .A(n9319), .B(n9330), .X(n9326) );
	nand3_1 U9478( .A(n32), .B(n9331), .C(n9303), .Y(n9330) );
	o22ai_1 U9479( .A1(n9307), .A2(n9292), .B1(g1910), .B2(n9308), .Y(n9329) );
	mux2i_1 U9480( .A0(n9309), .A1(n9310), .S(n6587), .Y(n9292) );
	nor2_1 U9481( .A(n9322), .B(n9306), .Y(n9310) );
	nor2_1 U9482( .A(n6662), .B(n9321), .Y(n9306) );
	nor2_1 U9483( .A(n9322), .B(n6662), .Y(n9309) );
	o221ai_1 U9484( .A1(n6721), .A2(n5344), .B1(n6748), .B2(n5554), .C1(n9332), .Y(n6662) );
	nand2_1 U9485( .A(n7660), .B(g7052), .Y(n9332) );
	a21oi_1 U9486( .A1(n9323), .A2(n9333), .B1(RST), .Y(n4187) );
	o221ai_1 U9487( .A1(n9307), .A2(n9293), .B1(g1909), .B2(n9308), .C1(n9281), .Y(n9333) );
	nand2_1 U9488( .A(n9334), .B(n9328), .Y(n9293) );
	inv_1 U9489( .A(n9322), .Y(n9328) );
	mux2i_1 U9490( .A0(n6653), .A1(n9315), .S(n6590), .Y(n9334) );
	o21ai_0 U9491( .A1(n9335), .A2(n9322), .B1(n9303), .Y(n9323) );
	inv_1 U9492( .A(n9331), .Y(n9335) );
	o221ai_1 U9493( .A1(n7522), .A2(n6598), .B1(n7499), .B2(n6597), .C1(n9336), .Y(n9331) );
	a21oi_1 U9494( .A1(g7229), .A2(n6560), .B1(n9321), .Y(n9336) );
	inv_1 U9495( .A(n7521), .Y(n6560) );
	o21ai_0 U9496( .A1(RST), .A2(n9337), .B1(n9338), .Y(n4186) );
	nand4_1 U9497( .A(n9865), .B(n9339), .C(n9340), .D(n6098), .Y(n9338) );
	a221oi_1 U9498( .A1(n7590), .A2(n9341), .B1(n7292), .B2(n9342), .C1(n9343), .Y(n9337) );
	and4_1 U9499( .A(g3229), .B(n9866), .C(n9340), .D(n9339), .X(n9343) );
	inv_1 U9500( .A(n9344), .Y(n9340) );
	xor2_1 U9501( .A(n9345), .B(n9346), .X(n9342) );
	xor2_1 U9502( .A(n9347), .B(n9348), .X(n9341) );
	xor2_1 U9503( .A(n9349), .B(n9350), .X(n9348) );
	xor2_1 U9504( .A(n9351), .B(n9352), .X(n9350) );
	xor2_1 U9505( .A(n9353), .B(n9354), .X(n9349) );
	xor2_1 U9506( .A(n9355), .B(n9356), .X(n9347) );
	xor2_1 U9507( .A(n9357), .B(n9358), .X(n9356) );
	xor2_1 U9508( .A(n9359), .B(n9360), .X(n9355) );
	a21oi_1 U9509( .A1(n9361), .A2(n9362), .B1(RST), .Y(n4185) );
	nand2_1 U9510( .A(n9363), .B(n9346), .Y(n9362) );
	nand2_1 U9511( .A(n9364), .B(n9365), .Y(n9346) );
	mux2i_1 U9512( .A0(n7812), .A1(n9366), .S(n7205), .Y(n9364) );
	o221ai_1 U9513( .A1(n9367), .A2(n9352), .B1(g1223), .B2(n9344), .C1(n9339), .Y(n9361) );
	mux2i_1 U9514( .A0(n9368), .A1(n9369), .S(n7209), .Y(n9352) );
	a21oi_1 U9515( .A1(n9370), .A2(n9371), .B1(RST), .Y(n4184) );
	nand2_1 U9516( .A(n9363), .B(n9345), .Y(n9371) );
	nand2_1 U9517( .A(n9372), .B(n9373), .Y(n9345) );
	mux2i_1 U9518( .A0(n7803), .A1(n9374), .S(n7204), .Y(n9372) );
	o221ai_1 U9519( .A1(n9367), .A2(n9353), .B1(g1222), .B2(n9344), .C1(n9339), .Y(n9370) );
	nand2_1 U9520( .A(n9375), .B(n9373), .Y(n9353) );
	mux2i_1 U9521( .A0(n7803), .A1(n9374), .S(n7199), .Y(n9375) );
	o21ai_0 U9522( .A1(n9376), .A2(n9377), .B1(n9378), .Y(n4183) );
	o22ai_1 U9523( .A1(n9367), .A2(n9358), .B1(g1220), .B2(n9344), .Y(n9377) );
	nand2_1 U9524( .A(n9379), .B(n9365), .Y(n9358) );
	a21oi_1 U9525( .A1(n7812), .A2(n9380), .B1(n9381), .Y(n9365) );
	mux2i_1 U9526( .A0(n9366), .A1(n7812), .S(n7203), .Y(n9379) );
	o21ai_0 U9527( .A1(n9376), .A2(n9382), .B1(n9378), .Y(n4182) );
	o22ai_1 U9528( .A1(n9367), .A2(n9357), .B1(g1219), .B2(n9344), .Y(n9382) );
	nand2_1 U9529( .A(n9383), .B(n9373), .Y(n9357) );
	a21oi_1 U9530( .A1(n7803), .A2(n9380), .B1(n9381), .Y(n9373) );
	mux2i_1 U9531( .A0(n7803), .A1(n9374), .S(n7211), .Y(n9383) );
	a21oi_1 U9532( .A1(n9384), .A2(n9385), .B1(RST), .Y(n4181) );
	o221ai_1 U9533( .A1(n9367), .A2(n9351), .B1(g1218), .B2(n9344), .C1(n9339), .Y(n9385) );
	mux2i_1 U9534( .A0(n9368), .A1(n9369), .S(n7198), .Y(n9351) );
	o21ai_0 U9535( .A1(n9376), .A2(n9386), .B1(n9387), .Y(n4180) );
	o22ai_1 U9536( .A1(n9367), .A2(n9360), .B1(g1217), .B2(n9344), .Y(n9386) );
	nand2_1 U9537( .A(n9388), .B(n9389), .Y(n9360) );
	mux2i_1 U9538( .A0(n7803), .A1(n9374), .S(n7213), .Y(n9388) );
	o21ai_0 U9539( .A1(n9376), .A2(n9390), .B1(n9387), .Y(n4179) );
	and2_0 U9540( .A(n9378), .B(n9391), .X(n9387) );
	nand3_1 U9541( .A(n44), .B(n9392), .C(n9363), .Y(n9391) );
	inv_1 U9542( .A(n8987), .Y(n44) );
	nand2_1 U9543( .A(g1186), .B(n5742), .Y(n8987) );
	nand3_1 U9544( .A(n9393), .B(n5740), .C(n9363), .Y(n9378) );
	inv_1 U9545( .A(n9394), .Y(n9393) );
	o22ai_1 U9546( .A1(n9367), .A2(n9354), .B1(g1216), .B2(n9344), .Y(n9390) );
	mux2i_1 U9547( .A0(n9368), .A1(n9369), .S(n7210), .Y(n9354) );
	nor2_1 U9548( .A(n9381), .B(n9366), .Y(n9369) );
	nor2_1 U9549( .A(n7812), .B(n9380), .Y(n9366) );
	nor2_1 U9550( .A(n9381), .B(n7812), .Y(n9368) );
	o221ai_1 U9551( .A1(n7871), .A2(n5345), .B1(n7898), .B2(n5555), .C1(n9395), .Y(n7812) );
	nand2_1 U9552( .A(n7662), .B(g6750), .Y(n9395) );
	nand2_1 U9553( .A(n9339), .B(n5742), .Y(n9376) );
	a21oi_1 U9554( .A1(n9384), .A2(n9396), .B1(RST), .Y(n4178) );
	o221ai_1 U9555( .A1(n9367), .A2(n9359), .B1(g1215), .B2(n9344), .C1(n9339), .Y(n9396) );
	nand2_1 U9556( .A(n9367), .B(n9394), .Y(n9344) );
	nand2_1 U9557( .A(n9397), .B(n9389), .Y(n9359) );
	inv_1 U9558( .A(n9381), .Y(n9389) );
	mux2i_1 U9559( .A0(n7803), .A1(n9374), .S(n7214), .Y(n9397) );
	nor2_1 U9560( .A(n7803), .B(n9380), .Y(n9374) );
	o221ai_1 U9561( .A1(n7871), .A2(n5346), .B1(n7898), .B2(n5556), .C1(n9398), .Y(n7803) );
	nand2_1 U9562( .A(n7663), .B(g6750), .Y(n9398) );
	o21ai_0 U9563( .A1(n9399), .A2(n9381), .B1(n9363), .Y(n9384) );
	nor2_1 U9564( .A(n9400), .B(n9339), .Y(n9363) );
	a21oi_1 U9565( .A1(n5517), .A2(n7788), .B1(n7292), .Y(n9339) );
	inv_1 U9566( .A(n7590), .Y(n7788) );
	inv_1 U9567( .A(n9367), .Y(n9400) );
	a21oi_1 U9568( .A1(n7919), .A2(n5517), .B1(n7590), .Y(n9367) );
	inv_1 U9569( .A(n7292), .Y(n7919) );
	nand2_1 U9570( .A(n9394), .B(g1186), .Y(n9381) );
	nor3_1 U9571( .A(n7288), .B(g1249), .C(n9401), .Y(n9394) );
	inv_1 U9572( .A(n9392), .Y(n9399) );
	o221ai_1 U9573( .A1(n7546), .A2(n7746), .B1(n7523), .B2(n7253), .C1(n9402), .Y(n9392) );
	a21oi_1 U9574( .A1(g6979), .A2(n7183), .B1(n9380), .Y(n9402) );
	and4_1 U9575( .A(n9403), .B(n9404), .C(n9405), .D(n9406), .X(n9380) );
	and3_1 U9576( .A(n7211), .B(n7199), .C(n7204), .X(n9406) );
	o221ai_1 U9577( .A1(n7524), .A2(n7746), .B1(n7525), .B2(n7253), .C1(n9407), .Y(n7204) );
	nand2_1 U9578( .A(g6979), .B(n5453), .Y(n9407) );
	o221ai_1 U9579( .A1(n7530), .A2(n7746), .B1(n7531), .B2(n7253), .C1(n9408), .Y(n7199) );
	nand2_1 U9580( .A(g6979), .B(n5454), .Y(n9408) );
	o221ai_1 U9581( .A1(n7532), .A2(n7746), .B1(n7533), .B2(n7253), .C1(n9409), .Y(n7211) );
	nand2_1 U9582( .A(g6979), .B(n5455), .Y(n9409) );
	nor3_1 U9583( .A(n9410), .B(n9411), .C(n7203), .Y(n9405) );
	a221oi_1 U9584( .A1(n7764), .A2(g7161), .B1(n7763), .B2(n7238), .C1(n9412), .Y(n7203) );
	nor2_1 U9585( .A(n7748), .B(n10035), .Y(n9412) );
	inv_1 U9586( .A(g6979), .Y(n7748) );
	inv_1 U9587( .A(n7529), .Y(n7763) );
	inv_1 U9588( .A(n7528), .Y(n7764) );
	inv_1 U9589( .A(n7205), .Y(n9411) );
	o221ai_1 U9590( .A1(n7526), .A2(n7746), .B1(n7527), .B2(n7253), .C1(n9413), .Y(n7205) );
	nand2_1 U9591( .A(g6979), .B(n5456), .Y(n9413) );
	a222oi_1 U9592( .A1(n7238), .A2(n7168), .B1(g6979), .B2(n5544), .C1(g7161), .C2(n5335), .Y(n9410) );
	inv_1 U9593( .A(n7317), .Y(n7168) );
	nor3_1 U9594( .A(n7210), .B(n9414), .C(n7198), .Y(n9404) );
	o221ai_1 U9595( .A1(n7541), .A2(n7746), .B1(n7542), .B2(n7253), .C1(n9415), .Y(n7198) );
	nand2_1 U9596( .A(g6979), .B(n5457), .Y(n9415) );
	inv_1 U9597( .A(n9416), .Y(n9414) );
	o211ai_1 U9598( .A1(n7253), .A2(n9867), .B1(n7186), .C1(n7185), .Y(n9416) );
	nand2_1 U9599( .A(g7161), .B(n7217), .Y(n7185) );
	inv_1 U9600( .A(n7534), .Y(n7217) );
	nand2_1 U9601( .A(g6979), .B(n5458), .Y(n7186) );
	o221ai_1 U9602( .A1(n7537), .A2(n7746), .B1(n7538), .B2(n7253), .C1(n9417), .Y(n7210) );
	nand2_1 U9603( .A(g6979), .B(n5459), .Y(n9417) );
	nor3_1 U9604( .A(n7214), .B(n7209), .C(n7213), .Y(n9403) );
	o221ai_1 U9605( .A1(n7539), .A2(n7746), .B1(n7540), .B2(n7253), .C1(n9418), .Y(n7213) );
	nand2_1 U9606( .A(g6979), .B(n5460), .Y(n9418) );
	o221ai_1 U9607( .A1(n7543), .A2(n7746), .B1(n7544), .B2(n7253), .C1(n9419), .Y(n7209) );
	nand2_1 U9608( .A(g6979), .B(n5461), .Y(n9419) );
	o221ai_1 U9609( .A1(n7535), .A2(n7746), .B1(n7536), .B2(n7253), .C1(n9420), .Y(n7214) );
	nand2_1 U9610( .A(g6979), .B(n5462), .Y(n9420) );
	inv_1 U9611( .A(n7545), .Y(n7183) );
	inv_1 U9612( .A(n7238), .Y(n7253) );
	inv_1 U9613( .A(g7161), .Y(n7746) );
	o21ai_0 U9614( .A1(RST), .A2(n9421), .B1(n9422), .Y(n4177) );
	nand4_1 U9615( .A(n9868), .B(n9423), .C(n9424), .D(n6098), .Y(n9422) );
	nor2_1 U9616( .A(g3229), .B(RST), .Y(n6098) );
	a221oi_1 U9617( .A1(n7591), .A2(n9425), .B1(n7293), .B2(n9426), .C1(n9427), .Y(n9421) );
	and4_1 U9618( .A(g3229), .B(n9869), .C(n9424), .D(n9423), .X(n9427) );
	xor2_1 U9619( .A(n9428), .B(n9429), .X(n9426) );
	xor2_1 U9620( .A(n9430), .B(n9431), .X(n9425) );
	xor2_1 U9621( .A(n9432), .B(n9433), .X(n9431) );
	xor2_1 U9622( .A(n9434), .B(n9435), .X(n9433) );
	xor2_1 U9623( .A(n9436), .B(n9437), .X(n9432) );
	xor2_1 U9624( .A(n9438), .B(n9439), .X(n9430) );
	xor2_1 U9625( .A(n9440), .B(n9441), .X(n9439) );
	xor2_1 U9626( .A(n9442), .B(n9443), .X(n9438) );
	a21oi_1 U9627( .A1(n9444), .A2(n9445), .B1(RST), .Y(n4176) );
	nand2_1 U9628( .A(n9446), .B(n9429), .Y(n9445) );
	nand2_1 U9629( .A(n9447), .B(n9448), .Y(n9429) );
	mux2i_1 U9630( .A0(n8441), .A1(n9449), .S(n8362), .Y(n9447) );
	o221ai_1 U9631( .A1(n9450), .A2(n9434), .B1(g537), .B2(n9451), .C1(n9423), .Y(n9444) );
	mux2i_1 U9632( .A0(n9452), .A1(n9453), .S(n8366), .Y(n9434) );
	a21oi_1 U9633( .A1(n9454), .A2(n9455), .B1(RST), .Y(n4175) );
	nand2_1 U9634( .A(n9446), .B(n9428), .Y(n9455) );
	nand2_1 U9635( .A(n9456), .B(n9457), .Y(n9428) );
	mux2i_1 U9636( .A0(n8432), .A1(n9458), .S(n8361), .Y(n9456) );
	o221ai_1 U9637( .A1(n9450), .A2(n9436), .B1(g536), .B2(n9451), .C1(n9423), .Y(n9454) );
	nand2_1 U9638( .A(n9459), .B(n9457), .Y(n9436) );
	mux2i_1 U9639( .A0(n8432), .A1(n9458), .S(n8356), .Y(n9459) );
	o21ai_0 U9640( .A1(n9460), .A2(n9461), .B1(n9462), .Y(n4174) );
	o22ai_1 U9641( .A1(n9450), .A2(n9441), .B1(g534), .B2(n9451), .Y(n9461) );
	nand2_1 U9642( .A(n9463), .B(n9448), .Y(n9441) );
	a21oi_1 U9643( .A1(n8441), .A2(n9464), .B1(n9465), .Y(n9448) );
	mux2i_1 U9644( .A0(n9449), .A1(n8441), .S(n8360), .Y(n9463) );
	o21ai_0 U9645( .A1(n9460), .A2(n9466), .B1(n9462), .Y(n4173) );
	o22ai_1 U9646( .A1(n9450), .A2(n9440), .B1(g533), .B2(n9451), .Y(n9466) );
	nand2_1 U9647( .A(n9467), .B(n9457), .Y(n9440) );
	a21oi_1 U9648( .A1(n8432), .A2(n9464), .B1(n9465), .Y(n9457) );
	mux2i_1 U9649( .A0(n8432), .A1(n9458), .S(n8368), .Y(n9467) );
	a21oi_1 U9650( .A1(n9468), .A2(n9469), .B1(RST), .Y(n4172) );
	o221ai_1 U9651( .A1(n9450), .A2(n9437), .B1(g532), .B2(n9451), .C1(n9423), .Y(n9469) );
	mux2i_1 U9652( .A0(n9452), .A1(n9453), .S(n8355), .Y(n9437) );
	o21ai_0 U9653( .A1(n9460), .A2(n9470), .B1(n9471), .Y(n4171) );
	o22ai_1 U9654( .A1(n9450), .A2(n9443), .B1(g531), .B2(n9451), .Y(n9470) );
	nand2_1 U9655( .A(n9472), .B(n9473), .Y(n9443) );
	mux2i_1 U9656( .A0(n8432), .A1(n9458), .S(n8370), .Y(n9472) );
	o21ai_0 U9657( .A1(n9460), .A2(n9474), .B1(n9471), .Y(n4170) );
	and2_0 U9658( .A(n9462), .B(n9475), .X(n9471) );
	nand3_1 U9659( .A(n35), .B(n9476), .C(n9446), .Y(n9475) );
	nand3_1 U9660( .A(n9477), .B(n5740), .C(n9446), .Y(n9462) );
	o22ai_1 U9661( .A1(n9450), .A2(n9435), .B1(g530), .B2(n9451), .Y(n9474) );
	mux2i_1 U9662( .A0(n9452), .A1(n9453), .S(n8367), .Y(n9435) );
	nor2_1 U9663( .A(n9465), .B(n9449), .Y(n9453) );
	nor2_1 U9664( .A(n8441), .B(n9464), .Y(n9449) );
	nor2_1 U9665( .A(n9465), .B(n8441), .Y(n9452) );
	o221ai_1 U9666( .A1(n8500), .A2(n5347), .B1(n8527), .B2(n5557), .C1(n9478), .Y(n8441) );
	nand2_1 U9667( .A(n7664), .B(g6485), .Y(n9478) );
	nand2_1 U9668( .A(n9423), .B(n5743), .Y(n9460) );
	a21oi_1 U9669( .A1(n9468), .A2(n9479), .B1(RST), .Y(n4169) );
	o221ai_1 U9670( .A1(n9450), .A2(n9442), .B1(g529), .B2(n9451), .C1(n9423), .Y(n9479) );
	inv_1 U9671( .A(n9424), .Y(n9451) );
	nor2_1 U9672( .A(n9480), .B(n9477), .Y(n9424) );
	nand2_1 U9673( .A(n9481), .B(n9473), .Y(n9442) );
	mux2i_1 U9674( .A0(n8432), .A1(n9458), .S(n8371), .Y(n9481) );
	nor2_1 U9675( .A(n8432), .B(n9464), .Y(n9458) );
	o221ai_1 U9676( .A1(n8500), .A2(n5348), .B1(n8527), .B2(n5558), .C1(n9482), .Y(n8432) );
	nand2_1 U9677( .A(n7665), .B(g6485), .Y(n9482) );
	o21ai_0 U9678( .A1(n9483), .A2(n9465), .B1(n9446), .Y(n9468) );
	nor2_1 U9679( .A(n9480), .B(n9423), .Y(n9446) );
	a21oi_1 U9680( .A1(n5518), .A2(n8417), .B1(n7293), .Y(n9423) );
	inv_1 U9681( .A(n7591), .Y(n8417) );
	inv_1 U9682( .A(n9450), .Y(n9480) );
	a21oi_1 U9683( .A1(n8548), .A2(n5518), .B1(n7591), .Y(n9450) );
	inv_1 U9684( .A(n7293), .Y(n8548) );
	inv_1 U9685( .A(n9473), .Y(n9465) );
	nor2_1 U9686( .A(n9477), .B(n9484), .Y(n9473) );
	inv_1 U9687( .A(g499), .Y(n9484) );
	o211ai_1 U9688( .A1(g499), .A2(n8495), .B1(n8998), .C1(n9485), .Y(n9477) );
	nor2_1 U9689( .A(n7272), .B(g563), .Y(n9485) );
	inv_1 U9690( .A(n9476), .Y(n9483) );
	o221ai_1 U9691( .A1(n7570), .A2(n8379), .B1(n7547), .B2(n8378), .C1(n9486), .Y(n9476) );
	a21oi_1 U9692( .A1(g6677), .A2(n8340), .B1(n9464), .Y(n9486) );
	and4_1 U9693( .A(n9487), .B(n9488), .C(n9489), .D(n9490), .X(n9464) );
	and3_1 U9694( .A(n8368), .B(n8356), .C(n8361), .X(n9490) );
	o221ai_1 U9695( .A1(n7548), .A2(n8379), .B1(n7549), .B2(n8378), .C1(n9491), .Y(n8361) );
	nand2_1 U9696( .A(g6677), .B(n5463), .Y(n9491) );
	o221ai_1 U9697( .A1(n7554), .A2(n8379), .B1(n7555), .B2(n8378), .C1(n9492), .Y(n8356) );
	nand2_1 U9698( .A(g6677), .B(n5464), .Y(n9492) );
	o221ai_1 U9699( .A1(n7556), .A2(n8379), .B1(n7557), .B2(n8378), .C1(n9493), .Y(n8368) );
	nand2_1 U9700( .A(g6677), .B(n5465), .Y(n9493) );
	nor3_1 U9701( .A(n9494), .B(n9495), .C(n8360), .Y(n9489) );
	a221oi_1 U9702( .A1(n8397), .A2(g6911), .B1(n8396), .B2(n7239), .C1(n9496), .Y(n8360) );
	nor2_1 U9703( .A(n8381), .B(n10036), .Y(n9496) );
	inv_1 U9704( .A(g6677), .Y(n8381) );
	inv_1 U9705( .A(n7553), .Y(n8396) );
	inv_1 U9706( .A(n7552), .Y(n8397) );
	inv_1 U9707( .A(n8362), .Y(n9495) );
	o221ai_1 U9708( .A1(n7550), .A2(n8379), .B1(n7551), .B2(n8378), .C1(n9497), .Y(n8362) );
	nand2_1 U9709( .A(g6677), .B(n5466), .Y(n9497) );
	a222oi_1 U9710( .A1(n7239), .A2(n8325), .B1(g6677), .B2(n5545), .C1(g6911), .C2(n5336), .Y(n9494) );
	inv_1 U9711( .A(n7318), .Y(n8325) );
	nor3_1 U9712( .A(n8367), .B(n9498), .C(n8355), .Y(n9488) );
	o221ai_1 U9713( .A1(n7565), .A2(n8379), .B1(n7566), .B2(n8378), .C1(n9499), .Y(n8355) );
	nand2_1 U9714( .A(g6677), .B(n5467), .Y(n9499) );
	inv_1 U9715( .A(n9500), .Y(n9498) );
	o211ai_1 U9716( .A1(n8378), .A2(n9870), .B1(n8343), .C1(n8342), .Y(n9500) );
	nand2_1 U9717( .A(g6911), .B(n8374), .Y(n8342) );
	inv_1 U9718( .A(n7558), .Y(n8374) );
	nand2_1 U9719( .A(g6677), .B(n5468), .Y(n8343) );
	o221ai_1 U9720( .A1(n7561), .A2(n8379), .B1(n7562), .B2(n8378), .C1(n9501), .Y(n8367) );
	nand2_1 U9721( .A(g6677), .B(n5469), .Y(n9501) );
	nor3_1 U9722( .A(n8371), .B(n8366), .C(n8370), .Y(n9487) );
	o221ai_1 U9723( .A1(n7563), .A2(n8379), .B1(n7564), .B2(n8378), .C1(n9502), .Y(n8370) );
	nand2_1 U9724( .A(g6677), .B(n5470), .Y(n9502) );
	o221ai_1 U9725( .A1(n7567), .A2(n8379), .B1(n7568), .B2(n8378), .C1(n9503), .Y(n8366) );
	nand2_1 U9726( .A(g6677), .B(n5471), .Y(n9503) );
	o221ai_1 U9727( .A1(n7559), .A2(n8379), .B1(n7560), .B2(n8378), .C1(n9504), .Y(n8371) );
	nand2_1 U9728( .A(g6677), .B(n5472), .Y(n9504) );
	inv_1 U9729( .A(n7569), .Y(n8340) );
	inv_1 U9730( .A(n7239), .Y(n8378) );
	inv_1 U9731( .A(g6911), .Y(n8379) );
	and2_0 U9732( .A(g2640), .B(n5763), .X(n4168) );
	and2_0 U9733( .A(g2462), .B(n5763), .X(n4167) );
	and2_0 U9734( .A(g2447), .B(n5763), .X(n4166) );
	and2_0 U9735( .A(g2417), .B(n5763), .X(n4165) );
	and2_0 U9736( .A(g1946), .B(n5763), .X(n4164) );
	and2_0 U9737( .A(g1768), .B(n5763), .X(n4163) );
	and2_0 U9738( .A(g1753), .B(n5763), .X(n4162) );
	and2_0 U9739( .A(g1723), .B(n5763), .X(n4161) );
	a221oi_1 U9740( .A1(n9505), .A2(n9506), .B1(n6839), .B2(n7075), .C1(RST), .Y(n4160) );
	and4_1 U9741( .A(n6979), .B(n7034), .C(n7133), .D(n9507), .X(n7075) );
	nor3_1 U9742( .A(n7029), .B(n7043), .C(n6976), .Y(n9507) );
	and4_1 U9743( .A(n7049), .B(n6996), .C(n9508), .D(n7021), .X(n7133) );
	inv_1 U9744( .A(n7016), .Y(n7021) );
	nor2_1 U9745( .A(n7009), .B(n6994), .Y(n9508) );
	inv_1 U9746( .A(n6995), .Y(n6996) );
	inv_1 U9747( .A(n7040), .Y(n7049) );
	nor4_1 U9748( .A(n9509), .B(n9510), .C(n6337), .D(n9133), .Y(n9506) );
	xor2_1 U9749( .A(n7700), .B(n7043), .X(n9510) );
	o221ai_1 U9750( .A1(n6904), .A2(n5530), .B1(n6903), .B2(n7044), .C1(n9511), .Y(n7043) );
	nand2_1 U9751( .A(n9936), .B(g6573), .Y(n9511) );
	inv_1 U9752( .A(n7682), .Y(n7044) );
	nand3_1 U9753( .A(n9512), .B(n9513), .C(n9514), .Y(n9509) );
	xnor2_1 U9754( .A(n9967), .B(n7040), .Y(n9514) );
	o221ai_1 U9755( .A1(n6904), .A2(n5396), .B1(n6903), .B2(n7050), .C1(n9515), .Y(n7040) );
	nand2_1 U9756( .A(n9939), .B(g6573), .Y(n9515) );
	inv_1 U9757( .A(n7681), .Y(n7050) );
	xnor2_1 U9758( .A(n10086), .B(n7016), .Y(n9513) );
	o21ai_0 U9759( .A1(n6903), .A2(n7017), .B1(n9516), .Y(n7016) );
	a22oi_1 U9760( .A1(n9941), .A2(g6573), .B1(n9940), .B2(g6782), .Y(n9516) );
	inv_1 U9761( .A(n7683), .Y(n7017) );
	xnor2_1 U9762( .A(n10088), .B(n6976), .Y(n9512) );
	o21ai_0 U9763( .A1(n6903), .A2(n6962), .B1(n9517), .Y(n6976) );
	a22oi_1 U9764( .A1(n9938), .A2(g6573), .B1(n9937), .B2(g6782), .Y(n9517) );
	inv_1 U9765( .A(n7684), .Y(n6962) );
	nor4_1 U9766( .A(n9518), .B(n9519), .C(n9520), .D(n9521), .Y(n9505) );
	xnor2_1 U9767( .A(n7710), .B(n7024), .Y(n9521) );
	inv_1 U9768( .A(n7029), .Y(n7024) );
	o221ai_1 U9769( .A1(n6904), .A2(n5531), .B1(n6903), .B2(n7026), .C1(n9522), .Y(n7029) );
	nand2_1 U9770( .A(n9947), .B(g6573), .Y(n9522) );
	inv_1 U9771( .A(n7678), .Y(n7026) );
	xnor2_1 U9772( .A(n10085), .B(n7034), .Y(n9520) );
	inv_1 U9773( .A(n7032), .Y(n7034) );
	o221ai_1 U9774( .A1(n6904), .A2(n5532), .B1(n6903), .B2(n7035), .C1(n9523), .Y(n7032) );
	nand2_1 U9775( .A(n9949), .B(g6573), .Y(n9523) );
	inv_1 U9776( .A(n7686), .Y(n7035) );
	xnor2_1 U9777( .A(n7308), .B(n6979), .Y(n9519) );
	inv_1 U9778( .A(n6989), .Y(n6979) );
	o221ai_1 U9779( .A1(n6904), .A2(n5533), .B1(n6903), .B2(n6981), .C1(n9524), .Y(n6989) );
	nand2_1 U9780( .A(n9948), .B(g6573), .Y(n9524) );
	inv_1 U9781( .A(n7687), .Y(n6981) );
	nand3_1 U9782( .A(n9525), .B(n9526), .C(n9527), .Y(n9518) );
	xnor2_1 U9783( .A(n7697), .B(n7009), .Y(n9527) );
	o21ai_0 U9784( .A1(n6903), .A2(n7010), .B1(n9528), .Y(n7009) );
	a22oi_1 U9785( .A1(n9944), .A2(g6573), .B1(n9943), .B2(g6782), .Y(n9528) );
	inv_1 U9786( .A(n7679), .Y(n7010) );
	xnor2_1 U9787( .A(n7706), .B(n6994), .Y(n9526) );
	o21ai_0 U9788( .A1(n6903), .A2(n6997), .B1(n9529), .Y(n6994) );
	a22oi_1 U9789( .A1(n9946), .A2(g6573), .B1(n9945), .B2(g6782), .Y(n9529) );
	inv_1 U9790( .A(n7685), .Y(n6997) );
	xnor2_1 U9791( .A(n10087), .B(n6995), .Y(n9525) );
	o221ai_1 U9792( .A1(n6904), .A2(n5534), .B1(n6903), .B2(n7003), .C1(n9530), .Y(n6995) );
	nand2_1 U9793( .A(n9942), .B(g6573), .Y(n9530) );
	inv_1 U9794( .A(n7680), .Y(n7003) );
	inv_1 U9795( .A(n7229), .Y(n6903) );
	and2_0 U9796( .A(g1252), .B(n5763), .X(n4159) );
	and2_0 U9797( .A(g1074), .B(n5763), .X(n4158) );
	and2_0 U9798( .A(g1059), .B(n5763), .X(n4157) );
	and2_0 U9799( .A(g1029), .B(n5763), .X(n4156) );
	a221oi_1 U9800( .A1(n9531), .A2(n9532), .B1(n7986), .B2(n8231), .C1(RST), .Y(n4155) );
	and4_1 U9801( .A(n8124), .B(n8185), .C(n8290), .D(n9533), .X(n8231) );
	nor3_1 U9802( .A(n8217), .B(n8194), .C(n8218), .Y(n9533) );
	and4_1 U9803( .A(n8196), .B(n8133), .C(n9534), .D(n8163), .X(n8290) );
	inv_1 U9804( .A(n8161), .Y(n8163) );
	nor2_1 U9805( .A(n8153), .B(n8134), .Y(n9534) );
	inv_1 U9806( .A(n8228), .Y(n8133) );
	nor4_1 U9807( .A(n9535), .B(n9536), .C(n9537), .D(n9538), .Y(n9532) );
	xnor2_1 U9808( .A(n7711), .B(n8171), .Y(n9538) );
	inv_1 U9809( .A(n8217), .Y(n8171) );
	o221ai_1 U9810( .A1(n8049), .A2(n5535), .B1(n8048), .B2(n8172), .C1(n9539), .Y(n8217) );
	nand2_1 U9811( .A(n9815), .B(g6368), .Y(n9539) );
	inv_1 U9812( .A(n7618), .Y(n8172) );
	xnor2_1 U9813( .A(n10001), .B(n8196), .Y(n9537) );
	inv_1 U9814( .A(n8187), .Y(n8196) );
	o221ai_1 U9815( .A1(n8049), .A2(n5397), .B1(n8048), .B2(n8198), .C1(n9540), .Y(n8187) );
	nand2_1 U9816( .A(n9817), .B(g6368), .Y(n9540) );
	inv_1 U9817( .A(n7643), .Y(n8198) );
	xor2_1 U9818( .A(n7707), .B(n8134), .X(n9536) );
	o221ai_1 U9819( .A1(n8049), .A2(n5536), .B1(n8048), .B2(n8138), .C1(n9541), .Y(n8134) );
	nand2_1 U9820( .A(n9816), .B(g6368), .Y(n9541) );
	inv_1 U9821( .A(n7646), .Y(n8138) );
	nand3_1 U9822( .A(n9158), .B(n6131), .C(n9542), .Y(n9535) );
	xnor2_1 U9823( .A(n10004), .B(n8218), .Y(n9542) );
	o21ai_0 U9824( .A1(n8048), .A2(n8107), .B1(n9543), .Y(n8218) );
	a22oi_1 U9825( .A1(n9814), .A2(g6368), .B1(n9813), .B2(g6518), .Y(n9543) );
	inv_1 U9826( .A(n7645), .Y(n8107) );
	inv_1 U9827( .A(n6337), .Y(n6131) );
	nor4_1 U9828( .A(n9544), .B(n9545), .C(n9546), .D(n9547), .Y(n9531) );
	xnor2_1 U9829( .A(n7305), .B(n8124), .Y(n9547) );
	inv_1 U9830( .A(n8132), .Y(n8124) );
	o221ai_1 U9831( .A1(n8049), .A2(n5537), .B1(n8048), .B2(n8125), .C1(n9548), .Y(n8132) );
	nand2_1 U9832( .A(n9822), .B(g6368), .Y(n9548) );
	inv_1 U9833( .A(n7648), .Y(n8125) );
	xnor2_1 U9834( .A(n7701), .B(n8186), .Y(n9546) );
	inv_1 U9835( .A(n8194), .Y(n8186) );
	o221ai_1 U9836( .A1(n8049), .A2(n5538), .B1(n8048), .B2(n8190), .C1(n9549), .Y(n8194) );
	nand2_1 U9837( .A(n9824), .B(g6368), .Y(n9549) );
	inv_1 U9838( .A(n7644), .Y(n8190) );
	xnor2_1 U9839( .A(n10007), .B(n8185), .Y(n9545) );
	inv_1 U9840( .A(n8177), .Y(n8185) );
	o221ai_1 U9841( .A1(n8049), .A2(n5539), .B1(n8048), .B2(n8178), .C1(n9550), .Y(n8177) );
	nand2_1 U9842( .A(n9823), .B(g6368), .Y(n9550) );
	inv_1 U9843( .A(n7647), .Y(n8178) );
	nand3_1 U9844( .A(n9551), .B(n9552), .C(n9553), .Y(n9544) );
	xnor2_1 U9845( .A(n10005), .B(n8228), .Y(n9553) );
	o221ai_1 U9846( .A1(n8049), .A2(n5540), .B1(n8048), .B2(n8146), .C1(n9554), .Y(n8228) );
	nand2_1 U9847( .A(n9820), .B(g6368), .Y(n9554) );
	inv_1 U9848( .A(n7642), .Y(n8146) );
	xnor2_1 U9849( .A(n10006), .B(n8161), .Y(n9552) );
	o221ai_1 U9850( .A1(n8049), .A2(n5541), .B1(n8048), .B2(n8164), .C1(n9555), .Y(n8161) );
	nand2_1 U9851( .A(n9821), .B(g6368), .Y(n9555) );
	inv_1 U9852( .A(n7619), .Y(n8164) );
	xnor2_1 U9853( .A(n7698), .B(n8153), .Y(n9551) );
	o21ai_0 U9854( .A1(n8048), .A2(n8154), .B1(n9556), .Y(n8153) );
	a22oi_1 U9855( .A1(n9819), .A2(g6368), .B1(n9818), .B2(g6518), .Y(n9556) );
	inv_1 U9856( .A(n7641), .Y(n8154) );
	inv_1 U9857( .A(n7231), .Y(n8048) );
	and2_0 U9858( .A(g543), .B(n5763), .X(n4154) );
	and2_0 U9859( .A(g566), .B(n5763), .X(n4153) );
	and2_0 U9860( .A(g387), .B(n5763), .X(n4152) );
	and2_0 U9861( .A(g372), .B(n5762), .X(n4151) );
	and2_0 U9862( .A(g342), .B(n5762), .X(n4150) );
	o21ai_0 U9863( .A1(n9317), .A2(n9557), .B1(n9319), .Y(n4149) );
	nand3_1 U9864( .A(n9558), .B(n5740), .C(n9303), .Y(n9319) );
	nor2_1 U9865( .A(n9559), .B(n9281), .Y(n9303) );
	o22ai_1 U9866( .A1(n9307), .A2(n9297), .B1(g1913), .B2(n9308), .Y(n9557) );
	inv_1 U9867( .A(n9280), .Y(n9308) );
	nor2_1 U9868( .A(n9559), .B(n9558), .Y(n9280) );
	inv_1 U9869( .A(n9560), .Y(n9558) );
	nand2_1 U9870( .A(n9561), .B(n9314), .Y(n9297) );
	a21oi_1 U9871( .A1(n6653), .A2(n9321), .B1(n9322), .Y(n9314) );
	nand2_1 U9872( .A(n9560), .B(g1880), .Y(n9322) );
	nor3_1 U9873( .A(n7289), .B(g1943), .C(n8993), .Y(n9560) );
	mux2i_1 U9874( .A0(n6653), .A1(n9315), .S(n6589), .Y(n9561) );
	nor2_1 U9875( .A(n6653), .B(n9321), .Y(n9315) );
	and4_1 U9876( .A(n9562), .B(n9563), .C(n9564), .D(n9565), .X(n9321) );
	and3_1 U9877( .A(n6589), .B(n6576), .C(n6581), .X(n9565) );
	o221ai_1 U9878( .A1(n7500), .A2(n6598), .B1(n7501), .B2(n6597), .C1(n9566), .Y(n6581) );
	nand2_1 U9879( .A(g7229), .B(n5473), .Y(n9566) );
	o221ai_1 U9880( .A1(n7506), .A2(n6598), .B1(n7507), .B2(n6597), .C1(n9567), .Y(n6576) );
	nand2_1 U9881( .A(g7229), .B(n5474), .Y(n9567) );
	o221ai_1 U9882( .A1(n7508), .A2(n6598), .B1(n7509), .B2(n6597), .C1(n9568), .Y(n6589) );
	nand2_1 U9883( .A(g7229), .B(n5475), .Y(n9568) );
	nor3_1 U9884( .A(n9569), .B(n9570), .C(n6580), .Y(n9564) );
	a221oi_1 U9885( .A1(n6617), .A2(g7357), .B1(n6616), .B2(n7237), .C1(n9571), .Y(n6580) );
	nor2_1 U9886( .A(n6600), .B(n10069), .Y(n9571) );
	inv_1 U9887( .A(g7229), .Y(n6600) );
	inv_1 U9888( .A(n7505), .Y(n6616) );
	inv_1 U9889( .A(n7504), .Y(n6617) );
	inv_1 U9890( .A(n6582), .Y(n9570) );
	o221ai_1 U9891( .A1(n7502), .A2(n6598), .B1(n7503), .B2(n6597), .C1(n9572), .Y(n6582) );
	nand2_1 U9892( .A(g7229), .B(n5476), .Y(n9572) );
	a222oi_1 U9893( .A1(n7237), .A2(n6545), .B1(g7229), .B2(n5546), .C1(g7357), .C2(n5337), .Y(n9569) );
	inv_1 U9894( .A(n7316), .Y(n6545) );
	nor3_1 U9895( .A(n6587), .B(n9573), .C(n6575), .Y(n9563) );
	o221ai_1 U9896( .A1(n7517), .A2(n6598), .B1(n7518), .B2(n6597), .C1(n9574), .Y(n6575) );
	nand2_1 U9897( .A(g7229), .B(n5477), .Y(n9574) );
	inv_1 U9898( .A(n9575), .Y(n9573) );
	o211ai_1 U9899( .A1(n6597), .A2(n9911), .B1(n6563), .C1(n6562), .Y(n9575) );
	nand2_1 U9900( .A(g7357), .B(n6593), .Y(n6562) );
	inv_1 U9901( .A(n7510), .Y(n6593) );
	nand2_1 U9902( .A(g7229), .B(n5478), .Y(n6563) );
	o221ai_1 U9903( .A1(n7513), .A2(n6598), .B1(n7514), .B2(n6597), .C1(n9576), .Y(n6587) );
	nand2_1 U9904( .A(g7229), .B(n5479), .Y(n9576) );
	nor3_1 U9905( .A(n6590), .B(n6586), .C(n6588), .Y(n9562) );
	o221ai_1 U9906( .A1(n7515), .A2(n6598), .B1(n7516), .B2(n6597), .C1(n9577), .Y(n6588) );
	nand2_1 U9907( .A(g7229), .B(n5480), .Y(n9577) );
	o221ai_1 U9908( .A1(n7519), .A2(n6598), .B1(n7520), .B2(n6597), .C1(n9578), .Y(n6586) );
	nand2_1 U9909( .A(g7229), .B(n5481), .Y(n9578) );
	o221ai_1 U9910( .A1(n7511), .A2(n6598), .B1(n7512), .B2(n6597), .C1(n9579), .Y(n6590) );
	nand2_1 U9911( .A(g7229), .B(n5482), .Y(n9579) );
	inv_1 U9912( .A(n7237), .Y(n6597) );
	inv_1 U9913( .A(g7357), .Y(n6598) );
	o221ai_1 U9914( .A1(n6721), .A2(n5349), .B1(n6748), .B2(n5559), .C1(n9580), .Y(n6653) );
	nand2_1 U9915( .A(n7661), .B(g7052), .Y(n9580) );
	inv_1 U9916( .A(n9559), .Y(n9307) );
	o21ai_0 U9917( .A1(n7291), .A2(n9964), .B1(n6638), .Y(n9559) );
	inv_1 U9918( .A(n7589), .Y(n6638) );
	nand2_1 U9919( .A(n9281), .B(n5743), .Y(n9317) );
	inv_1 U9920( .A(n9581), .Y(n9281) );
	o21ai_0 U9921( .A1(n9964), .A2(n7589), .B1(n6771), .Y(n9581) );
	inv_1 U9922( .A(n7291), .Y(n6771) );
	and2_0 U9923( .A(n5763), .B(n6096), .X(n4148) );
	o22ai_1 U9924( .A1(n6755), .A2(n5940), .B1(n9582), .B2(n5994), .Y(n6096) );
	o21ai_0 U9925( .A1(n6101), .A2(n5566), .B1(n9583), .Y(n5994) );
	a22oi_1 U9926( .A1(n7636), .A2(g7302), .B1(n9877), .B2(g7390), .Y(n9583) );
	a21oi_1 U9927( .A1(n7588), .A2(n5944), .B1(n5981), .Y(n9582) );
	inv_1 U9928( .A(n6755), .Y(n5981) );
	o221ai_1 U9929( .A1(n6071), .A2(n5350), .B1(n6101), .B2(n5560), .C1(n9584), .Y(n5944) );
	nand2_1 U9930( .A(n7658), .B(g7302), .Y(n9584) );
	o221ai_1 U9931( .A1(n6071), .A2(n5351), .B1(n6101), .B2(n5561), .C1(n9585), .Y(n5940) );
	nand2_1 U9932( .A(n7659), .B(g7302), .Y(n9585) );
	nor4_1 U9933( .A(n7249), .B(n7254), .C(n9586), .D(n7326), .Y(n6755) );
	or2_0 U9934( .A(n10082), .B(n10083), .X(n9586) );
	and2_0 U9935( .A(g2609), .B(n5762), .X(n4147) );
	and2_0 U9936( .A(g2644), .B(n5762), .X(n4146) );
	and2_0 U9937( .A(g2597), .B(n5762), .X(n4145) );
	and2_0 U9938( .A(g2432), .B(n5762), .X(n4144) );
	and2_0 U9939( .A(g1915), .B(n5762), .X(n4143) );
	and2_0 U9940( .A(g1950), .B(n5762), .X(n4142) );
	and2_0 U9941( .A(g1903), .B(n5762), .X(n4141) );
	and2_0 U9942( .A(g1738), .B(n5762), .X(n4140) );
	and2_0 U9943( .A(g1221), .B(n5762), .X(n4139) );
	and2_0 U9944( .A(g1256), .B(n5762), .X(n4138) );
	and2_0 U9945( .A(g1209), .B(n5762), .X(n4137) );
	and2_0 U9946( .A(g1044), .B(n5762), .X(n4136) );
	and2_0 U9947( .A(g535), .B(n5762), .X(n4135) );
	and2_0 U9948( .A(g570), .B(n5762), .X(n4134) );
	and2_0 U9949( .A(g523), .B(n5762), .X(n4133) );
	and2_0 U9950( .A(g357), .B(n5762), .X(n4132) );
	nor2_1 U9951( .A(n10043), .B(RST), .Y(n4130) );
	nor2_1 U9952( .A(n10044), .B(RST), .Y(n4129) );
	nor2_1 U9953( .A(n10045), .B(RST), .Y(n4128) );
	nor2_1 U9954( .A(n10046), .B(RST), .Y(n4127) );
	nor2_1 U9955( .A(n10047), .B(RST), .Y(n4126) );
	nor2_1 U9956( .A(n10048), .B(RST), .Y(n4125) );
	nor2_1 U9957( .A(n10049), .B(RST), .Y(n4124) );
	nor2_1 U9958( .A(n10050), .B(RST), .Y(n4123) );
	nor2_1 U9959( .A(n10073), .B(RST), .Y(n4122) );
	nor2_1 U9960( .A(n10074), .B(RST), .Y(n4121) );
	nor2_1 U9961( .A(n10075), .B(RST), .Y(n4120) );
	nor2_1 U9962( .A(n10076), .B(RST), .Y(n4119) );
	nor2_1 U9963( .A(n10077), .B(RST), .Y(n4118) );
	nor2_1 U9964( .A(n10078), .B(RST), .Y(n4117) );
	nor2_1 U9965( .A(n10079), .B(RST), .Y(n4116) );
	nor2_1 U9966( .A(n10080), .B(RST), .Y(n4115) );
	nor2_1 U9967( .A(n9993), .B(RST), .Y(n4114) );
	nor2_1 U9968( .A(n9994), .B(RST), .Y(n4113) );
	nor2_1 U9969( .A(n9995), .B(RST), .Y(n4112) );
	nor2_1 U9970( .A(n9996), .B(RST), .Y(n4111) );
	nor2_1 U9971( .A(n9997), .B(RST), .Y(n4110) );
	nor2_1 U9972( .A(n9998), .B(RST), .Y(n4109) );
	nor2_1 U9973( .A(n9999), .B(RST), .Y(n4108) );
	nor2_1 U9974( .A(n10000), .B(RST), .Y(n4107) );
	nor2_1 U9975( .A(n10015), .B(RST), .Y(n4106) );
	nor2_1 U9976( .A(n10016), .B(RST), .Y(n4105) );
	nor2_1 U9977( .A(n10017), .B(RST), .Y(n4104) );
	nor2_1 U9978( .A(n10018), .B(RST), .Y(n4103) );
	nor2_1 U9979( .A(n10019), .B(RST), .Y(n4102) );
	nor2_1 U9980( .A(n10020), .B(RST), .Y(n4101) );
	nor2_1 U9981( .A(n10021), .B(RST), .Y(n4100) );
	nor2_1 U9982( .A(RST), .B(n7235), .Y(n41) );
	nor2_1 U9983( .A(n10022), .B(RST), .Y(n4099) );
	nor2_1 U9984( .A(RST), .B(g25435), .Y(n4098) );
	nor2_1 U9985( .A(RST), .B(g26135), .Y(n4097) );
	mux2i_1 U9986( .A0(n9587), .A1(n9588), .S(n7725), .Y(n4096) );
	nand2_1 U9987( .A(g2581), .B(n5745), .Y(n9588) );
	a22oi_1 U9988( .A1(n9088), .A2(n59), .B1(n68), .B2(n6071), .Y(n9587) );
	and2_0 U9989( .A(g16437), .B(n5761), .X(n68) );
	nor2_1 U9990( .A(n6071), .B(RST), .Y(n59) );
	inv_1 U9991( .A(g7390), .Y(n6071) );
	mux2i_1 U9992( .A0(n9589), .A1(n15018), .S(n7730), .Y(n9088) );
	mux2i_1 U9993( .A0(n9089), .A1(g16399), .S(n6721), .Y(n9589) );
	mux2i_1 U9994( .A0(n9590), .A1(n15150), .S(n7741), .Y(n9089) );
	mux2i_1 U9995( .A0(n9591), .A1(g16355), .S(n7871), .Y(n9590) );
	o22ai_1 U9996( .A1(n7260), .A2(n5789), .B1(n6108), .B2(n9592), .Y(n4095) );
	nand2_1 U9997( .A(g2546), .B(n5745), .Y(n5789) );
	o22ai_1 U9998( .A1(g8167), .A2(n5790), .B1(n5787), .B2(n9592), .Y(n4094) );
	nand2_1 U9999( .A(g2543), .B(n5745), .Y(n5790) );
	o22ai_1 U10000( .A1(g8087), .A2(n5791), .B1(n5788), .B2(n9592), .Y(n4093) );
	inv_1 U10001( .A(n6121), .Y(n9592) );
	nor3_1 U10002( .A(n6187), .B(n6203), .C(n6198), .Y(n6121) );
	nand2_1 U10003( .A(g2540), .B(n5745), .Y(n5791) );
	o22ai_1 U10004( .A1(n7260), .A2(n5792), .B1(n6108), .B2(n6130), .Y(n4092) );
	nand2_1 U10005( .A(n7260), .B(n5745), .Y(n6108) );
	nand2_1 U10006( .A(g2536), .B(n5745), .Y(n5792) );
	o22ai_1 U10007( .A1(g8167), .A2(n5793), .B1(n5787), .B2(n6130), .Y(n4091) );
	nand2_1 U10008( .A(g8167), .B(n5745), .Y(n5787) );
	nand2_1 U10009( .A(g2533), .B(n5745), .Y(n5793) );
	o22ai_1 U10010( .A1(g8087), .A2(n5794), .B1(n5788), .B2(n6130), .Y(n4090) );
	nand3_1 U10011( .A(n6198), .B(n6203), .C(n6245), .Y(n6130) );
	inv_1 U10012( .A(n6187), .Y(n6245) );
	o221ai_1 U10013( .A1(n9892), .A2(n6281), .B1(n7571), .B2(n6264), .C1(n9593), .Y(n6187) );
	nand2_1 U10014( .A(n7780), .B(n6240), .Y(n9593) );
	inv_1 U10015( .A(n7572), .Y(n6240) );
	o221ai_1 U10016( .A1(n9893), .A2(n6281), .B1(n7575), .B2(n6264), .C1(n9594), .Y(n6203) );
	nand2_1 U10017( .A(n7780), .B(n6207), .Y(n9594) );
	inv_1 U10018( .A(n7576), .Y(n6207) );
	o221ai_1 U10019( .A1(n9894), .A2(n6281), .B1(n7573), .B2(n6264), .C1(n9595), .Y(n6198) );
	nand2_1 U10020( .A(n7780), .B(n6189), .Y(n9595) );
	inv_1 U10021( .A(n7574), .Y(n6189) );
	inv_1 U10022( .A(g7264), .Y(n6264) );
	nand2_1 U10023( .A(g8087), .B(n5745), .Y(n5788) );
	nand2_1 U10024( .A(g2530), .B(n5745), .Y(n5794) );
	o22ai_1 U10025( .A1(n7257), .A2(n9596), .B1(n6760), .B2(n9132), .Y(n4089) );
	o22ai_1 U10026( .A1(g8082), .A2(n9597), .B1(n6762), .B2(n9132), .Y(n4088) );
	o22ai_1 U10027( .A1(g8012), .A2(n9598), .B1(n6765), .B2(n9132), .Y(n4087) );
	inv_1 U10028( .A(n6839), .Y(n9132) );
	nor3_1 U10029( .A(n6823), .B(n6828), .C(n6812), .Y(n6839) );
	o22ai_1 U10030( .A1(n7257), .A2(n9599), .B1(n6760), .B2(n9600), .Y(n4086) );
	nand2_1 U10031( .A(n7257), .B(n5745), .Y(n6760) );
	o22ai_1 U10032( .A1(g8082), .A2(n9601), .B1(n6762), .B2(n9600), .Y(n4085) );
	o22ai_1 U10033( .A1(g8012), .A2(n9602), .B1(n6765), .B2(n9600), .Y(n4084) );
	inv_1 U10034( .A(n9133), .Y(n9600) );
	nor3_1 U10035( .A(n6836), .B(n6809), .C(n6812), .Y(n9133) );
	o221ai_1 U10036( .A1(n9933), .A2(n6939), .B1(n7577), .B2(n6774), .C1(n9603), .Y(n6812) );
	nand2_1 U10037( .A(n7782), .B(n6864), .Y(n9603) );
	inv_1 U10038( .A(n7578), .Y(n6864) );
	inv_1 U10039( .A(n6823), .Y(n6809) );
	o221ai_1 U10040( .A1(n9934), .A2(n6939), .B1(n7579), .B2(n6774), .C1(n9604), .Y(n6823) );
	nand2_1 U10041( .A(n7782), .B(n6814), .Y(n9604) );
	inv_1 U10042( .A(n7580), .Y(n6814) );
	inv_1 U10043( .A(n6828), .Y(n6836) );
	o221ai_1 U10044( .A1(n9935), .A2(n6939), .B1(n7581), .B2(n6774), .C1(n9605), .Y(n6828) );
	nand2_1 U10045( .A(n7782), .B(n6832), .Y(n9605) );
	inv_1 U10046( .A(n7582), .Y(n6832) );
	o22ai_1 U10047( .A1(n7258), .A2(n9606), .B1(n7908), .B2(n9607), .Y(n4083) );
	o22ai_1 U10048( .A1(g8007), .A2(n9608), .B1(n7910), .B2(n9607), .Y(n4082) );
	o22ai_1 U10049( .A1(g7961), .A2(n9609), .B1(n7913), .B2(n9607), .Y(n4081) );
	inv_1 U10050( .A(n7986), .Y(n9607) );
	nor3_1 U10051( .A(n7970), .B(n7975), .C(n7958), .Y(n7986) );
	o22ai_1 U10052( .A1(n7258), .A2(n9610), .B1(n7908), .B2(n9158), .Y(n4080) );
	nand2_1 U10053( .A(n7258), .B(n5746), .Y(n7908) );
	o22ai_1 U10054( .A1(g8007), .A2(n9611), .B1(n7910), .B2(n9158), .Y(n4079) );
	o22ai_1 U10055( .A1(g7961), .A2(n9612), .B1(n7913), .B2(n9158), .Y(n4078) );
	nand3_1 U10056( .A(n7970), .B(n7975), .C(n8016), .Y(n9158) );
	inv_1 U10057( .A(n7958), .Y(n8016) );
	o221ai_1 U10058( .A1(n9810), .A2(n7932), .B1(n7463), .B2(n8032), .C1(n9613), .Y(n7958) );
	nand2_1 U10059( .A(n7775), .B(n8012), .Y(n9613) );
	inv_1 U10060( .A(n7464), .Y(n8012) );
	o221ai_1 U10061( .A1(n9811), .A2(n7932), .B1(n7467), .B2(n8032), .C1(n9614), .Y(n7975) );
	nand2_1 U10062( .A(n7775), .B(n7980), .Y(n9614) );
	inv_1 U10063( .A(n7468), .Y(n7980) );
	o221ai_1 U10064( .A1(n9812), .A2(n7932), .B1(n7465), .B2(n8032), .C1(n9615), .Y(n7970) );
	nand2_1 U10065( .A(n7775), .B(n7962), .Y(n9615) );
	inv_1 U10066( .A(n7466), .Y(n7962) );
	o22ai_1 U10067( .A1(n7259), .A2(n9616), .B1(n8537), .B2(n9617), .Y(n4077) );
	o22ai_1 U10068( .A1(g7956), .A2(n9618), .B1(n8539), .B2(n9617), .Y(n4076) );
	o22ai_1 U10069( .A1(g7909), .A2(n9619), .B1(n8542), .B2(n9617), .Y(n4075) );
	inv_1 U10070( .A(n8554), .Y(n9617) );
	nor3_1 U10071( .A(n8617), .B(n8633), .C(n8628), .Y(n8554) );
	o22ai_1 U10072( .A1(n7259), .A2(n9620), .B1(n8537), .B2(n8563), .Y(n4074) );
	nand2_1 U10073( .A(n7259), .B(n5746), .Y(n8537) );
	o22ai_1 U10074( .A1(g7956), .A2(n9621), .B1(n8539), .B2(n8563), .Y(n4073) );
	o22ai_1 U10075( .A1(g7909), .A2(n9622), .B1(n8542), .B2(n8563), .Y(n4072) );
	nand3_1 U10076( .A(n8628), .B(n8633), .C(n8673), .Y(n8563) );
	inv_1 U10077( .A(n8617), .Y(n8673) );
	o221ai_1 U10078( .A1(n9840), .A2(n8709), .B1(n7470), .B2(n8692), .C1(n9623), .Y(n8617) );
	nand2_1 U10079( .A(n7784), .B(n8668), .Y(n9623) );
	inv_1 U10080( .A(n7469), .Y(n8668) );
	o221ai_1 U10081( .A1(n9841), .A2(n8709), .B1(n7474), .B2(n8692), .C1(n9624), .Y(n8633) );
	nand2_1 U10082( .A(n7784), .B(n8637), .Y(n9624) );
	inv_1 U10083( .A(n7473), .Y(n8637) );
	o221ai_1 U10084( .A1(n9842), .A2(n8709), .B1(n7472), .B2(n8692), .C1(n9625), .Y(n8628) );
	nand2_1 U10085( .A(n7784), .B(n8619), .Y(n9625) );
	inv_1 U10086( .A(n7471), .Y(n8619) );
	o22ai_1 U10087( .A1(n7587), .A2(n5795), .B1(n5822), .B2(n9626), .Y(n4071) );
	nand2_1 U10088( .A(g2878), .B(n5746), .Y(n5795) );
	o22ai_1 U10089( .A1(n5820), .A2(n9627), .B1(n5822), .B2(n9628), .Y(n4070) );
	o22ai_1 U10090( .A1(n5820), .A2(n5839), .B1(n5822), .B2(n9629), .Y(n4069) );
	inv_1 U10091( .A(n7598), .Y(n5839) );
	o22ai_1 U10092( .A1(n5820), .A2(n5841), .B1(n5822), .B2(n9630), .Y(n4068) );
	inv_1 U10093( .A(n7605), .Y(n5841) );
	o22ai_1 U10094( .A1(n5820), .A2(n5843), .B1(n5822), .B2(n9631), .Y(n4067) );
	inv_1 U10095( .A(n7599), .Y(n5843) );
	o22ai_1 U10096( .A1(n5820), .A2(n5845), .B1(n5822), .B2(n9632), .Y(n4066) );
	o22ai_1 U10097( .A1(n5820), .A2(n5847), .B1(n5822), .B2(n9633), .Y(n4065) );
	o22ai_1 U10098( .A1(n5820), .A2(n5849), .B1(n5822), .B2(n9634), .Y(n4064) );
	inv_1 U10099( .A(n7607), .Y(n5849) );
	o22ai_1 U10100( .A1(n5820), .A2(n5851), .B1(n5822), .B2(n9635), .Y(n4063) );
	o22ai_1 U10101( .A1(n5820), .A2(n5853), .B1(n5822), .B2(n9636), .Y(n4062) );
	inv_1 U10102( .A(n7280), .Y(n5853) );
	o22ai_1 U10103( .A1(n5820), .A2(n9626), .B1(n5822), .B2(n9637), .Y(n4061) );
	xnor2_1 U10104( .A(n9638), .B(n9007), .Y(n9626) );
	xnor2_1 U10105( .A(n9639), .B(n9640), .Y(n9007) );
	xor2_1 U10106( .A(n9641), .B(n9642), .X(n9640) );
	xnor2_1 U10107( .A(n5831), .B(n7601), .Y(n9642) );
	xnor2_1 U10108( .A(n5827), .B(n7603), .Y(n9641) );
	xor2_1 U10109( .A(n9643), .B(n9644), .X(n9639) );
	xnor2_1 U10110( .A(n5829), .B(n7596), .Y(n9644) );
	xnor2_1 U10111( .A(n7281), .B(n7595), .Y(n9643) );
	o22ai_1 U10112( .A1(n5823), .A2(n5820), .B1(n5822), .B2(n9645), .Y(n4060) );
	inv_1 U10113( .A(n7596), .Y(n5823) );
	o22ai_1 U10114( .A1(n5820), .A2(n5825), .B1(n5822), .B2(n9646), .Y(n4059) );
	inv_1 U10115( .A(n7281), .Y(n5825) );
	o22ai_1 U10116( .A1(n5820), .A2(n5827), .B1(n5822), .B2(n9647), .Y(n4058) );
	inv_1 U10117( .A(n7604), .Y(n5827) );
	o22ai_1 U10118( .A1(n5820), .A2(n5829), .B1(n5822), .B2(n9648), .Y(n4057) );
	inv_1 U10119( .A(n7597), .Y(n5829) );
	o22ai_1 U10120( .A1(n5820), .A2(n5831), .B1(n5822), .B2(n9649), .Y(n4056) );
	inv_1 U10121( .A(n7602), .Y(n5831) );
	o22ai_1 U10122( .A1(n5820), .A2(n5833), .B1(n5822), .B2(n9650), .Y(n4055) );
	inv_1 U10123( .A(n7601), .Y(n5833) );
	o22ai_1 U10124( .A1(n5820), .A2(n5835), .B1(n5822), .B2(n9651), .Y(n4054) );
	inv_1 U10125( .A(n7595), .Y(n5835) );
	o22ai_1 U10126( .A1(n5820), .A2(n5837), .B1(n5822), .B2(n9652), .Y(n4053) );
	inv_1 U10127( .A(n7603), .Y(n5837) );
	o22ai_1 U10128( .A1(n5820), .A2(n9653), .B1(n5822), .B2(n9627), .Y(n4052) );
	xnor2_1 U10129( .A(n9638), .B(n9009), .Y(n9627) );
	xnor2_1 U10130( .A(n9654), .B(n9655), .Y(n9009) );
	xor2_1 U10131( .A(n9656), .B(n9657), .X(n9655) );
	xnor2_1 U10132( .A(n5845), .B(n7605), .Y(n9657) );
	inv_1 U10133( .A(n7606), .Y(n5845) );
	xnor2_1 U10134( .A(n5851), .B(n7607), .Y(n9656) );
	inv_1 U10135( .A(n7608), .Y(n5851) );
	xor2_1 U10136( .A(n9658), .B(n9659), .X(n9654) );
	xnor2_1 U10137( .A(n5847), .B(n7599), .Y(n9659) );
	inv_1 U10138( .A(n7600), .Y(n5847) );
	xnor2_1 U10139( .A(n7280), .B(n7598), .Y(n9658) );
	or2_0 U10140( .A(n5567), .B(g3231), .X(n9638) );
	nand2_1 U10141( .A(n7587), .B(n5746), .Y(n5822) );
	and2_0 U10142( .A(g3232), .B(n5761), .X(n4051) );
	and2_0 U10143( .A(g3212), .B(n5761), .X(n4050) );
	and2_0 U10144( .A(n5762), .B(n9591), .X(n4049) );
	mux2i_1 U10145( .A0(n9660), .A1(n15423), .S(n7744), .Y(n9591) );
	nor2_1 U10146( .A(g6642), .B(g16297), .Y(n9660) );
	o21ai_0 U10147( .A1(RST), .A2(n14891), .B1(n9661), .Y(n4048) );
	o21ai_0 U10148( .A1(RST), .A2(n14915), .B1(n5871), .Y(n4047) );
	inv_1 U10149( .A(n70), .Y(n5871) );
	nor2_1 U10150( .A(n5867), .B(RST), .Y(n70) );
	inv_1 U10151( .A(g3234), .Y(n5867) );
	a211oi_1 U10152( .A1(g7390), .A2(n5415), .B1(n9662), .C1(RST), .Y(n4046) );
	o22ai_1 U10153( .A1(n9881), .A2(n6066), .B1(n7451), .B2(n6101), .Y(n9662) );
	a211oi_1 U10154( .A1(g7390), .A2(n5416), .B1(n9663), .C1(RST), .Y(n4045) );
	o22ai_1 U10155( .A1(n9879), .A2(n6066), .B1(n7459), .B2(n6101), .Y(n9663) );
	a211oi_1 U10156( .A1(g7390), .A2(n5417), .B1(n9664), .C1(RST), .Y(n4044) );
	o22ai_1 U10157( .A1(n9880), .A2(n6066), .B1(n7453), .B2(n6101), .Y(n9664) );
	nor2_1 U10158( .A(RST), .B(n6069), .Y(n4043) );
	o21ai_0 U10159( .A1(n6101), .A2(n15635), .B1(n9665), .Y(n6069) );
	a22oi_1 U10160( .A1(g2641), .A2(g7390), .B1(n9878), .B2(g7302), .Y(n9665) );
	nor2_1 U10161( .A(RST), .B(n6074), .Y(n4042) );
	o21ai_0 U10162( .A1(n6101), .A2(n15627), .B1(n9666), .Y(n6074) );
	a22oi_1 U10163( .A1(g2645), .A2(g7390), .B1(n9882), .B2(g7302), .Y(n9666) );
	inv_1 U10164( .A(n7224), .Y(n6101) );
	a211oi_1 U10165( .A1(g7194), .A2(n5418), .B1(n9667), .C1(RST), .Y(n4041) );
	o22ai_1 U10166( .A1(n9929), .A2(n6716), .B1(n7452), .B2(n6748), .Y(n9667) );
	a211oi_1 U10167( .A1(g7194), .A2(n5419), .B1(n9668), .C1(RST), .Y(n4040) );
	o22ai_1 U10168( .A1(n9926), .A2(n6716), .B1(n7460), .B2(n6748), .Y(n9668) );
	a211oi_1 U10169( .A1(g7194), .A2(n5420), .B1(n9669), .C1(RST), .Y(n4039) );
	o22ai_1 U10170( .A1(n9928), .A2(n6716), .B1(n7455), .B2(n6748), .Y(n9669) );
	nor2_1 U10171( .A(RST), .B(n6719), .Y(n4038) );
	o21ai_0 U10172( .A1(n6748), .A2(n15642), .B1(n9670), .Y(n6719) );
	a22oi_1 U10173( .A1(g1947), .A2(g7194), .B1(n9925), .B2(g7052), .Y(n9670) );
	nor2_1 U10174( .A(RST), .B(n6724), .Y(n4037) );
	o21ai_0 U10175( .A1(n6748), .A2(n15629), .B1(n9671), .Y(n6724) );
	a22oi_1 U10176( .A1(g1951), .A2(g7194), .B1(n9930), .B2(g7052), .Y(n9671) );
	inv_1 U10177( .A(n7225), .Y(n6748) );
	nor2_1 U10178( .A(RST), .B(n8963), .Y(n4036) );
	nand4_1 U10179( .A(n7703), .B(n6337), .C(n10081), .D(n9672), .Y(n8963) );
	nor4_1 U10180( .A(n10065), .B(n10066), .C(n7721), .D(n7303), .Y(n9672) );
	nor4_1 U10181( .A(n7247), .B(n7279), .C(n9673), .D(n7320), .Y(n6337) );
	or2_0 U10182( .A(n10084), .B(n7321), .X(n9673) );
	a211oi_1 U10183( .A1(g6944), .A2(n5421), .B1(n9674), .C1(RST), .Y(n4035) );
	o22ai_1 U10184( .A1(n9806), .A2(n7866), .B1(n7454), .B2(n7898), .Y(n9674) );
	a211oi_1 U10185( .A1(g6944), .A2(n5422), .B1(n9675), .C1(RST), .Y(n4034) );
	o22ai_1 U10186( .A1(n9804), .A2(n7866), .B1(n7461), .B2(n7898), .Y(n9675) );
	a211oi_1 U10187( .A1(g6944), .A2(n5423), .B1(n9676), .C1(RST), .Y(n4033) );
	o22ai_1 U10188( .A1(n9805), .A2(n7866), .B1(n7457), .B2(n7898), .Y(n9676) );
	nor2_1 U10189( .A(RST), .B(n7869), .Y(n4032) );
	o21ai_0 U10190( .A1(n7898), .A2(n15647), .B1(n9677), .Y(n7869) );
	a22oi_1 U10191( .A1(g1253), .A2(g6944), .B1(n9803), .B2(g6750), .Y(n9677) );
	nor2_1 U10192( .A(RST), .B(n7874), .Y(n4031) );
	o21ai_0 U10193( .A1(n7898), .A2(n15631), .B1(n9678), .Y(n7874) );
	a22oi_1 U10194( .A1(g1257), .A2(g6944), .B1(n9807), .B2(g6750), .Y(n9678) );
	inv_1 U10195( .A(n7226), .Y(n7898) );
	a211oi_1 U10196( .A1(g6642), .A2(n5424), .B1(n9679), .C1(RST), .Y(n4030) );
	o22ai_1 U10197( .A1(n9837), .A2(n8495), .B1(n7456), .B2(n8527), .Y(n9679) );
	a211oi_1 U10198( .A1(g6642), .A2(n5425), .B1(n9680), .C1(RST), .Y(n4029) );
	o22ai_1 U10199( .A1(n9835), .A2(n8495), .B1(n7462), .B2(n8527), .Y(n9680) );
	a211oi_1 U10200( .A1(g6642), .A2(n5426), .B1(n9681), .C1(RST), .Y(n4028) );
	o22ai_1 U10201( .A1(n9836), .A2(n8495), .B1(n7458), .B2(n8527), .Y(n9681) );
	nor2_1 U10202( .A(RST), .B(n8498), .Y(n4027) );
	o21ai_0 U10203( .A1(n8527), .A2(n15652), .B1(n9682), .Y(n8498) );
	a22oi_1 U10204( .A1(g567), .A2(g6642), .B1(n9834), .B2(g6485), .Y(n9682) );
	nor2_1 U10205( .A(RST), .B(n8503), .Y(n4026) );
	o21ai_0 U10206( .A1(n8527), .A2(n15638), .B1(n9683), .Y(n8503) );
	a22oi_1 U10207( .A1(g571), .A2(g6642), .B1(n9838), .B2(g6485), .Y(n9683) );
	inv_1 U10208( .A(n7227), .Y(n8527) );
	nor2_1 U10209( .A(RST), .B(n9684), .Y(n4025) );
	xor2_1 U10210( .A(n5855), .B(n9685), .X(n9684) );
	xor2_1 U10211( .A(n9686), .B(n9687), .X(n5855) );
	xor2_1 U10212( .A(n9688), .B(n9689), .X(n9687) );
	xnor2_1 U10213( .A(g8264), .B(g8263), .Y(n9689) );
	xnor2_1 U10214( .A(g8266), .B(g8265), .Y(n9688) );
	xor2_1 U10215( .A(n9690), .B(n9691), .X(n9686) );
	xor2_1 U10216( .A(g8262), .B(g8261), .X(n9691) );
	xnor2_1 U10217( .A(g8260), .B(g8259), .Y(n9690) );
	nor2_1 U10218( .A(RST), .B(n9692), .Y(n4024) );
	xor2_1 U10219( .A(n5857), .B(n9685), .X(n9692) );
	nor2_1 U10220( .A(n5414), .B(g3231), .Y(n9685) );
	xor2_1 U10221( .A(n9693), .B(n9694), .X(n5857) );
	xor2_1 U10222( .A(n9695), .B(n9696), .X(n9694) );
	xnor2_1 U10223( .A(g8273), .B(g8272), .Y(n9696) );
	xnor2_1 U10224( .A(g8275), .B(g8274), .Y(n9695) );
	xor2_1 U10225( .A(n9697), .B(n9698), .X(n9693) );
	xor2_1 U10226( .A(g8271), .B(g8270), .X(n9698) );
	xnor2_1 U10227( .A(g8269), .B(g8268), .Y(n9697) );
	and2_0 U10228( .A(g2363), .B(n5761), .X(n4023) );
	and2_0 U10229( .A(g2361), .B(n5754), .X(n4022) );
	and2_0 U10230( .A(g2359), .B(n5761), .X(n4021) );
	and2_0 U10231( .A(g2357), .B(n5761), .X(n4020) );
	and2_0 U10232( .A(g2355), .B(n5761), .X(n4019) );
	and2_0 U10233( .A(g2529), .B(n5761), .X(n4018) );
	and2_0 U10234( .A(g2527), .B(n5761), .X(n4017) );
	and2_0 U10235( .A(g2525), .B(n5761), .X(n4016) );
	and2_0 U10236( .A(g1669), .B(n5761), .X(n4015) );
	and2_0 U10237( .A(g1667), .B(n5761), .X(n4014) );
	and2_0 U10238( .A(g1665), .B(n5761), .X(n4013) );
	and2_0 U10239( .A(g1663), .B(n5761), .X(n4012) );
	and2_0 U10240( .A(g1661), .B(n5761), .X(n4011) );
	and2_0 U10241( .A(g1835), .B(n5761), .X(n4010) );
	and2_0 U10242( .A(g1833), .B(n5761), .X(n4009) );
	and2_0 U10243( .A(g1831), .B(n5760), .X(n4008) );
	and2_0 U10244( .A(g975), .B(n5760), .X(n4007) );
	and2_0 U10245( .A(g973), .B(n5760), .X(n4006) );
	and2_0 U10246( .A(g971), .B(n5760), .X(n4005) );
	and2_0 U10247( .A(g969), .B(n5760), .X(n4004) );
	and2_0 U10248( .A(g967), .B(n5760), .X(n4003) );
	and2_0 U10249( .A(g1141), .B(n5760), .X(n4002) );
	and2_0 U10250( .A(g1139), .B(n5760), .X(n4001) );
	and2_0 U10251( .A(g1137), .B(n5760), .X(n4000) );
	nor2_1 U10252( .A(RST), .B(n7250), .Y(n40) );
	nor2_1 U10253( .A(RST), .B(n7234), .Y(n4) );
	and2_0 U10254( .A(g288), .B(n5760), .X(n3999) );
	and2_0 U10255( .A(g286), .B(n5760), .X(n3998) );
	and2_0 U10256( .A(g284), .B(n5760), .X(n3997) );
	and2_0 U10257( .A(g282), .B(n5760), .X(n3996) );
	and2_0 U10258( .A(g280), .B(n5760), .X(n3995) );
	and2_0 U10259( .A(g454), .B(n5760), .X(n3994) );
	and2_0 U10260( .A(g452), .B(n5760), .X(n3993) );
	and2_0 U10261( .A(g450), .B(n5760), .X(n3992) );
	and2_0 U10262( .A(g2602), .B(n5760), .X(n3991) );
	and2_0 U10263( .A(g2587), .B(n5761), .X(n3990) );
	inv_1 U10264( .A(n9090), .Y(n3989) );
	nand2_1 U10265( .A(g2473), .B(n5749), .Y(n9090) );
	inv_1 U10266( .A(n9097), .Y(n3988) );
	nand2_1 U10267( .A(g2459), .B(n5749), .Y(n9097) );
	inv_1 U10268( .A(n9103), .Y(n3987) );
	nand2_1 U10269( .A(g2444), .B(n5749), .Y(n9103) );
	inv_1 U10270( .A(n9106), .Y(n3986) );
	nand2_1 U10271( .A(g2429), .B(n5749), .Y(n9106) );
	and2_0 U10272( .A(g1908), .B(n5763), .X(n3985) );
	and2_0 U10273( .A(g1893), .B(n5764), .X(n3984) );
	inv_1 U10274( .A(n9115), .Y(n3983) );
	nand2_1 U10275( .A(g1779), .B(n5749), .Y(n9115) );
	inv_1 U10276( .A(n9122), .Y(n3982) );
	nand2_1 U10277( .A(g1765), .B(n5749), .Y(n9122) );
	inv_1 U10278( .A(n9128), .Y(n3981) );
	nand2_1 U10279( .A(g1750), .B(n5749), .Y(n9128) );
	inv_1 U10280( .A(n9131), .Y(n3980) );
	nand2_1 U10281( .A(g1735), .B(n5749), .Y(n9131) );
	and2_0 U10282( .A(g1214), .B(n5765), .X(n3979) );
	and2_0 U10283( .A(g1199), .B(n5757), .X(n3978) );
	inv_1 U10284( .A(n9142), .Y(n3977) );
	nand2_1 U10285( .A(g1075), .B(n5750), .Y(n9142) );
	inv_1 U10286( .A(n9148), .Y(n3976) );
	nand2_1 U10287( .A(g1060), .B(n5750), .Y(n9148) );
	inv_1 U10288( .A(n9155), .Y(n3975) );
	nand2_1 U10289( .A(g1045), .B(n5750), .Y(n9155) );
	inv_1 U10290( .A(n9157), .Y(n3974) );
	nand2_1 U10291( .A(g1030), .B(n5750), .Y(n9157) );
	and2_0 U10292( .A(g2873), .B(n5756), .X(n3973) );
	and2_0 U10293( .A(g528), .B(n5755), .X(n3972) );
	and2_0 U10294( .A(g513), .B(n5745), .X(n3971) );
	inv_1 U10295( .A(n9170), .Y(n3970) );
	nand2_1 U10296( .A(g398), .B(n5750), .Y(n9170) );
	inv_1 U10297( .A(n9177), .Y(n3969) );
	nand2_1 U10298( .A(g384), .B(n5750), .Y(n9177) );
	inv_1 U10299( .A(n9183), .Y(n3968) );
	nand2_1 U10300( .A(g369), .B(n5750), .Y(n9183) );
	inv_1 U10301( .A(n9186), .Y(n3967) );
	nand2_1 U10302( .A(g354), .B(n5750), .Y(n9186) );
	and2_0 U10303( .A(g2857), .B(n5752), .X(n3966) );
	and2_0 U10304( .A(g2256), .B(n5748), .X(n3965) );
	and2_0 U10305( .A(g1562), .B(n5753), .X(n3964) );
	and2_0 U10306( .A(g868), .B(n5763), .X(n3963) );
	and2_0 U10307( .A(g180), .B(n5743), .X(n3962) );
	nor2_1 U10308( .A(n7932), .B(RST), .Y(n3961) );
	inv_1 U10309( .A(g6712), .Y(n7932) );
	nor2_1 U10310( .A(n6281), .B(RST), .Y(n3960) );
	inv_1 U10311( .A(g5555), .Y(n6281) );
	nor2_1 U10312( .A(n6939), .B(RST), .Y(n3959) );
	inv_1 U10313( .A(g5511), .Y(n6939) );
	nor2_1 U10314( .A(n8709), .B(RST), .Y(n3958) );
	inv_1 U10315( .A(g5437), .Y(n8709) );
	o21ai_0 U10316( .A1(n10032), .A2(n9005), .B1(n5820), .Y(n3957) );
	or2_0 U10317( .A(n7587), .B(RST), .X(n5820) );
	nand2_1 U10318( .A(g8021), .B(n5751), .Y(n9005) );
	nor2_1 U10319( .A(n7586), .B(RST), .Y(n39) );
	nor2_1 U10320( .A(n7242), .B(RST), .Y(n38) );
	nor2_1 U10321( .A(n6278), .B(RST), .Y(n37) );
	inv_1 U10322( .A(g7084), .Y(n6278) );
	nor2_1 U10323( .A(n6279), .B(RST), .Y(n36) );
	inv_1 U10324( .A(g6837), .Y(n6279) );
	inv_1 U10325( .A(n8988), .Y(n35) );
	nand2_1 U10326( .A(g499), .B(n5751), .Y(n8988) );
	nor2_1 U10327( .A(n8990), .B(RST), .Y(n34) );
	inv_1 U10328( .A(n9258), .Y(n8990) );
	mux2i_1 U10329( .A0(n9699), .A1(n14885), .S(g2574), .Y(n9258) );
	mux2i_1 U10330( .A0(n8993), .A1(n9913), .S(n6066), .Y(n9699) );
	inv_1 U10331( .A(g7302), .Y(n6066) );
	mux2i_1 U10332( .A0(n9700), .A1(n14880), .S(g1880), .Y(n8993) );
	mux2i_1 U10333( .A0(n9401), .A1(n9922), .S(n6716), .Y(n9700) );
	inv_1 U10334( .A(n6639), .Y(n33) );
	nand2_1 U10335( .A(n5755), .B(DFF_1153_D), .Y(n6639) );
	inv_1 U10336( .A(n8986), .Y(n32) );
	nand2_1 U10337( .A(g1880), .B(n5751), .Y(n8986) );
	nor2_1 U10338( .A(n8995), .B(RST), .Y(n31) );
	inv_1 U10339( .A(n9401), .Y(n8995) );
	mux2i_1 U10340( .A0(n9701), .A1(n14876), .S(g1186), .Y(n9401) );
	mux2i_1 U10341( .A0(n9702), .A1(n9923), .S(n7866), .Y(n9701) );
	inv_1 U10342( .A(n8998), .Y(n9702) );
	mux2i_1 U10343( .A0(n9703), .A1(g544), .S(g499), .Y(n8998) );
	nor2_1 U10344( .A(g6485), .B(n15417), .Y(n9703) );
	inv_1 U10345( .A(n9661), .Y(n3) );
	nand2_1 U10346( .A(g51), .B(n5751), .Y(n9661) );
	inv_1 U10347( .A(n6762), .Y(n29) );
	nand2_1 U10348( .A(g8082), .B(n5751), .Y(n6762) );
	inv_1 U10349( .A(n6765), .Y(n28) );
	nand2_1 U10350( .A(g8012), .B(n5751), .Y(n6765) );
	inv_1 U10351( .A(n9596), .Y(n27) );
	nand2_1 U10352( .A(g1852), .B(n5751), .Y(n9596) );
	inv_1 U10353( .A(n9597), .Y(n26) );
	nand2_1 U10354( .A(g1849), .B(n5751), .Y(n9597) );
	inv_1 U10355( .A(n9598), .Y(n25) );
	nand2_1 U10356( .A(g1846), .B(n5751), .Y(n9598) );
	inv_1 U10357( .A(n9599), .Y(n24) );
	nand2_1 U10358( .A(g1842), .B(n5751), .Y(n9599) );
	inv_1 U10359( .A(n9601), .Y(n23) );
	nand2_1 U10360( .A(g1839), .B(n5752), .Y(n9601) );
	inv_1 U10361( .A(n9602), .Y(n22) );
	nand2_1 U10362( .A(g1836), .B(n5752), .Y(n9602) );
	nor2_1 U10363( .A(n6721), .B(RST), .Y(n21) );
	inv_1 U10364( .A(g7194), .Y(n6721) );
	nor2_1 U10365( .A(n6716), .B(RST), .Y(n20) );
	inv_1 U10366( .A(g7052), .Y(n6716) );
	inv_1 U10367( .A(n9043), .Y(n19) );
	nand2_1 U10368( .A(g1772), .B(n5752), .Y(n9043) );
	inv_1 U10369( .A(n9046), .Y(n18) );
	nand2_1 U10370( .A(g1769), .B(n5752), .Y(n9046) );
	nor2_1 U10371( .A(n6774), .B(RST), .Y(n172) );
	inv_1 U10372( .A(g7014), .Y(n6774) );
	nor2_1 U10373( .A(RST), .B(n7268), .Y(n171) );
	nor2_1 U10374( .A(n6904), .B(RST), .Y(n170) );
	inv_1 U10375( .A(g6782), .Y(n6904) );
	inv_1 U10376( .A(n9048), .Y(n17) );
	nand2_1 U10377( .A(g1757), .B(n5752), .Y(n9048) );
	nor2_1 U10378( .A(n6905), .B(RST), .Y(n169) );
	inv_1 U10379( .A(g6573), .Y(n6905) );
	nor2_1 U10380( .A(RST), .B(n9628), .Y(n168) );
	inv_1 U10381( .A(g8096), .Y(n9628) );
	inv_1 U10382( .A(n7789), .Y(n167) );
	nand2_1 U10383( .A(n5755), .B(DFF_803_D), .Y(n7789) );
	nor2_1 U10384( .A(RST), .B(n9629), .Y(n166) );
	inv_1 U10385( .A(g4450), .Y(n9629) );
	nor2_1 U10386( .A(RST), .B(n9630), .Y(n165) );
	inv_1 U10387( .A(g4200), .Y(n9630) );
	nor2_1 U10388( .A(RST), .B(n9631), .Y(n164) );
	inv_1 U10389( .A(g3993), .Y(n9631) );
	nor2_1 U10390( .A(RST), .B(n9632), .Y(n163) );
	inv_1 U10391( .A(g8175), .Y(n9632) );
	inv_1 U10392( .A(n7910), .Y(n162) );
	nand2_1 U10393( .A(g8007), .B(n5752), .Y(n7910) );
	inv_1 U10394( .A(n7913), .Y(n161) );
	nand2_1 U10395( .A(g7961), .B(n5752), .Y(n7913) );
	inv_1 U10396( .A(n9606), .Y(n160) );
	nand2_1 U10397( .A(g1158), .B(n5752), .Y(n9606) );
	inv_1 U10398( .A(n9050), .Y(n16) );
	nand2_1 U10399( .A(g1754), .B(n5752), .Y(n9050) );
	inv_1 U10400( .A(n9608), .Y(n159) );
	nand2_1 U10401( .A(g1155), .B(n5752), .Y(n9608) );
	inv_1 U10402( .A(n9609), .Y(n158) );
	nand2_1 U10403( .A(g1152), .B(n5752), .Y(n9609) );
	nor2_1 U10404( .A(RST), .B(n9633), .Y(n157) );
	inv_1 U10405( .A(g8023), .Y(n9633) );
	inv_1 U10406( .A(n9610), .Y(n156) );
	nand2_1 U10407( .A(g1148), .B(n5752), .Y(n9610) );
	inv_1 U10408( .A(n9611), .Y(n155) );
	nand2_1 U10409( .A(g1145), .B(n5753), .Y(n9611) );
	inv_1 U10410( .A(n9612), .Y(n154) );
	nand2_1 U10411( .A(g1142), .B(n5753), .Y(n9612) );
	nor2_1 U10412( .A(n7871), .B(RST), .Y(n153) );
	inv_1 U10413( .A(g6944), .Y(n7871) );
	nor2_1 U10414( .A(n7866), .B(RST), .Y(n152) );
	inv_1 U10415( .A(g6750), .Y(n7866) );
	nor2_1 U10416( .A(RST), .B(n9634), .Y(n151) );
	inv_1 U10417( .A(g4321), .Y(n9634) );
	nor2_1 U10418( .A(RST), .B(n9635), .Y(n150) );
	inv_1 U10419( .A(g4088), .Y(n9635) );
	inv_1 U10420( .A(n9051), .Y(n15) );
	nand2_1 U10421( .A(g1742), .B(n5753), .Y(n9051) );
	nor2_1 U10422( .A(RST), .B(n9636), .Y(n149) );
	inv_1 U10423( .A(g8249), .Y(n9636) );
	nor2_1 U10424( .A(RST), .B(n9637), .Y(n148) );
	inv_1 U10425( .A(g7519), .Y(n9637) );
	nor2_1 U10426( .A(RST), .B(n9645), .Y(n147) );
	inv_1 U10427( .A(g7334), .Y(n9645) );
	inv_1 U10428( .A(n9058), .Y(n146) );
	nand2_1 U10429( .A(g1078), .B(n5753), .Y(n9058) );
	inv_1 U10430( .A(n9061), .Y(n145) );
	nand2_1 U10431( .A(g1085), .B(n5753), .Y(n9061) );
	inv_1 U10432( .A(n9063), .Y(n144) );
	nand2_1 U10433( .A(g1063), .B(n5753), .Y(n9063) );
	nor2_1 U10434( .A(n9164), .B(RST), .Y(n143) );
	inv_1 U10435( .A(g1071), .Y(n9164) );
	inv_1 U10436( .A(n9066), .Y(n142) );
	nand2_1 U10437( .A(g1048), .B(n5753), .Y(n9066) );
	nor2_1 U10438( .A(n9162), .B(RST), .Y(n141) );
	inv_1 U10439( .A(g1056), .Y(n9162) );
	inv_1 U10440( .A(n9069), .Y(n140) );
	nand2_1 U10441( .A(g1033), .B(n5753), .Y(n9069) );
	inv_1 U10442( .A(n9053), .Y(n14) );
	nand2_1 U10443( .A(g1739), .B(n5753), .Y(n9053) );
	nor2_1 U10444( .A(n9166), .B(RST), .Y(n139) );
	inv_1 U10445( .A(g1041), .Y(n9166) );
	nor2_1 U10446( .A(n8032), .B(RST), .Y(n138) );
	inv_1 U10447( .A(g5472), .Y(n8032) );
	nor2_1 U10448( .A(RST), .B(n9646), .Y(n137) );
	inv_1 U10449( .A(g6895), .Y(n9646) );
	nor2_1 U10450( .A(RST), .B(n9647), .Y(n136) );
	inv_1 U10451( .A(g6442), .Y(n9647) );
	nor2_1 U10452( .A(RST), .B(n9648), .Y(n135) );
	inv_1 U10453( .A(g6225), .Y(n9648) );
	nor2_1 U10454( .A(RST), .B(n9649), .Y(n134) );
	inv_1 U10455( .A(g4590), .Y(n9649) );
	nor2_1 U10456( .A(RST), .B(n7222), .Y(n133) );
	nor2_1 U10457( .A(RST), .B(n7240), .Y(n132) );
	nor2_1 U10458( .A(RST), .B(n7270), .Y(n131) );
	nor2_1 U10459( .A(RST), .B(n7245), .Y(n130) );
	inv_1 U10460( .A(n9054), .Y(n13) );
	nand2_1 U10461( .A(g1727), .B(n5753), .Y(n9054) );
	nor2_1 U10462( .A(RST), .B(n7248), .Y(n129) );
	nor2_1 U10463( .A(RST), .B(n7592), .Y(n128) );
	nor2_1 U10464( .A(RST), .B(n9650), .Y(n127) );
	inv_1 U10465( .A(g4323), .Y(n9650) );
	nor2_1 U10466( .A(n7251), .B(RST), .Y(n126) );
	nor2_1 U10467( .A(n7593), .B(RST), .Y(n125) );
	nor2_1 U10468( .A(n8049), .B(RST), .Y(n124) );
	inv_1 U10469( .A(g6518), .Y(n8049) );
	nor2_1 U10470( .A(n8050), .B(RST), .Y(n123) );
	inv_1 U10471( .A(g6368), .Y(n8050) );
	o22ai_1 U10472( .A1(n9032), .A2(n9035), .B1(RST), .B2(n9704), .Y(n122) );
	a21oi_1 U10473( .A1(n10081), .A2(n9705), .B1(n9034), .Y(n9704) );
	nand2_1 U10474( .A(n5361), .B(n9019), .Y(n9034) );
	nand2_1 U10475( .A(n9706), .B(n9707), .Y(n9019) );
	nor4_1 U10476( .A(n10081), .B(n10084), .C(n7320), .D(n9708), .Y(n9707) );
	and4_1 U10477( .A(n7247), .B(n7279), .C(n7321), .D(n7721), .X(n9706) );
	inv_1 U10478( .A(n4131), .Y(n9035) );
	nor2_1 U10479( .A(n9708), .B(RST), .Y(n4131) );
	inv_1 U10480( .A(g2950), .Y(n9708) );
	inv_1 U10481( .A(n9705), .Y(n9032) );
	nand2_1 U10482( .A(g2950), .B(n10081), .Y(n9705) );
	nor2_1 U10483( .A(RST), .B(n9651), .Y(n121) );
	inv_1 U10484( .A(g4090), .Y(n9651) );
	nor2_1 U10485( .A(RST), .B(n9652), .Y(n120) );
	inv_1 U10486( .A(g8251), .Y(n9652) );
	inv_1 U10487( .A(n9057), .Y(n12) );
	nand2_1 U10488( .A(g1724), .B(n5753), .Y(n9057) );
	inv_1 U10489( .A(n8418), .Y(n119) );
	nand2_1 U10490( .A(n5755), .B(DFF_453_D), .Y(n8418) );
	inv_1 U10491( .A(n8539), .Y(n118) );
	nand2_1 U10492( .A(g7956), .B(n5753), .Y(n8539) );
	inv_1 U10493( .A(n8542), .Y(n117) );
	nand2_1 U10494( .A(g7909), .B(n5754), .Y(n8542) );
	inv_1 U10495( .A(n9616), .Y(n116) );
	nand2_1 U10496( .A(g471), .B(n5754), .Y(n9616) );
	inv_1 U10497( .A(n9618), .Y(n115) );
	nand2_1 U10498( .A(g468), .B(n5754), .Y(n9618) );
	inv_1 U10499( .A(n9619), .Y(n114) );
	nand2_1 U10500( .A(g465), .B(n5754), .Y(n9619) );
	inv_1 U10501( .A(n9620), .Y(n113) );
	nand2_1 U10502( .A(g461), .B(n5754), .Y(n9620) );
	inv_1 U10503( .A(n9621), .Y(n112) );
	nand2_1 U10504( .A(g458), .B(n5754), .Y(n9621) );
	inv_1 U10505( .A(n9622), .Y(n111) );
	nand2_1 U10506( .A(g455), .B(n5754), .Y(n9622) );
	nor2_1 U10507( .A(n8500), .B(RST), .Y(n110) );
	inv_1 U10508( .A(g6642), .Y(n8500) );
	nor2_1 U10509( .A(RST), .B(n9653), .Y(n11) );
	inv_1 U10510( .A(g2877), .Y(n9653) );
	nor2_1 U10511( .A(n8495), .B(RST), .Y(n109) );
	inv_1 U10512( .A(g6485), .Y(n8495) );
	inv_1 U10513( .A(n9073), .Y(n108) );
	nand2_1 U10514( .A(g391), .B(n5754), .Y(n9073) );
	inv_1 U10515( .A(n9076), .Y(n107) );
	nand2_1 U10516( .A(g388), .B(n5754), .Y(n9076) );
	inv_1 U10517( .A(n9078), .Y(n106) );
	nand2_1 U10518( .A(g376), .B(n5754), .Y(n9078) );
	inv_1 U10519( .A(n9080), .Y(n105) );
	nand2_1 U10520( .A(g373), .B(n5754), .Y(n9080) );
	inv_1 U10521( .A(n9081), .Y(n104) );
	nand2_1 U10522( .A(g361), .B(n5754), .Y(n9081) );
	inv_1 U10523( .A(n9083), .Y(n103) );
	nand2_1 U10524( .A(g358), .B(n5754), .Y(n9083) );
	inv_1 U10525( .A(n9084), .Y(n102) );
	nand2_1 U10526( .A(g346), .B(n5755), .Y(n9084) );
	inv_1 U10527( .A(n9087), .Y(n101) );
	nand2_1 U10528( .A(g343), .B(n5741), .Y(n9087) );
	nor2_1 U10529( .A(n8692), .B(RST), .Y(n100) );
	inv_1 U10530( .A(g6447), .Y(n8692) );
	nor2_1 U10531( .A(n7243), .B(RST), .Y(n10) );
	inv_1 U10532( .A(n8979), .Y(g27380) );
	nor4_1 U10533( .A(n9709), .B(n9710), .C(n9711), .D(n9712), .Y(n8979) );
	o32ai_1 U10534( .A1(n9713), .A2(n7262), .A3(n9714), .B1(n9715), .B2(n5567), .Y(n9712) );
	a21oi_1 U10535( .A1(n9716), .A2(n9717), .B1(n9718), .Y(n9714) );
	mux2i_1 U10536( .A0(n7256), .A1(n9719), .S(n5352), .Y(n9716) );
	inv_1 U10537( .A(n9720), .Y(n9719) );
	a22oi_1 U10538( .A1(n9721), .A2(n7724), .B1(n9722), .B2(n7723), .Y(n9720) );
	nor2_1 U10539( .A(n9723), .B(n5382), .Y(n9711) );
	o22ai_1 U10540( .A1(n9883), .A2(n9724), .B1(n9725), .B2(n9726), .Y(n9710) );
	nand4_1 U10541( .A(n9727), .B(n9728), .C(n9729), .D(n9730), .Y(g26149) );
	a221oi_1 U10542( .A1(n9731), .A2(n9732), .B1(n9888), .B2(n9733), .C1(n9734), .Y(n9730) );
	o22ai_1 U10543( .A1(n9735), .A2(n5307), .B1(n9736), .B2(n5383), .Y(n9734) );
	inv_1 U10544( .A(n9715), .Y(n9733) );
	o22ai_1 U10545( .A1(n9737), .A2(n5308), .B1(n9738), .B2(n5384), .Y(n9732) );
	a221oi_1 U10546( .A1(n9890), .A2(n9739), .B1(n9981), .B2(n9740), .C1(n9741), .Y(n9729) );
	o22ai_1 U10547( .A1(n9742), .A2(n5309), .B1(n9743), .B2(n5385), .Y(n9741) );
	a221oi_1 U10548( .A1(n9891), .A2(n9744), .B1(n9906), .B2(n9745), .C1(n9746), .Y(n9728) );
	o22ai_1 U10549( .A1(n9747), .A2(n5310), .B1(n9748), .B2(n5386), .Y(n9746) );
	inv_1 U10550( .A(n9749), .Y(n9744) );
	a221oi_1 U10551( .A1(n9886), .A2(n9750), .B1(n9887), .B2(n9751), .C1(n9709), .Y(n9727) );
	inv_1 U10552( .A(n9752), .Y(n9709) );
	inv_1 U10553( .A(n9724), .Y(n9751) );
	nand4_1 U10554( .A(n9753), .B(n9754), .C(n9755), .D(n9756), .Y(g26135) );
	a221oi_1 U10555( .A1(n9924), .A2(n9757), .B1(n9927), .B2(n9758), .C1(n9759), .Y(n9756) );
	o22ai_1 U10556( .A1(n9715), .A2(n15162), .B1(n9760), .B2(n9725), .Y(n9759) );
	a222oi_1 U10557( .A1(n9718), .A2(n9722), .B1(n9983), .B2(n9761), .C1(n7666), .C2(n9717), .Y(n9760) );
	a221oi_1 U10558( .A1(n7722), .A2(n9762), .B1(n9982), .B2(n9739), .C1(n9763), .Y(n9755) );
	o22ai_1 U10559( .A1(n9742), .A2(n5311), .B1(n9743), .B2(n5387), .Y(n9763) );
	a221oi_1 U10560( .A1(n9916), .A2(n9745), .B1(n9912), .B2(n9764), .C1(n9765), .Y(n9754) );
	o22ai_1 U10561( .A1(n9749), .A2(n5312), .B1(n9766), .B2(n5388), .Y(n9765) );
	a221oi_1 U10562( .A1(n9915), .A2(n9767), .B1(n9750), .B2(n7723), .C1(n9768), .Y(n9753) );
	o21ai_0 U10563( .A1(g3128), .A2(n9724), .B1(n9752), .Y(n9768) );
	nand4_1 U10564( .A(n9769), .B(n9770), .C(n9771), .D(n9772), .Y(g26104) );
	a221oi_1 U10565( .A1(n9884), .A2(n9757), .B1(n9885), .B2(n9758), .C1(n9773), .Y(n9772) );
	o22ai_1 U10566( .A1(n9715), .A2(n5414), .B1(n9774), .B2(n9725), .Y(n9773) );
	inv_1 U10567( .A(n9731), .Y(n9725) );
	a222oi_1 U10568( .A1(n9718), .A2(n9721), .B1(n9985), .B2(n9761), .C1(n7640), .C2(n9717), .Y(n9774) );
	inv_1 U10569( .A(n9738), .Y(n9761) );
	nand3_1 U10570( .A(n9775), .B(n9776), .C(n9777), .Y(n9715) );
	inv_1 U10571( .A(n9735), .Y(n9758) );
	nand2_1 U10572( .A(n9778), .B(n9779), .Y(n9735) );
	inv_1 U10573( .A(n9736), .Y(n9757) );
	nand3_1 U10574( .A(n9713), .B(n5352), .C(n9780), .Y(n9736) );
	a221oi_1 U10575( .A1(n9979), .A2(n9762), .B1(n9984), .B2(n9739), .C1(n9781), .Y(n9771) );
	o22ai_1 U10576( .A1(n9742), .A2(n5313), .B1(n9743), .B2(n5500), .Y(n9781) );
	nand2_1 U10577( .A(n9779), .B(n9777), .Y(n9743) );
	nand2_1 U10578( .A(n9778), .B(n9780), .Y(n9742) );
	and3_1 U10579( .A(n7319), .B(n10054), .C(n9780), .X(n9739) );
	inv_1 U10580( .A(n9723), .Y(n9762) );
	nand3_1 U10581( .A(n9777), .B(n9775), .C(n7262), .Y(n9723) );
	a221oi_1 U10582( .A1(n9950), .A2(n9745), .B1(n9931), .B2(n9764), .C1(n9782), .Y(n9770) );
	o22ai_1 U10583( .A1(n9749), .A2(n5314), .B1(n9766), .B2(n5389), .Y(n9782) );
	inv_1 U10584( .A(n9740), .Y(n9766) );
	nor4_1 U10585( .A(n9776), .B(n9737), .C(n7319), .D(n10054), .Y(n9740) );
	nand3_1 U10586( .A(n7319), .B(n10054), .C(n9779), .Y(n9749) );
	nor2_1 U10587( .A(n9738), .B(n7262), .Y(n9779) );
	inv_1 U10588( .A(n9748), .Y(n9764) );
	nand2_1 U10589( .A(n9780), .B(n9777), .Y(n9748) );
	nor2_1 U10590( .A(n9738), .B(n9776), .Y(n9780) );
	nand2_1 U10591( .A(n9783), .B(n5483), .Y(n9738) );
	and3_1 U10592( .A(n9717), .B(n9776), .C(n9778), .X(n9745) );
	inv_1 U10593( .A(n7262), .Y(n9776) );
	a221oi_1 U10594( .A1(n9932), .A2(n9767), .B1(n9750), .B2(n7724), .C1(n9784), .Y(n9769) );
	o21ai_0 U10595( .A1(n9724), .A2(n15165), .B1(n9752), .Y(n9784) );
	inv_1 U10596( .A(n9785), .Y(n9750) );
	inv_1 U10597( .A(n9747), .Y(n9767) );
	nand3_1 U10598( .A(n7262), .B(n9717), .C(n9778), .Y(n9747) );
	nor2_1 U10599( .A(n5352), .B(n7319), .Y(n9778) );
	inv_1 U10600( .A(n9737), .Y(n9717) );
	nand2_1 U10601( .A(n10055), .B(n9783), .Y(n9737) );
	nor4_1 U10602( .A(n5739), .B(g3194), .C(g3198), .D(n10057), .Y(n9783) );
	mux2i_1 U10603( .A0(n9786), .A1(n9787), .S(n7722), .Y(g25489) );
	nand3_1 U10604( .A(n9983), .B(n9980), .C(n9979), .Y(n9787) );
	a21oi_1 U10605( .A1(n9722), .A2(n5382), .B1(n9788), .Y(n9786) );
	a21oi_1 U10606( .A1(n9789), .A2(n9980), .B1(n9979), .Y(n9788) );
	inv_1 U10607( .A(n9721), .Y(n9789) );
	nand2_1 U10608( .A(n15168), .B(n15169), .Y(n9721) );
	nand2_1 U10609( .A(n15172), .B(n15173), .Y(n9722) );
	o221ai_1 U10610( .A1(n9785), .A2(n15211), .B1(n9724), .B2(n15212), .C1( n9752), .Y(g25442) );
	o221ai_1 U10611( .A1(n9785), .A2(n15213), .B1(g3125), .B2(n9724), .C1(n9752), .Y(g25435) );
	o221ai_1 U10612( .A1(n9785), .A2(n15214), .B1(n9724), .B2(n15217), .C1( n9752), .Y(g25420) );
	nand2_1 U10613( .A(n9731), .B(n9775), .Y(n9785) );
	and2_0 U10614( .A(n9790), .B(n10055), .X(n9775) );
	nor3_1 U10615( .A(n7319), .B(n10054), .C(n7262), .Y(n9731) );
	o21ai_0 U10616( .A1(n10053), .A2(n9724), .B1(n9752), .Y(g24734) );
	nor2_1 U10617( .A(n9791), .B(g3230), .Y(n9752) );
	inv_1 U10618( .A(g3233), .Y(n9791) );
	nand3_1 U10619( .A(n7262), .B(n9777), .C(n9718), .Y(n9724) );
	inv_1 U10620( .A(n9726), .Y(n9718) );
	nand2_1 U10621( .A(n9790), .B(n5483), .Y(n9726) );
	nor4_1 U10622( .A(g3194), .B(g3198), .C(n10057), .D(n10056), .Y(n9790) );
	nor2_1 U10623( .A(n9713), .B(n10054), .Y(n9777) );
	inv_1 U10624( .A(n7319), .Y(n9713) );
	o21ai_0 U10625( .A1(n10033), .A2(n5858), .B1(n7255), .Y(g16496) );
	inv_1 U10626( .A(g5388), .Y(n5858) );
	xor2_1 troj6_0_U1( .A(tempn4402), .B(Trigger_en_6_0), .X(n4402) );
	inv_1 troj6_0_U2( .A(troj6_0_n1), .Y(Trigger_en_6_0) );
	or4_1 troj6_0_U3( .A(n5055), .B(n4530), .C(n4040), .D(troj6_0_n2), .X(troj6_0_n1) );
	or3_1 troj6_0_U4( .A(n7068), .B(n6976), .C(n5075), .X(troj6_0_n2) );
endmodule
