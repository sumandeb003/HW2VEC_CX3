
module c5315 (N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81,
N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631, N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128);

input N1, N4, N11, N14, N17, N20, N23, N24, N25, N26, N27, N31, N34, N37, N40, N43, N46, N49, N52, N53, N54, N61, N64, N67, N70, N73, N76, N79, N80, N81, N82, N83, N86, N87, N88, N91, N94, N97, N100, N103, N106, N109, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N140, N141, N145, N146, N149, N152, N155, N158, N161, N164, N167, N170, N173, N176, N179, N182, N185, N188, N191, N194, N197, N200, N203, N206, N209, N210, N217, N218, N225, N226, N233, N234, N241, N242, N245, N248, N251, N254, N257, N264, N265, N272, N273, N280, N281, N288, N289, N292, N293, N299, N302, N307, N308, N315, N316, N323, N324, N331, N332, N335, N338, N341, N348, N351, N358, N361, N366, N369, N372, N373, N374, N386, N389, N400, N411, N422, N435, N446, N457, N468, N479, N490, N503, N514, N523, N534, N545, N549, N552, N556, N559, N562, N566, N571, N574, N577, N580, N583, N588, N591, N592, N595, N596, N597, N598, N599, N603, N607, N610, N613, N616, N619, N625, N631;

output N709, N816, N1066, N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1147, N1152, N1153, N1154, N1155, N1972, N2054, N2060, N2061, N2139, N2142, N2309, N2387, N2527, N2584, N2590, N2623, N3357, N3358, N3359, N3360, N3604, N3613, N4272, N4275, N4278, N4279, N4737, N4738, N4739, N4740, N5240, N5388, N6641, N6643, N6646, N6648, N6716, N6877, N6924, N6925, N6926, N6927, N7015, N7363, N7365, N7432, N7449, N7465, N7466, N7467, N7469, N7470, N7471, N7472, N7473, N7474, N7476, N7503, N7504, N7506, N7511, N7515, N7516, N7517, N7518, N7519, N7520, N7521, N7522, N7600, N7601, N7602, N7603, N7604, N7605, N7606, N7607, N7626, N7698, N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7735, N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7754, N7755, N7756, N7757, N7758, N7759, N7760, N7761, N8075, N8076, N8123, N8124, N8127, N8128;

wire N1042, N1043, N1067, N1080, N1092, N1104, N1146, N1148, N1149, N1150, N1151, N1156, N1157, N1161, N1173, N1185, N1197, N1209, N1213, N1216, N1219, N1223, N1235, N1247, N1259, N1271, N1280, N1292, N1303, N1315, N1327, N1339, N1351, N1363, N1375, N1378, N1381, N1384, N1387, N1390, N1393, N1396, N1415, N1418, N1421, N1424, N1427, N1430, N1433, N1436, N1455, N1462, N1469, N1475, N1479, N1482, N1492, N1495, N1498, N1501, N1504, N1507, N1510, N1513, N1516, N1519, N1522, N1525, N1542, N1545, N1548, N1551, N1554, N1557, N1560, N1563, N1566, N1573, N1580, N1583, N1588, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, N1621, N1624, N1627, N1630, N1633, N1636, N1639, N1642, N1645, N1648, N1651, N1654, N1657, N1660, N1663, N1675, N1685, N1697, N1709, N1721, N1727, N1731, N1743, N1755, N1758, N1761, N1769, N1777, N1785, N1793, N1800, N1807, N1814, N1821, N1824, N1827, N1830, N1833, N1836, N1839, N1842, N1845, N1848, N1851, N1854, N1857, N1860, N1863, N1866, N1869, N1872, N1875, N1878, N1881, N1884, N1887, N1890, N1893, N1896, N1899, N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938, N1941, N1944, N1947, N1950, N1953, N1956, N1959, N1962, N1965, N1968, N2349, N2350, N2585, N2586, N2587, N2588, N2589, N2591, N2592, N2593, N2594, N2595, N2596, N2597, N2598, N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608, N2609, N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2617, N2618, N2619, N2620, N2621, N2622, N2624, N2625, N2626, N2627, N2628, N2629, N2630, N2631, N2632, N2633, N2634, N2635, N2636, N2637, N2638, N2639, N2640, N2641, N2642, N2643, N2644, N2645, N2646, N2647, N2653, N2664, N2675, N2681, N2692, N2703, N2704, N2709, N2710, N2711, N2712, N2713, N2714, N2715, N2716, N2717, N2718, N2719, N2720, N2721, N2722, N2728, N2739, N2750, N2756, N2767, N2778, N2779, N2790, N2801, N2812, N2823, N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2831, N2832, N2833, N2834, N2835, N2836, N2837, N2838, N2839, N2840, N2841, N2842, N2843, N2844, N2845, N2846, N2847, N2848, N2849, N2850, N2851, N2852, N2853, N2854, N2855, N2861, N2867, N2868, N2869, N2870, N2871, N2872, N2873, N2874, N2875, N2876, N2877, N2882, N2891, N2901, N2902, N2903, N2904, N2905, N2906, N2907, N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917, N2918, N2919, N2920, N2921, N2922, N2923, N2924, N2925, N2926, N2927, N2928, N2929, N2930, N2931, N2932, N2933, N2934, N2935, N2936, N2937, N2938, N2939, N2940, N2941, N2942, N2948, N2954, N2955, N2956, N2957, N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2969, N2970, N2971, N2972, N2973, N2974, N2975, N2976, N2977, N2978, N2979, N2980, N2981, N2982, N2983, N2984, N2985, N2986, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3003, N3006, N3007, N3010, N3013, N3014, N3015, N3016, N3017, N3018, N3019, N3020, N3021, N3022, N3023, N3024, N3025, N3026, N3027, N3028, N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3038, N3041, N3052, N3063, N3068, N3071, N3072, N3073, N3074, N3075, N3086, N3097, N3108, N3119, N3130, N3141, N3142, N3143, N3144, N3145, N3146, N3147, N3158, N3169, N3180, N3191, N3194, N3195, N3196, N3197, N3198, N3199, N3200, N3203, N3401, N3402, N3403, N3404, N3405, N3406, N3407, N3408, N3409, N3410, N3411, N3412, N3413, N3414, N3415, N3416, N3444, N3445, N3446, N3447, N3448, N3449, N3450, N3451, N3452, N3453, N3454, N3455, N3456, N3459, N3460, N3461, N3462, N3463, N3464, N3465, N3466, N3481, N3482, N3483, N3484, N3485, N3486, N3487, N3488, N3489, N3490, N3491, N3492, N3493, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509, N3510, N3511, N3512, N3513, N3514, N3515, N3558, N3559, N3560, N3561, N3562, N3563, N3605, N3606, N3607, N3608, N3609, N3610, N3614, N3615, N3616, N3617, N3618, N3619, N3620, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628, N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638, N3639, N3640, N3641, N3642, N3643, N3644, N3645, N3646, N3647, N3648, N3649, N3650, N3651, N3652, N3653, N3654, N3655, N3656, N3657, N3658, N3659, N3660, N3661, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3683, N3684, N3685, N3686, N3687, N3688, N3689, N3691, N3700, N3701, N3702, N3703, N3704, N3705, N3708, N3709, N3710, N3711, N3712, N3713, N3715, N3716, N3717, N3718, N3719, N3720, N3721, N3722, N3723, N3724, N3725, N3726, N3727, N3728, N3729, N3730, N3731, N3732, N3738, N3739, N3740, N3741, N3742, N3743, N3744, N3745, N3746, N3747, N3748, N3749, N3750, N3751, N3752, N3753, N3754, N3755, N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765, N3766, N3767, N3768, N3769, N3770, N3771, N3775, N3779, N3780, N3781, N3782, N3783, N3784, N3785, N3786, N3787, N3788, N3789, N3793, N3797, N3800, N3801, N3802, N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3810, N3813, N3816, N3819, N3822, N3823, N3824, N3827, N3828, N3829, N3830, N3831, N3834, N3835, N3836, N3837, N3838, N3839, N3840, N3841, N3842, N3849, N3855, N3861, N3867, N3873, N3881, N3887, N3893, N3908, N3909, N3911, N3914, N3915, N3916, N3917, N3918, N3919, N3920, N3921, N3927, N3933, N3942, N3948, N3956, N3962, N3968, N3975, N3976, N3977, N3978, N3979, N3980, N3981, N3982, N3983, N3984, N3987, N3988, N3989, N3990, N3991, N3998, N4008, N4011, N4021, N4024, N4027, N4031, N4032, N4033, N4034, N4035, N4036, N4037, N4038, N4039, N4040, N4041, N4042, N4067, N4080, N4088, N4091, N4094, N4097, N4100, N4103, N4106, N4109, N4144, N4147, N4150, N4153, N4156, N4159, N4183, N4184, N4185, N4186, N4188, N4191, N4196, N4197, N4198, N4199, N4200, N4203, N4206, N4209, N4212, N4215, N4219, N4223, N4224, N4225, N4228, N4231, N4234, N4237, N4240, N4243, N4246, N4249, N4252, N4255, N4258, N4263, N4264, N4267, N4268, N4269, N4270, N4271, N4273, N4274, N4276, N4277, N4280, N4284, N4290, N4297, N4298, N4301, N4305, N4310, N4316, N4320, N4325, N4331, N4332, N4336, N4342, N4349, N4357, N4364, N4375, N4379, N4385, N4392, N4396, N4400, N4405, N4412, N4418, N4425, N4436, N4440, N4445, N4451, N4456, N4462, N4469, N4477, N4512, N4515, N4516, N4521, N4523, N4524, N4532, N4547, N4548, N4551, N4554, N4557, N4560, N4563, N4566, N4569, N4572, N4575, N4578, N4581, N4584, N4587, N4590, N4593, N4596, N4599, N4602, N4605, N4608, N4611, N4614, N4617, N4621, N4624, N4627, N4630, N4633, N4637, N4640, N4643, N4646, N4649, N4652, N4655, N4658, N4662, N4665, N4668, N4671, N4674, N4677, N4680, N4683, N4686, N4689, N4692, N4695, N4698, N4701, N4702, N4720, N4721, N4724, N4725, N4726, N4727, N4728, N4729, N4730, N4731, N4732, N4733, N4734, N4735, N4736, N4741, N4855, N4856, N4908, N4909, N4939, N4942, N4947, N4953, N4954, N4955, N4956, N4957, N4958, N4959, N4960, N4961, N4965, N4966, N4967, N4968, N4972, N4973, N4974, N4975, N4976, N4977, N4978, N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N5049, N5052, N5053, N5054, N5055, N5056, N5057, N5058, N5059, N5060, N5061, N5062, N5063, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5074, N5075, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083, N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093, N5094, N5095, N5096, N5097, N5098, N5099, N5100, N5101, N5102, N5103, N5104, N5105, N5106, N5107, N5108, N5109, N5110, N5111, N5112, N5113, N5114, N5115, N5116, N5117, N5118, N5119, N5120, N5121, N5122, N5123, N5124, N5125, N5126, N5127, N5128, N5129, N5130, N5131, N5132, N5133, N5135, N5136, N5137, N5138, N5139, N5140, N5141, N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5150, N5153, N5154, N5155, N5156, N5157, N5160, N5161, N5162, N5163, N5164, N5165, N5166, N5169, N5172, N5173, N5176, N5177, N5180, N5183, N5186, N5189, N5192, N5195, N5198, N5199, N5202, N5205, N5208, N5211, N5214, N5217, N5220, N5223, N5224, N5225, N5226, N5227, N5228, N5229, N5230, N5232, N5233, N5234, N5235, N5236, N5239, N5241, N5242, N5243, N5244, N5245, N5246, N5247, N5248, N5249, N5250, N5252, N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262, N5263, N5264, N5274, N5275, N5282, N5283, N5284, N5298, N5299, N5300, N5303, N5304, N5305, N5306, N5307, N5308, N5309, N5310, N5311, N5312, N5315, N5319, N5324, N5328, N5331, N5332, N5346, N5363, N5364, N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5374, N5377, N5382, N5385, N5389, N5396, N5407, N5418, N5424, N5431, N5441, N5452, N5462, N5469, N5470, N5477, N5488, N5498, N5506, N5520, N5536, N5549, N5555, N5562, N5573, N5579, N5595, N5606, N5616, N5617, N5618, N5619, N5620, N5621, N5622, N5624, N5634, N5655, N5671, N5684, N5690, N5691, N5692, N5696, N5700, N5703, N5707, N5711, N5726, N5727, N5728, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5739, N5742, N5745, N5755, N5756, N5954, N5955, N5956, N6005, N6006, N6023, N6024, N6025, N6028, N6031, N6034, N6037, N6040, N6044, N6045, N6048, N6051, N6054, N6065, N6066, N6067, N6068, N6069, N6071, N6072, N6073, N6074, N6075, N6076, N6077, N6078, N6079, N6080, N6083, N6084, N6085, N6086, N6087, N6088, N6089, N6090, N6091, N6094, N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104, N6105, N6106, N6107, N6108, N6111, N6112, N6113, N6114, N6115, N6116, N6117, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128, N6129, N6130, N6131, N6132, N6133, N6134, N6135, N6136, N6137, N6138, N6139, N6140, N6143, N6144, N6145, N6146, N6147, N6148, N6149, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159, N6160, N6161, N6162, N6163, N6164, N6168, N6171, N6172, N6173, N6174, N6175, N6178, N6179, N6180, N6181, N6182, N6183, N6184, N6185, N6186, N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6197, N6200, N6203, N6206, N6209, N6212, N6215, N6218, N6221, N6234, N6235, N6238, N6241, N6244, N6247, N6250, N6253, N6256, N6259, N6262, N6265, N6268, N6271, N6274, N6277, N6280, N6283, N6286, N6289, N6292, N6295, N6298, N6301, N6304, N6307, N6310, N6313, N6316, N6319, N6322, N6325, N6328, N6331, N6335, N6338, N6341, N6344, N6347, N6350, N6353, N6356, N6359, N6364, N6367, N6370, N6373, N6374, N6375, N6376, N6377, N6378, N6382, N6386, N6388, N6392, N6397, N6411, N6415, N6419, N6427, N6434, N6437, N6441, N6445, N6448, N6449, N6466, N6469, N6470, N6471, N6472, N6473, N6474, N6475, N6476, N6477, N6478, N6482, N6486, N6490, N6494, N6500, N6504, N6508, N6512, N6516, N6526, N6536, N6539, N6553, N6556, N6566, N6569, N6572, N6575, N6580, N6584, N6587, N6592, N6599, N6606, N6609, N6619, N6622, N6630, N6631, N6632, N6633, N6634, N6637, N6640, N6650, N6651, N6653, N6655, N6657, N6659, N6660, N6661, N6662, N6663, N6664, N6666, N6668, N6670, N6672, N6675, N6680, N6681, N6682, N6683, N6689, N6690, N6691, N6692, N6693, N6695, N6698, N6699, N6700, N6703, N6708, N6709, N6710, N6711, N6712, N6713, N6714, N6715, N6718, N6719, N6720, N6721, N6722, N6724, N6739, N6740, N6741, N6744, N6745, N6746, N6751, N6752, N6753, N6754, N6755, N6760, N6761, N6762, N6772, N6773, N6776, N6777, N6782, N6783, N6784, N6785, N6790, N6791, N6792, N6795, N6801, N6802, N6803, N6804, N6805, N6806, N6807, N6808, N6809, N6810, N6811, N6812, N6813, N6814, N6815, N6816, N6817, N6823, N6824, N6825, N6826, N6827, N6828, N6829, N6830, N6831, N6834, N6835, N6836, N6837, N6838, N6839, N6840, N6841, N6842, N6843, N6844, N6850, N6851, N6852, N6853, N6854, N6855, N6856, N6857, N6860, N6861, N6862, N6863, N6866, N6872, N6873, N6874, N6875, N6876, N6879, N6880, N6881, N6884, N6885, N6888, N6889, N6890, N6891, N6894, N6895, N6896, N6897, N6900, N6901, N6904, N6905, N6908, N6909, N6912, N6913, N6914, N6915, N6916, N6919, N6922, N6923, N6930, N6932, N6935, N6936, N6937, N6938, N6939, N6940, N6946, N6947, N6948, N6949, N6953, N6954, N6955, N6956, N6957, N6958, N6964, N6965, N6966, N6967, N6973, N6974, N6975, N6976, N6977, N6978, N6979, N6987, N6990, N6999, N7002, N7003, N7006, N7011, N7012, N7013, N7016, N7018, N7019, N7020, N7021, N7022, N7023, N7028, N7031, N7034, N7037, N7040, N7041, N7044, N7045, N7046, N7047, N7048, N7049, N7054, N7057, N7060, N7064, N7065, N7072, N7073, N7074, N7075, N7076, N7079, N7080, N7083, N7084, N7085, N7086, N7087, N7088, N7089, N7090, N7093, N7094, N7097, N7101, N7105, N7110, N7114, N7115, N7116, N7125, N7126, N7127, N7130, N7131, N7139, N7140, N7141, N7146, N7147, N7149, N7150, N7151, N7152, N7153, N7158, N7159, N7160, N7166, N7167, N7168, N7169, N7170, N7171, N7172, N7173, N7174, N7175, N7176, N7177, N7178, N7179, N7180, N7181, N7182, N7183, N7184, N7185, N7186, N7187, N7188, N7189, N7190, N7196, N7197, N7198, N7204, N7205, N7206, N7207, N7208, N7209, N7212, N7215, N7216, N7217, N7218, N7219, N7222, N7225, N7228, N7229, N7236, N7239, N7242, N7245, N7250, N7257, N7260, N7263, N7268, N7269, N7270, N7276, N7282, N7288, N7294, N7300, N7301, N7304, N7310, N7320, N7321, N7328, N7338, N7339, N7340, N7341, N7342, N7349, N7357, N7364, N7394, N7397, N7402, N7405, N7406, N7407, N7408, N7409, N7412, N7415, N7416, N7417, N7418, N7419, N7420, N7421, N7424, N7425, N7426, N7427, N7428, N7429, N7430, N7431, N7433, N7434, N7435, N7436, N7437, N7438, N7439, N7440, N7441, N7442, N7443, N7444, N7445, N7446, N7447, N7448, N7450, N7451, N7452, N7453, N7454, N7455, N7456, N7457, N7458, N7459, N7460, N7461, N7462, N7463, N7464, N7468, N7479, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489, N7492, N7493, N7498, N7499, N7500, N7505, N7507, N7508, N7509, N7510, N7512, N7513, N7514, N7525, N7526, N7527, N7528, N7529, N7530, N7531, N7537, N7543, N7549, N7555, N7561, N7567, N7573, N7579, N7582, N7585, N7586, N7587, N7588, N7589, N7592, N7595, N7598, N7599, N7624, N7625, N7631, N7636, N7657, N7658, N7665, N7666, N7667, N7668, N7669, N7670, N7671, N7672, N7673, N7674, N7675, N7676, N7677, N7678, N7679, N7680, N7681, N7682, N7683, N7684, N7685, N7686, N7687, N7688, N7689, N7690, N7691, N7692, N7693, N7694, N7695, N7696, N7697, N7708, N7709, N7710, N7711, N7712, N7715, N7718, N7719, N7720, N7721, N7722, N7723, N7724, N7727, N7728, N7729, N7730, N7731, N7732, N7733, N7734, N7743, N7744, N7749, N7750, N7751, N7762, N7765, N7768, N7769, N7770, N7771, N7772, N7775, N7778, N7781, N7782, N7787, N7788, N7795, N7796, N7797, N7798, N7799, N7800, N7803, N7806, N7807, N7808, N7809, N7810, N7811, N7812, N7815, N7816, N7821, N7822, N7823, N7826, N7829, N7832, N7833, N7834, N7835, N7836, N7839, N7842, N7845, N7846, N7851, N7852, N7859, N7860, N7861, N7862, N7863, N7864, N7867, N7870, N7871, N7872, N7873, N7874, N7875, N7876, N7879, N7880, N7885, N7886, N7887, N7890, N7893, N7896, N7897, N7898, N7899, N7900, N7903, N7906, N7909, N7910, N7917, N7918, N7923, N7924, N7925, N7926, N7927, N7928, N7929, N7930, N7931, N7932, N7935, N7938, N7939, N7940, N7943, N7944, N7945, N7946, N7951, N7954, N7957, N7960, N7963, N7966, N7967, N7968, N7969, N7970, N7973, N7974, N7984, N7985, N7987, N7988, N7989, N7990, N7991, N7992, N7993, N7994, N7995, N7996, N7997, N7998, N8001, N8004, N8009, N8013, N8017, N8020, N8021, N8022, N8023, N8025, N8026, N8027, N8031, N8032, N8033, N8034, N8035, N8036, N8037, N8038, N8039, N8040, N8041, N8042, N8043, N8044, N8045, N8048, N8055, N8056, N8057, N8058, N8059, N8060, N8061, N8064, N8071, N8072, N8073, N8074, N8077, N8078, N8079, N8082, N8089, N8090, N8091, N8092, N8093, N8096, N8099, N8102, N8113, N8114, N8115, N8116, N8117, N8118, N8119, N8120, N8121, N8122, N8125, N8126;


wire Trigger_en52_0,  troj52_0n1,  troj52_0n2,  troj52_0n3,  troj52_0n4,  tempN7709;

nb1s1 U1 (.Q(N709), .DIN(N141));
nb1s1 U2 (.Q(N816), .DIN(N293));
and2s1 U3 (.Q(N1042), .DIN1(N135), .DIN2(N631));
hi1s1 U4 (.Q(N1043), .DIN(N591));
nb1s1 U5 (.Q(N1066), .DIN(N592));
hi1s1 U6 (.Q(N1067), .DIN(N595));
hi1s1 U7 (.Q(N1080), .DIN(N596));
hi1s1 U8 (.Q(N1092), .DIN(N597));
hi1s1 U9 (.Q(N1104), .DIN(N598));
hi1s1 U10 (.Q(N1137), .DIN(N545));
hi1s1 U11 (.Q(N1138), .DIN(N348));
hi1s1 U12 (.Q(N1139), .DIN(N366));
and2s1 U13 (.Q(N1140), .DIN1(N552), .DIN2(N562));
hi1s1 U14 (.Q(N1141), .DIN(N549));
hi1s1 U15 (.Q(N1142), .DIN(N545));
hi1s1 U16 (.Q(N1143), .DIN(N545));
hi1s1 U17 (.Q(N1144), .DIN(N338));
hi1s1 U18 (.Q(N1145), .DIN(N358));
nnd2s1 U19 (.Q(N1146), .DIN1(N373), .DIN2(N1));
and2s1 U20 (.Q(N1147), .DIN1(N141), .DIN2(N145));
hi1s1 U21 (.Q(N1148), .DIN(N592));
hi1s1 U22 (.Q(N1149), .DIN(N1042));
and2s1 U23 (.Q(N1150), .DIN1(N1043), .DIN2(N27));
and2s1 U24 (.Q(N1151), .DIN1(N386), .DIN2(N556));
hi1s1 U25 (.Q(N1152), .DIN(N245));
hi1s1 U26 (.Q(N1153), .DIN(N552));
hi1s1 U27 (.Q(N1154), .DIN(N562));
hi1s1 U28 (.Q(N1155), .DIN(N559));
and4s1 U29 (.Q(N1156), .DIN1(N386), .DIN2(N559), .DIN3(N556), .DIN4(N552));
hi1s1 U30 (.Q(N1157), .DIN(N566));
nb1s1 U31 (.Q(N1161), .DIN(N571));
nb1s1 U32 (.Q(N1173), .DIN(N574));
nb1s1 U33 (.Q(N1185), .DIN(N571));
nb1s1 U34 (.Q(N1197), .DIN(N574));
nb1s1 U35 (.Q(N1209), .DIN(N137));
nb1s1 U36 (.Q(N1213), .DIN(N137));
nb1s1 U37 (.Q(N1216), .DIN(N141));
hi1s1 U38 (.Q(N1219), .DIN(N583));
nb1s1 U39 (.Q(N1223), .DIN(N577));
nb1s1 U40 (.Q(N1235), .DIN(N580));
nb1s1 U41 (.Q(N1247), .DIN(N577));
nb1s1 U42 (.Q(N1259), .DIN(N580));
nb1s1 U43 (.Q(N1271), .DIN(N254));
nb1s1 U44 (.Q(N1280), .DIN(N251));
nb1s1 U45 (.Q(N1292), .DIN(N251));
nb1s1 U46 (.Q(N1303), .DIN(N248));
nb1s1 U47 (.Q(N1315), .DIN(N248));
nb1s1 U48 (.Q(N1327), .DIN(N610));
nb1s1 U49 (.Q(N1339), .DIN(N607));
nb1s1 U50 (.Q(N1351), .DIN(N613));
nb1s1 U51 (.Q(N1363), .DIN(N616));
nb1s1 U52 (.Q(N1375), .DIN(N210));
nb1s1 U53 (.Q(N1378), .DIN(N210));
nb1s1 U54 (.Q(N1381), .DIN(N218));
nb1s1 U55 (.Q(N1384), .DIN(N218));
nb1s1 U56 (.Q(N1387), .DIN(N226));
nb1s1 U57 (.Q(N1390), .DIN(N226));
nb1s1 U58 (.Q(N1393), .DIN(N234));
nb1s1 U59 (.Q(N1396), .DIN(N234));
nb1s1 U60 (.Q(N1415), .DIN(N257));
nb1s1 U61 (.Q(N1418), .DIN(N257));
nb1s1 U62 (.Q(N1421), .DIN(N265));
nb1s1 U63 (.Q(N1424), .DIN(N265));
nb1s1 U64 (.Q(N1427), .DIN(N273));
nb1s1 U65 (.Q(N1430), .DIN(N273));
nb1s1 U66 (.Q(N1433), .DIN(N281));
nb1s1 U67 (.Q(N1436), .DIN(N281));
nb1s1 U68 (.Q(N1455), .DIN(N335));
nb1s1 U69 (.Q(N1462), .DIN(N335));
nb1s1 U70 (.Q(N1469), .DIN(N206));
and2s1 U71 (.Q(N1475), .DIN1(N27), .DIN2(N31));
nb1s1 U72 (.Q(N1479), .DIN(N1));
nb1s1 U73 (.Q(N1482), .DIN(N588));
nb1s1 U74 (.Q(N1492), .DIN(N293));
nb1s1 U75 (.Q(N1495), .DIN(N302));
nb1s1 U76 (.Q(N1498), .DIN(N308));
nb1s1 U77 (.Q(N1501), .DIN(N308));
nb1s1 U78 (.Q(N1504), .DIN(N316));
nb1s1 U79 (.Q(N1507), .DIN(N316));
nb1s1 U80 (.Q(N1510), .DIN(N324));
nb1s1 U81 (.Q(N1513), .DIN(N324));
nb1s1 U82 (.Q(N1516), .DIN(N341));
nb1s1 U83 (.Q(N1519), .DIN(N341));
nb1s1 U84 (.Q(N1522), .DIN(N351));
nb1s1 U85 (.Q(N1525), .DIN(N351));
nb1s1 U86 (.Q(N1542), .DIN(N257));
nb1s1 U87 (.Q(N1545), .DIN(N257));
nb1s1 U88 (.Q(N1548), .DIN(N265));
nb1s1 U89 (.Q(N1551), .DIN(N265));
nb1s1 U90 (.Q(N1554), .DIN(N273));
nb1s1 U91 (.Q(N1557), .DIN(N273));
nb1s1 U92 (.Q(N1560), .DIN(N281));
nb1s1 U93 (.Q(N1563), .DIN(N281));
nb1s1 U94 (.Q(N1566), .DIN(N332));
nb1s1 U95 (.Q(N1573), .DIN(N332));
nb1s1 U96 (.Q(N1580), .DIN(N549));
and2s1 U97 (.Q(N1583), .DIN1(N31), .DIN2(N27));
hi1s1 U98 (.Q(N1588), .DIN(N588));
nb1s1 U99 (.Q(N1594), .DIN(N324));
nb1s1 U100 (.Q(N1597), .DIN(N324));
nb1s1 U101 (.Q(N1600), .DIN(N341));
nb1s1 U102 (.Q(N1603), .DIN(N341));
nb1s1 U103 (.Q(N1606), .DIN(N351));
nb1s1 U104 (.Q(N1609), .DIN(N351));
nb1s1 U105 (.Q(N1612), .DIN(N293));
nb1s1 U106 (.Q(N1615), .DIN(N302));
nb1s1 U107 (.Q(N1618), .DIN(N308));
nb1s1 U108 (.Q(N1621), .DIN(N308));
nb1s1 U109 (.Q(N1624), .DIN(N316));
nb1s1 U110 (.Q(N1627), .DIN(N316));
nb1s1 U111 (.Q(N1630), .DIN(N361));
nb1s1 U112 (.Q(N1633), .DIN(N361));
nb1s1 U113 (.Q(N1636), .DIN(N210));
nb1s1 U114 (.Q(N1639), .DIN(N210));
nb1s1 U115 (.Q(N1642), .DIN(N218));
nb1s1 U116 (.Q(N1645), .DIN(N218));
nb1s1 U117 (.Q(N1648), .DIN(N226));
nb1s1 U118 (.Q(N1651), .DIN(N226));
nb1s1 U119 (.Q(N1654), .DIN(N234));
nb1s1 U120 (.Q(N1657), .DIN(N234));
hi1s1 U121 (.Q(N1660), .DIN(N324));
nb1s1 U122 (.Q(N1663), .DIN(N242));
nb1s1 U123 (.Q(N1675), .DIN(N242));
nb1s1 U124 (.Q(N1685), .DIN(N254));
nb1s1 U125 (.Q(N1697), .DIN(N610));
nb1s1 U126 (.Q(N1709), .DIN(N607));
nb1s1 U127 (.Q(N1721), .DIN(N625));
nb1s1 U128 (.Q(N1727), .DIN(N619));
nb1s1 U129 (.Q(N1731), .DIN(N613));
nb1s1 U130 (.Q(N1743), .DIN(N616));
hi1s1 U131 (.Q(N1755), .DIN(N599));
hi1s1 U132 (.Q(N1758), .DIN(N603));
nb1s1 U133 (.Q(N1761), .DIN(N619));
nb1s1 U134 (.Q(N1769), .DIN(N625));
nb1s1 U135 (.Q(N1777), .DIN(N619));
nb1s1 U136 (.Q(N1785), .DIN(N625));
nb1s1 U137 (.Q(N1793), .DIN(N619));
nb1s1 U138 (.Q(N1800), .DIN(N625));
nb1s1 U139 (.Q(N1807), .DIN(N619));
nb1s1 U140 (.Q(N1814), .DIN(N625));
nb1s1 U141 (.Q(N1821), .DIN(N299));
nb1s1 U142 (.Q(N1824), .DIN(N446));
nb1s1 U143 (.Q(N1827), .DIN(N457));
nb1s1 U144 (.Q(N1830), .DIN(N468));
nb1s1 U145 (.Q(N1833), .DIN(N422));
nb1s1 U146 (.Q(N1836), .DIN(N435));
nb1s1 U147 (.Q(N1839), .DIN(N389));
nb1s1 U148 (.Q(N1842), .DIN(N400));
nb1s1 U149 (.Q(N1845), .DIN(N411));
nb1s1 U150 (.Q(N1848), .DIN(N374));
nb1s1 U151 (.Q(N1851), .DIN(N4));
nb1s1 U152 (.Q(N1854), .DIN(N446));
nb1s1 U153 (.Q(N1857), .DIN(N457));
nb1s1 U154 (.Q(N1860), .DIN(N468));
nb1s1 U155 (.Q(N1863), .DIN(N435));
nb1s1 U156 (.Q(N1866), .DIN(N389));
nb1s1 U157 (.Q(N1869), .DIN(N400));
nb1s1 U158 (.Q(N1872), .DIN(N411));
nb1s1 U159 (.Q(N1875), .DIN(N422));
nb1s1 U160 (.Q(N1878), .DIN(N374));
nb1s1 U161 (.Q(N1881), .DIN(N479));
nb1s1 U162 (.Q(N1884), .DIN(N490));
nb1s1 U163 (.Q(N1887), .DIN(N503));
nb1s1 U164 (.Q(N1890), .DIN(N514));
nb1s1 U165 (.Q(N1893), .DIN(N523));
nb1s1 U166 (.Q(N1896), .DIN(N534));
nb1s1 U167 (.Q(N1899), .DIN(N54));
nb1s1 U168 (.Q(N1902), .DIN(N479));
nb1s1 U169 (.Q(N1905), .DIN(N503));
nb1s1 U170 (.Q(N1908), .DIN(N514));
nb1s1 U171 (.Q(N1911), .DIN(N523));
nb1s1 U172 (.Q(N1914), .DIN(N534));
nb1s1 U173 (.Q(N1917), .DIN(N490));
nb1s1 U174 (.Q(N1920), .DIN(N361));
nb1s1 U175 (.Q(N1923), .DIN(N369));
nb1s1 U176 (.Q(N1926), .DIN(N341));
nb1s1 U177 (.Q(N1929), .DIN(N351));
nb1s1 U178 (.Q(N1932), .DIN(N308));
nb1s1 U179 (.Q(N1935), .DIN(N316));
nb1s1 U180 (.Q(N1938), .DIN(N293));
nb1s1 U181 (.Q(N1941), .DIN(N302));
nb1s1 U182 (.Q(N1944), .DIN(N281));
nb1s1 U183 (.Q(N1947), .DIN(N289));
nb1s1 U184 (.Q(N1950), .DIN(N265));
nb1s1 U185 (.Q(N1953), .DIN(N273));
nb1s1 U186 (.Q(N1956), .DIN(N234));
nb1s1 U187 (.Q(N1959), .DIN(N257));
nb1s1 U188 (.Q(N1962), .DIN(N218));
nb1s1 U189 (.Q(N1965), .DIN(N226));
nb1s1 U190 (.Q(N1968), .DIN(N210));
hi1s1 U191 (.Q(N1972), .DIN(N1146));
and2s1 U192 (.Q(N2054), .DIN1(N136), .DIN2(N1148));
hi1s1 U193 (.Q(N2060), .DIN(N1150));
hi1s1 U194 (.Q(N2061), .DIN(N1151));
nb1s1 U195 (.Q(N2139), .DIN(N1209));
nb1s1 U196 (.Q(N2142), .DIN(N1216));
nb1s1 U197 (.Q(N2309), .DIN(N1479));
and2s1 U198 (.Q(N2349), .DIN1(N1104), .DIN2(N514));
or2s1 U199 (.Q(N2350), .DIN1(N1067), .DIN2(N514));
nb1s1 U200 (.Q(N2387), .DIN(N1580));
nb1s1 U201 (.Q(N2527), .DIN(N1821));
hi1s1 U202 (.Q(N2584), .DIN(N1580));
and3s1 U203 (.Q(N2585), .DIN1(N170), .DIN2(N1161), .DIN3(N1173));
and3s1 U204 (.Q(N2586), .DIN1(N173), .DIN2(N1161), .DIN3(N1173));
and3s1 U205 (.Q(N2587), .DIN1(N167), .DIN2(N1161), .DIN3(N1173));
and3s1 U206 (.Q(N2588), .DIN1(N164), .DIN2(N1161), .DIN3(N1173));
and3s1 U207 (.Q(N2589), .DIN1(N161), .DIN2(N1161), .DIN3(N1173));
nnd2s1 U208 (.Q(N2590), .DIN1(N1475), .DIN2(N140));
and3s1 U209 (.Q(N2591), .DIN1(N185), .DIN2(N1185), .DIN3(N1197));
and3s1 U210 (.Q(N2592), .DIN1(N158), .DIN2(N1185), .DIN3(N1197));
and3s1 U211 (.Q(N2593), .DIN1(N152), .DIN2(N1185), .DIN3(N1197));
and3s1 U212 (.Q(N2594), .DIN1(N146), .DIN2(N1185), .DIN3(N1197));
and3s1 U213 (.Q(N2595), .DIN1(N170), .DIN2(N1223), .DIN3(N1235));
and3s1 U214 (.Q(N2596), .DIN1(N173), .DIN2(N1223), .DIN3(N1235));
and3s1 U215 (.Q(N2597), .DIN1(N167), .DIN2(N1223), .DIN3(N1235));
and3s1 U216 (.Q(N2598), .DIN1(N164), .DIN2(N1223), .DIN3(N1235));
and3s1 U217 (.Q(N2599), .DIN1(N161), .DIN2(N1223), .DIN3(N1235));
and3s1 U218 (.Q(N2600), .DIN1(N185), .DIN2(N1247), .DIN3(N1259));
and3s1 U219 (.Q(N2601), .DIN1(N158), .DIN2(N1247), .DIN3(N1259));
and3s1 U220 (.Q(N2602), .DIN1(N152), .DIN2(N1247), .DIN3(N1259));
and3s1 U221 (.Q(N2603), .DIN1(N146), .DIN2(N1247), .DIN3(N1259));
and3s1 U222 (.Q(N2604), .DIN1(N106), .DIN2(N1731), .DIN3(N1743));
and3s1 U223 (.Q(N2605), .DIN1(N61), .DIN2(N1327), .DIN3(N1339));
and3s1 U224 (.Q(N2606), .DIN1(N106), .DIN2(N1697), .DIN3(N1709));
and3s1 U225 (.Q(N2607), .DIN1(N49), .DIN2(N1697), .DIN3(N1709));
and3s1 U226 (.Q(N2608), .DIN1(N103), .DIN2(N1697), .DIN3(N1709));
and3s1 U227 (.Q(N2609), .DIN1(N40), .DIN2(N1697), .DIN3(N1709));
and3s1 U228 (.Q(N2610), .DIN1(N37), .DIN2(N1697), .DIN3(N1709));
and3s1 U229 (.Q(N2611), .DIN1(N20), .DIN2(N1327), .DIN3(N1339));
and3s1 U230 (.Q(N2612), .DIN1(N17), .DIN2(N1327), .DIN3(N1339));
and3s1 U231 (.Q(N2613), .DIN1(N70), .DIN2(N1327), .DIN3(N1339));
and3s1 U232 (.Q(N2614), .DIN1(N64), .DIN2(N1327), .DIN3(N1339));
and3s1 U233 (.Q(N2615), .DIN1(N49), .DIN2(N1731), .DIN3(N1743));
and3s1 U234 (.Q(N2616), .DIN1(N103), .DIN2(N1731), .DIN3(N1743));
and3s1 U235 (.Q(N2617), .DIN1(N40), .DIN2(N1731), .DIN3(N1743));
and3s1 U236 (.Q(N2618), .DIN1(N37), .DIN2(N1731), .DIN3(N1743));
and3s1 U237 (.Q(N2619), .DIN1(N20), .DIN2(N1351), .DIN3(N1363));
and3s1 U238 (.Q(N2620), .DIN1(N17), .DIN2(N1351), .DIN3(N1363));
and3s1 U239 (.Q(N2621), .DIN1(N70), .DIN2(N1351), .DIN3(N1363));
and3s1 U240 (.Q(N2622), .DIN1(N64), .DIN2(N1351), .DIN3(N1363));
hi1s1 U241 (.Q(N2623), .DIN(N1475));
and3s1 U242 (.Q(N2624), .DIN1(N123), .DIN2(N1758), .DIN3(N599));
and2s1 U243 (.Q(N2625), .DIN1(N1777), .DIN2(N1785));
and3s1 U244 (.Q(N2626), .DIN1(N61), .DIN2(N1351), .DIN3(N1363));
and2s1 U245 (.Q(N2627), .DIN1(N1761), .DIN2(N1769));
hi1s1 U246 (.Q(N2628), .DIN(N1824));
hi1s1 U247 (.Q(N2629), .DIN(N1827));
hi1s1 U248 (.Q(N2630), .DIN(N1830));
hi1s1 U249 (.Q(N2631), .DIN(N1833));
hi1s1 U250 (.Q(N2632), .DIN(N1836));
hi1s1 U251 (.Q(N2633), .DIN(N1839));
hi1s1 U252 (.Q(N2634), .DIN(N1842));
hi1s1 U253 (.Q(N2635), .DIN(N1845));
hi1s1 U254 (.Q(N2636), .DIN(N1848));
hi1s1 U255 (.Q(N2637), .DIN(N1851));
hi1s1 U256 (.Q(N2638), .DIN(N1854));
hi1s1 U257 (.Q(N2639), .DIN(N1857));
hi1s1 U258 (.Q(N2640), .DIN(N1860));
hi1s1 U259 (.Q(N2641), .DIN(N1863));
hi1s1 U260 (.Q(N2642), .DIN(N1866));
hi1s1 U261 (.Q(N2643), .DIN(N1869));
hi1s1 U262 (.Q(N2644), .DIN(N1872));
hi1s1 U263 (.Q(N2645), .DIN(N1875));
hi1s1 U264 (.Q(N2646), .DIN(N1878));
nb1s1 U265 (.Q(N2647), .DIN(N1209));
hi1s1 U266 (.Q(N2653), .DIN(N1161));
hi1s1 U267 (.Q(N2664), .DIN(N1173));
nb1s1 U268 (.Q(N2675), .DIN(N1209));
hi1s1 U269 (.Q(N2681), .DIN(N1185));
hi1s1 U270 (.Q(N2692), .DIN(N1197));
and3s1 U271 (.Q(N2703), .DIN1(N179), .DIN2(N1185), .DIN3(N1197));
nb1s1 U272 (.Q(N2704), .DIN(N1479));
hi1s1 U273 (.Q(N2709), .DIN(N1881));
hi1s1 U274 (.Q(N2710), .DIN(N1884));
hi1s1 U275 (.Q(N2711), .DIN(N1887));
hi1s1 U276 (.Q(N2712), .DIN(N1890));
hi1s1 U277 (.Q(N2713), .DIN(N1893));
hi1s1 U278 (.Q(N2714), .DIN(N1896));
hi1s1 U279 (.Q(N2715), .DIN(N1899));
hi1s1 U280 (.Q(N2716), .DIN(N1902));
hi1s1 U281 (.Q(N2717), .DIN(N1905));
hi1s1 U282 (.Q(N2718), .DIN(N1908));
hi1s1 U283 (.Q(N2719), .DIN(N1911));
hi1s1 U284 (.Q(N2720), .DIN(N1914));
hi1s1 U285 (.Q(N2721), .DIN(N1917));
nb1s1 U286 (.Q(N2722), .DIN(N1213));
hi1s1 U287 (.Q(N2728), .DIN(N1223));
hi1s1 U288 (.Q(N2739), .DIN(N1235));
nb1s1 U289 (.Q(N2750), .DIN(N1213));
hi1s1 U290 (.Q(N2756), .DIN(N1247));
hi1s1 U291 (.Q(N2767), .DIN(N1259));
and3s1 U292 (.Q(N2778), .DIN1(N179), .DIN2(N1247), .DIN3(N1259));
hi1s1 U293 (.Q(N2779), .DIN(N1327));
hi1s1 U294 (.Q(N2790), .DIN(N1339));
hi1s1 U295 (.Q(N2801), .DIN(N1351));
hi1s1 U296 (.Q(N2812), .DIN(N1363));
hi1s1 U297 (.Q(N2823), .DIN(N1375));
hi1s1 U298 (.Q(N2824), .DIN(N1378));
hi1s1 U299 (.Q(N2825), .DIN(N1381));
hi1s1 U300 (.Q(N2826), .DIN(N1384));
hi1s1 U301 (.Q(N2827), .DIN(N1387));
hi1s1 U302 (.Q(N2828), .DIN(N1390));
hi1s1 U303 (.Q(N2829), .DIN(N1393));
hi1s1 U304 (.Q(N2830), .DIN(N1396));
and3s1 U305 (.Q(N2831), .DIN1(N1104), .DIN2(N457), .DIN3(N1378));
and3s1 U306 (.Q(N2832), .DIN1(N1104), .DIN2(N468), .DIN3(N1384));
and3s1 U307 (.Q(N2833), .DIN1(N1104), .DIN2(N422), .DIN3(N1390));
and3s1 U308 (.Q(N2834), .DIN1(N1104), .DIN2(N435), .DIN3(N1396));
and2s1 U309 (.Q(N2835), .DIN1(N1067), .DIN2(N1375));
and2s1 U310 (.Q(N2836), .DIN1(N1067), .DIN2(N1381));
and2s1 U311 (.Q(N2837), .DIN1(N1067), .DIN2(N1387));
and2s1 U312 (.Q(N2838), .DIN1(N1067), .DIN2(N1393));
hi1s1 U313 (.Q(N2839), .DIN(N1415));
hi1s1 U314 (.Q(N2840), .DIN(N1418));
hi1s1 U315 (.Q(N2841), .DIN(N1421));
hi1s1 U316 (.Q(N2842), .DIN(N1424));
hi1s1 U317 (.Q(N2843), .DIN(N1427));
hi1s1 U318 (.Q(N2844), .DIN(N1430));
hi1s1 U319 (.Q(N2845), .DIN(N1433));
hi1s1 U320 (.Q(N2846), .DIN(N1436));
and3s1 U321 (.Q(N2847), .DIN1(N1104), .DIN2(N389), .DIN3(N1418));
and3s1 U322 (.Q(N2848), .DIN1(N1104), .DIN2(N400), .DIN3(N1424));
and3s1 U323 (.Q(N2849), .DIN1(N1104), .DIN2(N411), .DIN3(N1430));
and3s1 U324 (.Q(N2850), .DIN1(N1104), .DIN2(N374), .DIN3(N1436));
and2s1 U325 (.Q(N2851), .DIN1(N1067), .DIN2(N1415));
and2s1 U326 (.Q(N2852), .DIN1(N1067), .DIN2(N1421));
and2s1 U327 (.Q(N2853), .DIN1(N1067), .DIN2(N1427));
and2s1 U328 (.Q(N2854), .DIN1(N1067), .DIN2(N1433));
hi1s1 U329 (.Q(N2855), .DIN(N1455));
hi1s1 U330 (.Q(N2861), .DIN(N1462));
and2s1 U331 (.Q(N2867), .DIN1(N292), .DIN2(N1455));
and2s1 U332 (.Q(N2868), .DIN1(N288), .DIN2(N1455));
and2s1 U333 (.Q(N2869), .DIN1(N280), .DIN2(N1455));
and2s1 U334 (.Q(N2870), .DIN1(N272), .DIN2(N1455));
and2s1 U335 (.Q(N2871), .DIN1(N264), .DIN2(N1455));
and2s1 U336 (.Q(N2872), .DIN1(N241), .DIN2(N1462));
and2s1 U337 (.Q(N2873), .DIN1(N233), .DIN2(N1462));
and2s1 U338 (.Q(N2874), .DIN1(N225), .DIN2(N1462));
and2s1 U339 (.Q(N2875), .DIN1(N217), .DIN2(N1462));
and2s1 U340 (.Q(N2876), .DIN1(N209), .DIN2(N1462));
nb1s1 U341 (.Q(N2877), .DIN(N1216));
hi1s1 U342 (.Q(N2882), .DIN(N1482));
hi1s1 U343 (.Q(N2891), .DIN(N1475));
hi1s1 U344 (.Q(N2901), .DIN(N1492));
hi1s1 U345 (.Q(N2902), .DIN(N1495));
hi1s1 U346 (.Q(N2903), .DIN(N1498));
hi1s1 U347 (.Q(N2904), .DIN(N1501));
hi1s1 U348 (.Q(N2905), .DIN(N1504));
hi1s1 U349 (.Q(N2906), .DIN(N1507));
and2s1 U350 (.Q(N2907), .DIN1(N1303), .DIN2(N1495));
and3s1 U351 (.Q(N2908), .DIN1(N1303), .DIN2(N479), .DIN3(N1501));
and3s1 U352 (.Q(N2909), .DIN1(N1303), .DIN2(N490), .DIN3(N1507));
and2s1 U353 (.Q(N2910), .DIN1(N1663), .DIN2(N1492));
and2s1 U354 (.Q(N2911), .DIN1(N1663), .DIN2(N1498));
and2s1 U355 (.Q(N2912), .DIN1(N1663), .DIN2(N1504));
hi1s1 U356 (.Q(N2913), .DIN(N1510));
hi1s1 U357 (.Q(N2914), .DIN(N1513));
hi1s1 U358 (.Q(N2915), .DIN(N1516));
hi1s1 U359 (.Q(N2916), .DIN(N1519));
hi1s1 U360 (.Q(N2917), .DIN(N1522));
hi1s1 U361 (.Q(N2918), .DIN(N1525));
and3s1 U362 (.Q(N2919), .DIN1(N1104), .DIN2(N503), .DIN3(N1513));
hi1s1 U363 (.Q(N2920), .DIN(N2349));
and3s1 U364 (.Q(N2921), .DIN1(N1104), .DIN2(N523), .DIN3(N1519));
and3s1 U365 (.Q(N2922), .DIN1(N1104), .DIN2(N534), .DIN3(N1525));
and2s1 U366 (.Q(N2923), .DIN1(N1067), .DIN2(N1510));
and2s1 U367 (.Q(N2924), .DIN1(N1067), .DIN2(N1516));
and2s1 U368 (.Q(N2925), .DIN1(N1067), .DIN2(N1522));
hi1s1 U369 (.Q(N2926), .DIN(N1542));
hi1s1 U370 (.Q(N2927), .DIN(N1545));
hi1s1 U371 (.Q(N2928), .DIN(N1548));
hi1s1 U372 (.Q(N2929), .DIN(N1551));
hi1s1 U373 (.Q(N2930), .DIN(N1554));
hi1s1 U374 (.Q(N2931), .DIN(N1557));
hi1s1 U375 (.Q(N2932), .DIN(N1560));
hi1s1 U376 (.Q(N2933), .DIN(N1563));
and3s1 U377 (.Q(N2934), .DIN1(N1303), .DIN2(N389), .DIN3(N1545));
and3s1 U378 (.Q(N2935), .DIN1(N1303), .DIN2(N400), .DIN3(N1551));
and3s1 U379 (.Q(N2936), .DIN1(N1303), .DIN2(N411), .DIN3(N1557));
and3s1 U380 (.Q(N2937), .DIN1(N1303), .DIN2(N374), .DIN3(N1563));
and2s1 U381 (.Q(N2938), .DIN1(N1663), .DIN2(N1542));
and2s1 U382 (.Q(N2939), .DIN1(N1663), .DIN2(N1548));
and2s1 U383 (.Q(N2940), .DIN1(N1663), .DIN2(N1554));
and2s1 U384 (.Q(N2941), .DIN1(N1663), .DIN2(N1560));
hi1s1 U385 (.Q(N2942), .DIN(N1566));
hi1s1 U386 (.Q(N2948), .DIN(N1573));
and2s1 U387 (.Q(N2954), .DIN1(N372), .DIN2(N1566));
and2s1 U388 (.Q(N2955), .DIN1(N366), .DIN2(N1566));
and2s1 U389 (.Q(N2956), .DIN1(N358), .DIN2(N1566));
and2s1 U390 (.Q(N2957), .DIN1(N348), .DIN2(N1566));
and2s1 U391 (.Q(N2958), .DIN1(N338), .DIN2(N1566));
and2s1 U392 (.Q(N2959), .DIN1(N331), .DIN2(N1573));
and2s1 U393 (.Q(N2960), .DIN1(N323), .DIN2(N1573));
and2s1 U394 (.Q(N2961), .DIN1(N315), .DIN2(N1573));
and2s1 U395 (.Q(N2962), .DIN1(N307), .DIN2(N1573));
and2s1 U396 (.Q(N2963), .DIN1(N299), .DIN2(N1573));
hi1s1 U397 (.Q(N2964), .DIN(N1588));
and2s1 U398 (.Q(N2969), .DIN1(N83), .DIN2(N1588));
and2s1 U399 (.Q(N2970), .DIN1(N86), .DIN2(N1588));
and2s1 U400 (.Q(N2971), .DIN1(N88), .DIN2(N1588));
and2s1 U401 (.Q(N2972), .DIN1(N88), .DIN2(N1588));
hi1s1 U402 (.Q(N2973), .DIN(N1594));
hi1s1 U403 (.Q(N2974), .DIN(N1597));
hi1s1 U404 (.Q(N2975), .DIN(N1600));
hi1s1 U405 (.Q(N2976), .DIN(N1603));
hi1s1 U406 (.Q(N2977), .DIN(N1606));
hi1s1 U407 (.Q(N2978), .DIN(N1609));
and3s1 U408 (.Q(N2979), .DIN1(N1315), .DIN2(N503), .DIN3(N1597));
and2s1 U409 (.Q(N2980), .DIN1(N1315), .DIN2(N514));
and3s1 U410 (.Q(N2981), .DIN1(N1315), .DIN2(N523), .DIN3(N1603));
and3s1 U411 (.Q(N2982), .DIN1(N1315), .DIN2(N534), .DIN3(N1609));
and2s1 U412 (.Q(N2983), .DIN1(N1675), .DIN2(N1594));
or2s1 U413 (.Q(N2984), .DIN1(N1675), .DIN2(N514));
and2s1 U414 (.Q(N2985), .DIN1(N1675), .DIN2(N1600));
and2s1 U415 (.Q(N2986), .DIN1(N1675), .DIN2(N1606));
hi1s1 U416 (.Q(N2987), .DIN(N1612));
hi1s1 U417 (.Q(N2988), .DIN(N1615));
hi1s1 U418 (.Q(N2989), .DIN(N1618));
hi1s1 U419 (.Q(N2990), .DIN(N1621));
hi1s1 U420 (.Q(N2991), .DIN(N1624));
hi1s1 U421 (.Q(N2992), .DIN(N1627));
and2s1 U422 (.Q(N2993), .DIN1(N1315), .DIN2(N1615));
and3s1 U423 (.Q(N2994), .DIN1(N1315), .DIN2(N479), .DIN3(N1621));
and3s1 U424 (.Q(N2995), .DIN1(N1315), .DIN2(N490), .DIN3(N1627));
and2s1 U425 (.Q(N2996), .DIN1(N1675), .DIN2(N1612));
and2s1 U426 (.Q(N2997), .DIN1(N1675), .DIN2(N1618));
and2s1 U427 (.Q(N2998), .DIN1(N1675), .DIN2(N1624));
hi1s1 U428 (.Q(N2999), .DIN(N1630));
nb1s1 U429 (.Q(N3000), .DIN(N1469));
nb1s1 U430 (.Q(N3003), .DIN(N1469));
hi1s1 U431 (.Q(N3006), .DIN(N1633));
nb1s1 U432 (.Q(N3007), .DIN(N1469));
nb1s1 U433 (.Q(N3010), .DIN(N1469));
and2s1 U434 (.Q(N3013), .DIN1(N1315), .DIN2(N1630));
and2s1 U435 (.Q(N3014), .DIN1(N1315), .DIN2(N1633));
hi1s1 U436 (.Q(N3015), .DIN(N1636));
hi1s1 U437 (.Q(N3016), .DIN(N1639));
hi1s1 U438 (.Q(N3017), .DIN(N1642));
hi1s1 U439 (.Q(N3018), .DIN(N1645));
hi1s1 U440 (.Q(N3019), .DIN(N1648));
hi1s1 U441 (.Q(N3020), .DIN(N1651));
hi1s1 U442 (.Q(N3021), .DIN(N1654));
hi1s1 U443 (.Q(N3022), .DIN(N1657));
and3s1 U444 (.Q(N3023), .DIN1(N1303), .DIN2(N457), .DIN3(N1639));
and3s1 U445 (.Q(N3024), .DIN1(N1303), .DIN2(N468), .DIN3(N1645));
and3s1 U446 (.Q(N3025), .DIN1(N1303), .DIN2(N422), .DIN3(N1651));
and3s1 U447 (.Q(N3026), .DIN1(N1303), .DIN2(N435), .DIN3(N1657));
and2s1 U448 (.Q(N3027), .DIN1(N1663), .DIN2(N1636));
and2s1 U449 (.Q(N3028), .DIN1(N1663), .DIN2(N1642));
and2s1 U450 (.Q(N3029), .DIN1(N1663), .DIN2(N1648));
and2s1 U451 (.Q(N3030), .DIN1(N1663), .DIN2(N1654));
hi1s1 U452 (.Q(N3031), .DIN(N1920));
hi1s1 U453 (.Q(N3032), .DIN(N1923));
hi1s1 U454 (.Q(N3033), .DIN(N1926));
hi1s1 U455 (.Q(N3034), .DIN(N1929));
nb1s1 U456 (.Q(N3035), .DIN(N1660));
nb1s1 U457 (.Q(N3038), .DIN(N1660));
hi1s1 U458 (.Q(N3041), .DIN(N1697));
hi1s1 U459 (.Q(N3052), .DIN(N1709));
hi1s1 U460 (.Q(N3063), .DIN(N1721));
hi1s1 U461 (.Q(N3068), .DIN(N1727));
and2s1 U462 (.Q(N3071), .DIN1(N97), .DIN2(N1721));
and2s1 U463 (.Q(N3072), .DIN1(N94), .DIN2(N1721));
and2s1 U464 (.Q(N3073), .DIN1(N97), .DIN2(N1721));
and2s1 U465 (.Q(N3074), .DIN1(N94), .DIN2(N1721));
hi1s1 U466 (.Q(N3075), .DIN(N1731));
hi1s1 U467 (.Q(N3086), .DIN(N1743));
hi1s1 U468 (.Q(N3097), .DIN(N1761));
hi1s1 U469 (.Q(N3108), .DIN(N1769));
hi1s1 U470 (.Q(N3119), .DIN(N1777));
hi1s1 U471 (.Q(N3130), .DIN(N1785));
hi1s1 U472 (.Q(N3141), .DIN(N1944));
hi1s1 U473 (.Q(N3142), .DIN(N1947));
hi1s1 U474 (.Q(N3143), .DIN(N1950));
hi1s1 U475 (.Q(N3144), .DIN(N1953));
hi1s1 U476 (.Q(N3145), .DIN(N1956));
hi1s1 U477 (.Q(N3146), .DIN(N1959));
hi1s1 U478 (.Q(N3147), .DIN(N1793));
hi1s1 U479 (.Q(N3158), .DIN(N1800));
hi1s1 U480 (.Q(N3169), .DIN(N1807));
hi1s1 U481 (.Q(N3180), .DIN(N1814));
nb1s1 U482 (.Q(N3191), .DIN(N1821));
hi1s1 U483 (.Q(N3194), .DIN(N1932));
hi1s1 U484 (.Q(N3195), .DIN(N1935));
hi1s1 U485 (.Q(N3196), .DIN(N1938));
hi1s1 U486 (.Q(N3197), .DIN(N1941));
hi1s1 U487 (.Q(N3198), .DIN(N1962));
hi1s1 U488 (.Q(N3199), .DIN(N1965));
nb1s1 U489 (.Q(N3200), .DIN(N1469));
hi1s1 U490 (.Q(N3203), .DIN(N1968));
nb1s1 U491 (.Q(N3357), .DIN(N2704));
nb1s1 U492 (.Q(N3358), .DIN(N2704));
nb1s1 U493 (.Q(N3359), .DIN(N2704));
nb1s1 U494 (.Q(N3360), .DIN(N2704));
and3s1 U495 (.Q(N3401), .DIN1(N457), .DIN2(N1092), .DIN3(N2824));
and3s1 U496 (.Q(N3402), .DIN1(N468), .DIN2(N1092), .DIN3(N2826));
and3s1 U497 (.Q(N3403), .DIN1(N422), .DIN2(N1092), .DIN3(N2828));
and3s1 U498 (.Q(N3404), .DIN1(N435), .DIN2(N1092), .DIN3(N2830));
and2s1 U499 (.Q(N3405), .DIN1(N1080), .DIN2(N2823));
and2s1 U500 (.Q(N3406), .DIN1(N1080), .DIN2(N2825));
and2s1 U501 (.Q(N3407), .DIN1(N1080), .DIN2(N2827));
and2s1 U502 (.Q(N3408), .DIN1(N1080), .DIN2(N2829));
and3s1 U503 (.Q(N3409), .DIN1(N389), .DIN2(N1092), .DIN3(N2840));
and3s1 U504 (.Q(N3410), .DIN1(N400), .DIN2(N1092), .DIN3(N2842));
and3s1 U505 (.Q(N3411), .DIN1(N411), .DIN2(N1092), .DIN3(N2844));
and3s1 U506 (.Q(N3412), .DIN1(N374), .DIN2(N1092), .DIN3(N2846));
and2s1 U507 (.Q(N3413), .DIN1(N1080), .DIN2(N2839));
and2s1 U508 (.Q(N3414), .DIN1(N1080), .DIN2(N2841));
and2s1 U509 (.Q(N3415), .DIN1(N1080), .DIN2(N2843));
and2s1 U510 (.Q(N3416), .DIN1(N1080), .DIN2(N2845));
and2s1 U511 (.Q(N3444), .DIN1(N1280), .DIN2(N2902));
and3s1 U512 (.Q(N3445), .DIN1(N479), .DIN2(N1280), .DIN3(N2904));
and3s1 U513 (.Q(N3446), .DIN1(N490), .DIN2(N1280), .DIN3(N2906));
and2s1 U514 (.Q(N3447), .DIN1(N1685), .DIN2(N2901));
and2s1 U515 (.Q(N3448), .DIN1(N1685), .DIN2(N2903));
and2s1 U516 (.Q(N3449), .DIN1(N1685), .DIN2(N2905));
and3s1 U517 (.Q(N3450), .DIN1(N503), .DIN2(N1092), .DIN3(N2914));
and3s1 U518 (.Q(N3451), .DIN1(N523), .DIN2(N1092), .DIN3(N2916));
and3s1 U519 (.Q(N3452), .DIN1(N534), .DIN2(N1092), .DIN3(N2918));
and2s1 U520 (.Q(N3453), .DIN1(N1080), .DIN2(N2913));
and2s1 U521 (.Q(N3454), .DIN1(N1080), .DIN2(N2915));
and2s1 U522 (.Q(N3455), .DIN1(N1080), .DIN2(N2917));
and2s1 U523 (.Q(N3456), .DIN1(N2920), .DIN2(N2350));
and3s1 U524 (.Q(N3459), .DIN1(N389), .DIN2(N1280), .DIN3(N2927));
and3s1 U525 (.Q(N3460), .DIN1(N400), .DIN2(N1280), .DIN3(N2929));
and3s1 U526 (.Q(N3461), .DIN1(N411), .DIN2(N1280), .DIN3(N2931));
and3s1 U527 (.Q(N3462), .DIN1(N374), .DIN2(N1280), .DIN3(N2933));
and2s1 U528 (.Q(N3463), .DIN1(N1685), .DIN2(N2926));
and2s1 U529 (.Q(N3464), .DIN1(N1685), .DIN2(N2928));
and2s1 U530 (.Q(N3465), .DIN1(N1685), .DIN2(N2930));
and2s1 U531 (.Q(N3466), .DIN1(N1685), .DIN2(N2932));
and3s1 U532 (.Q(N3481), .DIN1(N503), .DIN2(N1292), .DIN3(N2974));
hi1s1 U533 (.Q(N3482), .DIN(N2980));
and3s1 U534 (.Q(N3483), .DIN1(N523), .DIN2(N1292), .DIN3(N2976));
and3s1 U535 (.Q(N3484), .DIN1(N534), .DIN2(N1292), .DIN3(N2978));
and2s1 U536 (.Q(N3485), .DIN1(N1271), .DIN2(N2973));
and2s1 U537 (.Q(N3486), .DIN1(N1271), .DIN2(N2975));
and2s1 U538 (.Q(N3487), .DIN1(N1271), .DIN2(N2977));
and2s1 U539 (.Q(N3488), .DIN1(N1292), .DIN2(N2988));
and3s1 U540 (.Q(N3489), .DIN1(N479), .DIN2(N1292), .DIN3(N2990));
and3s1 U541 (.Q(N3490), .DIN1(N490), .DIN2(N1292), .DIN3(N2992));
and2s1 U542 (.Q(N3491), .DIN1(N1271), .DIN2(N2987));
and2s1 U543 (.Q(N3492), .DIN1(N1271), .DIN2(N2989));
and2s1 U544 (.Q(N3493), .DIN1(N1271), .DIN2(N2991));
and2s1 U545 (.Q(N3502), .DIN1(N1292), .DIN2(N2999));
and2s1 U546 (.Q(N3503), .DIN1(N1292), .DIN2(N3006));
and3s1 U547 (.Q(N3504), .DIN1(N457), .DIN2(N1280), .DIN3(N3016));
and3s1 U548 (.Q(N3505), .DIN1(N468), .DIN2(N1280), .DIN3(N3018));
and3s1 U549 (.Q(N3506), .DIN1(N422), .DIN2(N1280), .DIN3(N3020));
and3s1 U550 (.Q(N3507), .DIN1(N435), .DIN2(N1280), .DIN3(N3022));
and2s1 U551 (.Q(N3508), .DIN1(N1685), .DIN2(N3015));
and2s1 U552 (.Q(N3509), .DIN1(N1685), .DIN2(N3017));
and2s1 U553 (.Q(N3510), .DIN1(N1685), .DIN2(N3019));
and2s1 U554 (.Q(N3511), .DIN1(N1685), .DIN2(N3021));
nnd2s1 U555 (.Q(N3512), .DIN1(N1923), .DIN2(N3031));
nnd2s1 U556 (.Q(N3513), .DIN1(N1920), .DIN2(N3032));
nnd2s1 U557 (.Q(N3514), .DIN1(N1929), .DIN2(N3033));
nnd2s1 U558 (.Q(N3515), .DIN1(N1926), .DIN2(N3034));
nnd2s1 U559 (.Q(N3558), .DIN1(N1947), .DIN2(N3141));
nnd2s1 U560 (.Q(N3559), .DIN1(N1944), .DIN2(N3142));
nnd2s1 U561 (.Q(N3560), .DIN1(N1953), .DIN2(N3143));
nnd2s1 U562 (.Q(N3561), .DIN1(N1950), .DIN2(N3144));
nnd2s1 U563 (.Q(N3562), .DIN1(N1959), .DIN2(N3145));
nnd2s1 U564 (.Q(N3563), .DIN1(N1956), .DIN2(N3146));
nb1s1 U565 (.Q(N3604), .DIN(N3191));
nnd2s1 U566 (.Q(N3605), .DIN1(N1935), .DIN2(N3194));
nnd2s1 U567 (.Q(N3606), .DIN1(N1932), .DIN2(N3195));
nnd2s1 U568 (.Q(N3607), .DIN1(N1941), .DIN2(N3196));
nnd2s1 U569 (.Q(N3608), .DIN1(N1938), .DIN2(N3197));
nnd2s1 U570 (.Q(N3609), .DIN1(N1965), .DIN2(N3198));
nnd2s1 U571 (.Q(N3610), .DIN1(N1962), .DIN2(N3199));
hi1s1 U572 (.Q(N3613), .DIN(N3191));
and2s1 U573 (.Q(N3614), .DIN1(N2882), .DIN2(N2891));
and2s1 U574 (.Q(N3615), .DIN1(N1482), .DIN2(N2891));
and3s1 U575 (.Q(N3616), .DIN1(N200), .DIN2(N2653), .DIN3(N1173));
and3s1 U576 (.Q(N3617), .DIN1(N203), .DIN2(N2653), .DIN3(N1173));
and3s1 U577 (.Q(N3618), .DIN1(N197), .DIN2(N2653), .DIN3(N1173));
and3s1 U578 (.Q(N3619), .DIN1(N194), .DIN2(N2653), .DIN3(N1173));
and3s1 U579 (.Q(N3620), .DIN1(N191), .DIN2(N2653), .DIN3(N1173));
and3s1 U580 (.Q(N3621), .DIN1(N182), .DIN2(N2681), .DIN3(N1197));
and3s1 U581 (.Q(N3622), .DIN1(N188), .DIN2(N2681), .DIN3(N1197));
and3s1 U582 (.Q(N3623), .DIN1(N155), .DIN2(N2681), .DIN3(N1197));
and3s1 U583 (.Q(N3624), .DIN1(N149), .DIN2(N2681), .DIN3(N1197));
and2s1 U584 (.Q(N3625), .DIN1(N2882), .DIN2(N2891));
and2s1 U585 (.Q(N3626), .DIN1(N1482), .DIN2(N2891));
and3s1 U586 (.Q(N3627), .DIN1(N200), .DIN2(N2728), .DIN3(N1235));
and3s1 U587 (.Q(N3628), .DIN1(N203), .DIN2(N2728), .DIN3(N1235));
and3s1 U588 (.Q(N3629), .DIN1(N197), .DIN2(N2728), .DIN3(N1235));
and3s1 U589 (.Q(N3630), .DIN1(N194), .DIN2(N2728), .DIN3(N1235));
and3s1 U590 (.Q(N3631), .DIN1(N191), .DIN2(N2728), .DIN3(N1235));
and3s1 U591 (.Q(N3632), .DIN1(N182), .DIN2(N2756), .DIN3(N1259));
and3s1 U592 (.Q(N3633), .DIN1(N188), .DIN2(N2756), .DIN3(N1259));
and3s1 U593 (.Q(N3634), .DIN1(N155), .DIN2(N2756), .DIN3(N1259));
and3s1 U594 (.Q(N3635), .DIN1(N149), .DIN2(N2756), .DIN3(N1259));
and2s1 U595 (.Q(N3636), .DIN1(N2882), .DIN2(N2891));
and2s1 U596 (.Q(N3637), .DIN1(N1482), .DIN2(N2891));
and3s1 U597 (.Q(N3638), .DIN1(N109), .DIN2(N3075), .DIN3(N1743));
and2s1 U598 (.Q(N3639), .DIN1(N2882), .DIN2(N2891));
and2s1 U599 (.Q(N3640), .DIN1(N1482), .DIN2(N2891));
and3s1 U600 (.Q(N3641), .DIN1(N11), .DIN2(N2779), .DIN3(N1339));
and3s1 U601 (.Q(N3642), .DIN1(N109), .DIN2(N3041), .DIN3(N1709));
and3s1 U602 (.Q(N3643), .DIN1(N46), .DIN2(N3041), .DIN3(N1709));
and3s1 U603 (.Q(N3644), .DIN1(N100), .DIN2(N3041), .DIN3(N1709));
and3s1 U604 (.Q(N3645), .DIN1(N91), .DIN2(N3041), .DIN3(N1709));
and3s1 U605 (.Q(N3646), .DIN1(N43), .DIN2(N3041), .DIN3(N1709));
and3s1 U606 (.Q(N3647), .DIN1(N76), .DIN2(N2779), .DIN3(N1339));
and3s1 U607 (.Q(N3648), .DIN1(N73), .DIN2(N2779), .DIN3(N1339));
and3s1 U608 (.Q(N3649), .DIN1(N67), .DIN2(N2779), .DIN3(N1339));
and3s1 U609 (.Q(N3650), .DIN1(N14), .DIN2(N2779), .DIN3(N1339));
and3s1 U610 (.Q(N3651), .DIN1(N46), .DIN2(N3075), .DIN3(N1743));
and3s1 U611 (.Q(N3652), .DIN1(N100), .DIN2(N3075), .DIN3(N1743));
and3s1 U612 (.Q(N3653), .DIN1(N91), .DIN2(N3075), .DIN3(N1743));
and3s1 U613 (.Q(N3654), .DIN1(N43), .DIN2(N3075), .DIN3(N1743));
and3s1 U614 (.Q(N3655), .DIN1(N76), .DIN2(N2801), .DIN3(N1363));
and3s1 U615 (.Q(N3656), .DIN1(N73), .DIN2(N2801), .DIN3(N1363));
and3s1 U616 (.Q(N3657), .DIN1(N67), .DIN2(N2801), .DIN3(N1363));
and3s1 U617 (.Q(N3658), .DIN1(N14), .DIN2(N2801), .DIN3(N1363));
and3s1 U618 (.Q(N3659), .DIN1(N120), .DIN2(N3119), .DIN3(N1785));
and3s1 U619 (.Q(N3660), .DIN1(N11), .DIN2(N2801), .DIN3(N1363));
and3s1 U620 (.Q(N3661), .DIN1(N118), .DIN2(N3097), .DIN3(N1769));
and3s1 U621 (.Q(N3662), .DIN1(N176), .DIN2(N2681), .DIN3(N1197));
and3s1 U622 (.Q(N3663), .DIN1(N176), .DIN2(N2756), .DIN3(N1259));
or2s1 U623 (.Q(N3664), .DIN1(N2831), .DIN2(N3401));
or2s1 U624 (.Q(N3665), .DIN1(N2832), .DIN2(N3402));
or2s1 U625 (.Q(N3666), .DIN1(N2833), .DIN2(N3403));
or2s1 U626 (.Q(N3667), .DIN1(N2834), .DIN2(N3404));
or3s1 U627 (.Q(N3668), .DIN1(N2835), .DIN2(N3405), .DIN3(N457));
or3s1 U628 (.Q(N3669), .DIN1(N2836), .DIN2(N3406), .DIN3(N468));
or3s1 U629 (.Q(N3670), .DIN1(N2837), .DIN2(N3407), .DIN3(N422));
or3s1 U630 (.Q(N3671), .DIN1(N2838), .DIN2(N3408), .DIN3(N435));
or2s1 U631 (.Q(N3672), .DIN1(N2847), .DIN2(N3409));
or2s1 U632 (.Q(N3673), .DIN1(N2848), .DIN2(N3410));
or2s1 U633 (.Q(N3674), .DIN1(N2849), .DIN2(N3411));
or2s1 U634 (.Q(N3675), .DIN1(N2850), .DIN2(N3412));
or3s1 U635 (.Q(N3676), .DIN1(N2851), .DIN2(N3413), .DIN3(N389));
or3s1 U636 (.Q(N3677), .DIN1(N2852), .DIN2(N3414), .DIN3(N400));
or3s1 U637 (.Q(N3678), .DIN1(N2853), .DIN2(N3415), .DIN3(N411));
or3s1 U638 (.Q(N3679), .DIN1(N2854), .DIN2(N3416), .DIN3(N374));
and2s1 U639 (.Q(N3680), .DIN1(N289), .DIN2(N2855));
and2s1 U640 (.Q(N3681), .DIN1(N281), .DIN2(N2855));
and2s1 U641 (.Q(N3682), .DIN1(N273), .DIN2(N2855));
and2s1 U642 (.Q(N3683), .DIN1(N265), .DIN2(N2855));
and2s1 U643 (.Q(N3684), .DIN1(N257), .DIN2(N2855));
and2s1 U644 (.Q(N3685), .DIN1(N234), .DIN2(N2861));
and2s1 U645 (.Q(N3686), .DIN1(N226), .DIN2(N2861));
and2s1 U646 (.Q(N3687), .DIN1(N218), .DIN2(N2861));
and2s1 U647 (.Q(N3688), .DIN1(N210), .DIN2(N2861));
and2s1 U648 (.Q(N3689), .DIN1(N206), .DIN2(N2861));
hi1s1 U649 (.Q(N3691), .DIN(N2891));
or2s1 U650 (.Q(N3700), .DIN1(N2907), .DIN2(N3444));
or2s1 U651 (.Q(N3701), .DIN1(N2908), .DIN2(N3445));
or2s1 U652 (.Q(N3702), .DIN1(N2909), .DIN2(N3446));
or3s1 U653 (.Q(N3703), .DIN1(N2911), .DIN2(N3448), .DIN3(N479));
or3s1 U654 (.Q(N3704), .DIN1(N2912), .DIN2(N3449), .DIN3(N490));
or2s1 U655 (.Q(N3705), .DIN1(N2910), .DIN2(N3447));
or2s1 U656 (.Q(N3708), .DIN1(N2919), .DIN2(N3450));
or2s1 U657 (.Q(N3709), .DIN1(N2921), .DIN2(N3451));
or2s1 U658 (.Q(N3710), .DIN1(N2922), .DIN2(N3452));
or3s1 U659 (.Q(N3711), .DIN1(N2923), .DIN2(N3453), .DIN3(N503));
or3s1 U660 (.Q(N3712), .DIN1(N2924), .DIN2(N3454), .DIN3(N523));
or3s1 U661 (.Q(N3713), .DIN1(N2925), .DIN2(N3455), .DIN3(N534));
or2s1 U662 (.Q(N3715), .DIN1(N2934), .DIN2(N3459));
or2s1 U663 (.Q(N3716), .DIN1(N2935), .DIN2(N3460));
or2s1 U664 (.Q(N3717), .DIN1(N2936), .DIN2(N3461));
or2s1 U665 (.Q(N3718), .DIN1(N2937), .DIN2(N3462));
or3s1 U666 (.Q(N3719), .DIN1(N2938), .DIN2(N3463), .DIN3(N389));
or3s1 U667 (.Q(N3720), .DIN1(N2939), .DIN2(N3464), .DIN3(N400));
or3s1 U668 (.Q(N3721), .DIN1(N2940), .DIN2(N3465), .DIN3(N411));
or3s1 U669 (.Q(N3722), .DIN1(N2941), .DIN2(N3466), .DIN3(N374));
and2s1 U670 (.Q(N3723), .DIN1(N369), .DIN2(N2942));
and2s1 U671 (.Q(N3724), .DIN1(N361), .DIN2(N2942));
and2s1 U672 (.Q(N3725), .DIN1(N351), .DIN2(N2942));
and2s1 U673 (.Q(N3726), .DIN1(N341), .DIN2(N2942));
and2s1 U674 (.Q(N3727), .DIN1(N324), .DIN2(N2948));
and2s1 U675 (.Q(N3728), .DIN1(N316), .DIN2(N2948));
and2s1 U676 (.Q(N3729), .DIN1(N308), .DIN2(N2948));
and2s1 U677 (.Q(N3730), .DIN1(N302), .DIN2(N2948));
and2s1 U678 (.Q(N3731), .DIN1(N293), .DIN2(N2948));
or2s1 U679 (.Q(N3732), .DIN1(N2942), .DIN2(N2958));
and2s1 U680 (.Q(N3738), .DIN1(N83), .DIN2(N2964));
and2s1 U681 (.Q(N3739), .DIN1(N87), .DIN2(N2964));
and2s1 U682 (.Q(N3740), .DIN1(N34), .DIN2(N2964));
and2s1 U683 (.Q(N3741), .DIN1(N34), .DIN2(N2964));
or2s1 U684 (.Q(N3742), .DIN1(N2979), .DIN2(N3481));
or2s1 U685 (.Q(N3743), .DIN1(N2981), .DIN2(N3483));
or2s1 U686 (.Q(N3744), .DIN1(N2982), .DIN2(N3484));
or3s1 U687 (.Q(N3745), .DIN1(N2983), .DIN2(N3485), .DIN3(N503));
or3s1 U688 (.Q(N3746), .DIN1(N2985), .DIN2(N3486), .DIN3(N523));
or3s1 U689 (.Q(N3747), .DIN1(N2986), .DIN2(N3487), .DIN3(N534));
or2s1 U690 (.Q(N3748), .DIN1(N2993), .DIN2(N3488));
or2s1 U691 (.Q(N3749), .DIN1(N2994), .DIN2(N3489));
or2s1 U692 (.Q(N3750), .DIN1(N2995), .DIN2(N3490));
or3s1 U693 (.Q(N3751), .DIN1(N2997), .DIN2(N3492), .DIN3(N479));
or3s1 U694 (.Q(N3752), .DIN1(N2998), .DIN2(N3493), .DIN3(N490));
hi1s1 U695 (.Q(N3753), .DIN(N3000));
hi1s1 U696 (.Q(N3754), .DIN(N3003));
hi1s1 U697 (.Q(N3755), .DIN(N3007));
hi1s1 U698 (.Q(N3756), .DIN(N3010));
or2s1 U699 (.Q(N3757), .DIN1(N3013), .DIN2(N3502));
and3s1 U700 (.Q(N3758), .DIN1(N1315), .DIN2(N446), .DIN3(N3003));
or2s1 U701 (.Q(N3759), .DIN1(N3014), .DIN2(N3503));
and3s1 U702 (.Q(N3760), .DIN1(N1315), .DIN2(N446), .DIN3(N3010));
and2s1 U703 (.Q(N3761), .DIN1(N1675), .DIN2(N3000));
and2s1 U704 (.Q(N3762), .DIN1(N1675), .DIN2(N3007));
or2s1 U705 (.Q(N3763), .DIN1(N3023), .DIN2(N3504));
or2s1 U706 (.Q(N3764), .DIN1(N3024), .DIN2(N3505));
or2s1 U707 (.Q(N3765), .DIN1(N3025), .DIN2(N3506));
or2s1 U708 (.Q(N3766), .DIN1(N3026), .DIN2(N3507));
or3s1 U709 (.Q(N3767), .DIN1(N3027), .DIN2(N3508), .DIN3(N457));
or3s1 U710 (.Q(N3768), .DIN1(N3028), .DIN2(N3509), .DIN3(N468));
or3s1 U711 (.Q(N3769), .DIN1(N3029), .DIN2(N3510), .DIN3(N422));
or3s1 U712 (.Q(N3770), .DIN1(N3030), .DIN2(N3511), .DIN3(N435));
nnd2s1 U713 (.Q(N3771), .DIN1(N3512), .DIN2(N3513));
nnd2s1 U714 (.Q(N3775), .DIN1(N3514), .DIN2(N3515));
hi1s1 U715 (.Q(N3779), .DIN(N3035));
hi1s1 U716 (.Q(N3780), .DIN(N3038));
and3s1 U717 (.Q(N3781), .DIN1(N117), .DIN2(N3097), .DIN3(N1769));
and3s1 U718 (.Q(N3782), .DIN1(N126), .DIN2(N3097), .DIN3(N1769));
and3s1 U719 (.Q(N3783), .DIN1(N127), .DIN2(N3097), .DIN3(N1769));
and3s1 U720 (.Q(N3784), .DIN1(N128), .DIN2(N3097), .DIN3(N1769));
and3s1 U721 (.Q(N3785), .DIN1(N131), .DIN2(N3119), .DIN3(N1785));
and3s1 U722 (.Q(N3786), .DIN1(N129), .DIN2(N3119), .DIN3(N1785));
and3s1 U723 (.Q(N3787), .DIN1(N119), .DIN2(N3119), .DIN3(N1785));
and3s1 U724 (.Q(N3788), .DIN1(N130), .DIN2(N3119), .DIN3(N1785));
nnd2s1 U725 (.Q(N3789), .DIN1(N3558), .DIN2(N3559));
nnd2s1 U726 (.Q(N3793), .DIN1(N3560), .DIN2(N3561));
nnd2s1 U727 (.Q(N3797), .DIN1(N3562), .DIN2(N3563));
and3s1 U728 (.Q(N3800), .DIN1(N122), .DIN2(N3147), .DIN3(N1800));
and3s1 U729 (.Q(N3801), .DIN1(N113), .DIN2(N3147), .DIN3(N1800));
and3s1 U730 (.Q(N3802), .DIN1(N53), .DIN2(N3147), .DIN3(N1800));
and3s1 U731 (.Q(N3803), .DIN1(N114), .DIN2(N3147), .DIN3(N1800));
and3s1 U732 (.Q(N3804), .DIN1(N115), .DIN2(N3147), .DIN3(N1800));
and3s1 U733 (.Q(N3805), .DIN1(N52), .DIN2(N3169), .DIN3(N1814));
and3s1 U734 (.Q(N3806), .DIN1(N112), .DIN2(N3169), .DIN3(N1814));
and3s1 U735 (.Q(N3807), .DIN1(N116), .DIN2(N3169), .DIN3(N1814));
and3s1 U736 (.Q(N3808), .DIN1(N121), .DIN2(N3169), .DIN3(N1814));
and3s1 U737 (.Q(N3809), .DIN1(N123), .DIN2(N3169), .DIN3(N1814));
nnd2s1 U738 (.Q(N3810), .DIN1(N3607), .DIN2(N3608));
nnd2s1 U739 (.Q(N3813), .DIN1(N3605), .DIN2(N3606));
and2s1 U740 (.Q(N3816), .DIN1(N3482), .DIN2(N2984));
or2s1 U741 (.Q(N3819), .DIN1(N2996), .DIN2(N3491));
hi1s1 U742 (.Q(N3822), .DIN(N3200));
nnd2s1 U743 (.Q(N3823), .DIN1(N3200), .DIN2(N3203));
nnd2s1 U744 (.Q(N3824), .DIN1(N3609), .DIN2(N3610));
hi1s1 U745 (.Q(N3827), .DIN(N3456));
or2s1 U746 (.Q(N3828), .DIN1(N3739), .DIN2(N2970));
or2s1 U747 (.Q(N3829), .DIN1(N3740), .DIN2(N2971));
or2s1 U748 (.Q(N3830), .DIN1(N3741), .DIN2(N2972));
or2s1 U749 (.Q(N3831), .DIN1(N3738), .DIN2(N2969));
hi1s1 U750 (.Q(N3834), .DIN(N3664));
hi1s1 U751 (.Q(N3835), .DIN(N3665));
hi1s1 U752 (.Q(N3836), .DIN(N3666));
hi1s1 U753 (.Q(N3837), .DIN(N3667));
hi1s1 U754 (.Q(N3838), .DIN(N3672));
hi1s1 U755 (.Q(N3839), .DIN(N3673));
hi1s1 U756 (.Q(N3840), .DIN(N3674));
hi1s1 U757 (.Q(N3841), .DIN(N3675));
or2s1 U758 (.Q(N3842), .DIN1(N3681), .DIN2(N2868));
or2s1 U759 (.Q(N3849), .DIN1(N3682), .DIN2(N2869));
or2s1 U760 (.Q(N3855), .DIN1(N3683), .DIN2(N2870));
or2s1 U761 (.Q(N3861), .DIN1(N3684), .DIN2(N2871));
or2s1 U762 (.Q(N3867), .DIN1(N3685), .DIN2(N2872));
or2s1 U763 (.Q(N3873), .DIN1(N3686), .DIN2(N2873));
or2s1 U764 (.Q(N3881), .DIN1(N3687), .DIN2(N2874));
or2s1 U765 (.Q(N3887), .DIN1(N3688), .DIN2(N2875));
or2s1 U766 (.Q(N3893), .DIN1(N3689), .DIN2(N2876));
hi1s1 U767 (.Q(N3908), .DIN(N3701));
hi1s1 U768 (.Q(N3909), .DIN(N3702));
hi1s1 U769 (.Q(N3911), .DIN(N3700));
hi1s1 U770 (.Q(N3914), .DIN(N3708));
hi1s1 U771 (.Q(N3915), .DIN(N3709));
hi1s1 U772 (.Q(N3916), .DIN(N3710));
hi1s1 U773 (.Q(N3917), .DIN(N3715));
hi1s1 U774 (.Q(N3918), .DIN(N3716));
hi1s1 U775 (.Q(N3919), .DIN(N3717));
hi1s1 U776 (.Q(N3920), .DIN(N3718));
or2s1 U777 (.Q(N3921), .DIN1(N3724), .DIN2(N2955));
or2s1 U778 (.Q(N3927), .DIN1(N3725), .DIN2(N2956));
or2s1 U779 (.Q(N3933), .DIN1(N3726), .DIN2(N2957));
or2s1 U780 (.Q(N3942), .DIN1(N3727), .DIN2(N2959));
or2s1 U781 (.Q(N3948), .DIN1(N3728), .DIN2(N2960));
or2s1 U782 (.Q(N3956), .DIN1(N3729), .DIN2(N2961));
or2s1 U783 (.Q(N3962), .DIN1(N3730), .DIN2(N2962));
or2s1 U784 (.Q(N3968), .DIN1(N3731), .DIN2(N2963));
hi1s1 U785 (.Q(N3975), .DIN(N3742));
hi1s1 U786 (.Q(N3976), .DIN(N3743));
hi1s1 U787 (.Q(N3977), .DIN(N3744));
hi1s1 U788 (.Q(N3978), .DIN(N3749));
hi1s1 U789 (.Q(N3979), .DIN(N3750));
and3s1 U790 (.Q(N3980), .DIN1(N446), .DIN2(N1292), .DIN3(N3754));
and3s1 U791 (.Q(N3981), .DIN1(N446), .DIN2(N1292), .DIN3(N3756));
and2s1 U792 (.Q(N3982), .DIN1(N1271), .DIN2(N3753));
and2s1 U793 (.Q(N3983), .DIN1(N1271), .DIN2(N3755));
hi1s1 U794 (.Q(N3984), .DIN(N3757));
hi1s1 U795 (.Q(N3987), .DIN(N3759));
hi1s1 U796 (.Q(N3988), .DIN(N3763));
hi1s1 U797 (.Q(N3989), .DIN(N3764));
hi1s1 U798 (.Q(N3990), .DIN(N3765));
hi1s1 U799 (.Q(N3991), .DIN(N3766));
and3s1 U800 (.Q(N3998), .DIN1(N3456), .DIN2(N3119), .DIN3(N3130));
or2s1 U801 (.Q(N4008), .DIN1(N3723), .DIN2(N2954));
or2s1 U802 (.Q(N4011), .DIN1(N3680), .DIN2(N2867));
hi1s1 U803 (.Q(N4021), .DIN(N3748));
nnd2s1 U804 (.Q(N4024), .DIN1(N1968), .DIN2(N3822));
hi1s1 U805 (.Q(N4027), .DIN(N3705));
and2s1 U806 (.Q(N4031), .DIN1(N3828), .DIN2(N1583));
and3s1 U807 (.Q(N4032), .DIN1(N24), .DIN2(N2882), .DIN3(N3691));
and3s1 U808 (.Q(N4033), .DIN1(N25), .DIN2(N1482), .DIN3(N3691));
and3s1 U809 (.Q(N4034), .DIN1(N26), .DIN2(N2882), .DIN3(N3691));
and3s1 U810 (.Q(N4035), .DIN1(N81), .DIN2(N1482), .DIN3(N3691));
and2s1 U811 (.Q(N4036), .DIN1(N3829), .DIN2(N1583));
and3s1 U812 (.Q(N4037), .DIN1(N79), .DIN2(N2882), .DIN3(N3691));
and3s1 U813 (.Q(N4038), .DIN1(N23), .DIN2(N1482), .DIN3(N3691));
and3s1 U814 (.Q(N4039), .DIN1(N82), .DIN2(N2882), .DIN3(N3691));
and3s1 U815 (.Q(N4040), .DIN1(N80), .DIN2(N1482), .DIN3(N3691));
and2s1 U816 (.Q(N4041), .DIN1(N3830), .DIN2(N1583));
and2s1 U817 (.Q(N4042), .DIN1(N3831), .DIN2(N1583));
and2s1 U818 (.Q(N4067), .DIN1(N3732), .DIN2(N514));
and2s1 U819 (.Q(N4080), .DIN1(N514), .DIN2(N3732));
and2s1 U820 (.Q(N4088), .DIN1(N3834), .DIN2(N3668));
and2s1 U821 (.Q(N4091), .DIN1(N3835), .DIN2(N3669));
and2s1 U822 (.Q(N4094), .DIN1(N3836), .DIN2(N3670));
and2s1 U823 (.Q(N4097), .DIN1(N3837), .DIN2(N3671));
and2s1 U824 (.Q(N4100), .DIN1(N3838), .DIN2(N3676));
and2s1 U825 (.Q(N4103), .DIN1(N3839), .DIN2(N3677));
and2s1 U826 (.Q(N4106), .DIN1(N3840), .DIN2(N3678));
and2s1 U827 (.Q(N4109), .DIN1(N3841), .DIN2(N3679));
and2s1 U828 (.Q(N4144), .DIN1(N3908), .DIN2(N3703));
and2s1 U829 (.Q(N4147), .DIN1(N3909), .DIN2(N3704));
nb1s1 U830 (.Q(N4150), .DIN(N3705));
and2s1 U831 (.Q(N4153), .DIN1(N3914), .DIN2(N3711));
and2s1 U832 (.Q(N4156), .DIN1(N3915), .DIN2(N3712));
and2s1 U833 (.Q(N4159), .DIN1(N3916), .DIN2(N3713));
or2s1 U834 (.Q(N4183), .DIN1(N3758), .DIN2(N3980));
or2s1 U835 (.Q(N4184), .DIN1(N3760), .DIN2(N3981));
or3s1 U836 (.Q(N4185), .DIN1(N3761), .DIN2(N3982), .DIN3(N446));
or3s1 U837 (.Q(N4186), .DIN1(N3762), .DIN2(N3983), .DIN3(N446));
hi1s1 U838 (.Q(N4188), .DIN(N3771));
hi1s1 U839 (.Q(N4191), .DIN(N3775));
and3s1 U840 (.Q(N4196), .DIN1(N3775), .DIN2(N3771), .DIN3(N3035));
and3s1 U841 (.Q(N4197), .DIN1(N3987), .DIN2(N3119), .DIN3(N3130));
and2s1 U842 (.Q(N4198), .DIN1(N3920), .DIN2(N3722));
hi1s1 U843 (.Q(N4199), .DIN(N3816));
hi1s1 U844 (.Q(N4200), .DIN(N3789));
hi1s1 U845 (.Q(N4203), .DIN(N3793));
nb1s1 U846 (.Q(N4206), .DIN(N3797));
nb1s1 U847 (.Q(N4209), .DIN(N3797));
nb1s1 U848 (.Q(N4212), .DIN(N3732));
nb1s1 U849 (.Q(N4215), .DIN(N3732));
nb1s1 U850 (.Q(N4219), .DIN(N3732));
hi1s1 U851 (.Q(N4223), .DIN(N3810));
hi1s1 U852 (.Q(N4224), .DIN(N3813));
and2s1 U853 (.Q(N4225), .DIN1(N3918), .DIN2(N3720));
and2s1 U854 (.Q(N4228), .DIN1(N3919), .DIN2(N3721));
and2s1 U855 (.Q(N4231), .DIN1(N3991), .DIN2(N3770));
and2s1 U856 (.Q(N4234), .DIN1(N3917), .DIN2(N3719));
and2s1 U857 (.Q(N4237), .DIN1(N3989), .DIN2(N3768));
and2s1 U858 (.Q(N4240), .DIN1(N3990), .DIN2(N3769));
and2s1 U859 (.Q(N4243), .DIN1(N3988), .DIN2(N3767));
and2s1 U860 (.Q(N4246), .DIN1(N3976), .DIN2(N3746));
and2s1 U861 (.Q(N4249), .DIN1(N3977), .DIN2(N3747));
and2s1 U862 (.Q(N4252), .DIN1(N3975), .DIN2(N3745));
and2s1 U863 (.Q(N4255), .DIN1(N3978), .DIN2(N3751));
and2s1 U864 (.Q(N4258), .DIN1(N3979), .DIN2(N3752));
hi1s1 U865 (.Q(N4263), .DIN(N3819));
nnd2s1 U866 (.Q(N4264), .DIN1(N4024), .DIN2(N3823));
hi1s1 U867 (.Q(N4267), .DIN(N3824));
and2s1 U868 (.Q(N4268), .DIN1(N446), .DIN2(N3893));
hi1s1 U869 (.Q(N4269), .DIN(N3911));
hi1s1 U870 (.Q(N4270), .DIN(N3984));
and2s1 U871 (.Q(N4271), .DIN1(N3893), .DIN2(N446));
hi1s1 U872 (.Q(N4272), .DIN(N4031));
or4s1 U873 (.Q(N4273), .DIN1(N4032), .DIN2(N4033), .DIN3(N3614), .DIN4(N3615));
or4s1 U874 (.Q(N4274), .DIN1(N4034), .DIN2(N4035), .DIN3(N3625), .DIN4(N3626));
hi1s1 U875 (.Q(N4275), .DIN(N4036));
or4s1 U876 (.Q(N4276), .DIN1(N4037), .DIN2(N4038), .DIN3(N3636), .DIN4(N3637));
or4s1 U877 (.Q(N4277), .DIN1(N4039), .DIN2(N4040), .DIN3(N3639), .DIN4(N3640));
hi1s1 U878 (.Q(N4278), .DIN(N4041));
hi1s1 U879 (.Q(N4279), .DIN(N4042));
and2s1 U880 (.Q(N4280), .DIN1(N3887), .DIN2(N457));
and2s1 U881 (.Q(N4284), .DIN1(N3881), .DIN2(N468));
and2s1 U882 (.Q(N4290), .DIN1(N422), .DIN2(N3873));
and2s1 U883 (.Q(N4297), .DIN1(N3867), .DIN2(N435));
and2s1 U884 (.Q(N4298), .DIN1(N3861), .DIN2(N389));
and2s1 U885 (.Q(N4301), .DIN1(N3855), .DIN2(N400));
and2s1 U886 (.Q(N4305), .DIN1(N3849), .DIN2(N411));
and2s1 U887 (.Q(N4310), .DIN1(N3842), .DIN2(N374));
and2s1 U888 (.Q(N4316), .DIN1(N457), .DIN2(N3887));
and2s1 U889 (.Q(N4320), .DIN1(N468), .DIN2(N3881));
and2s1 U890 (.Q(N4325), .DIN1(N422), .DIN2(N3873));
and2s1 U891 (.Q(N4331), .DIN1(N435), .DIN2(N3867));
and2s1 U892 (.Q(N4332), .DIN1(N389), .DIN2(N3861));
and2s1 U893 (.Q(N4336), .DIN1(N400), .DIN2(N3855));
and2s1 U894 (.Q(N4342), .DIN1(N411), .DIN2(N3849));
and2s1 U895 (.Q(N4349), .DIN1(N374), .DIN2(N3842));
hi1s1 U896 (.Q(N4357), .DIN(N3968));
hi1s1 U897 (.Q(N4364), .DIN(N3962));
nb1s1 U898 (.Q(N4375), .DIN(N3962));
and2s1 U899 (.Q(N4379), .DIN1(N3956), .DIN2(N479));
and2s1 U900 (.Q(N4385), .DIN1(N490), .DIN2(N3948));
and2s1 U901 (.Q(N4392), .DIN1(N3942), .DIN2(N503));
and2s1 U902 (.Q(N4396), .DIN1(N3933), .DIN2(N523));
and2s1 U903 (.Q(N4400), .DIN1(N3927), .DIN2(N534));
hi1s1 U904 (.Q(N4405), .DIN(N3921));
nb1s1 U905 (.Q(N4412), .DIN(N3921));
hi1s1 U906 (.Q(N4418), .DIN(N3968));
hi1s1 U907 (.Q(N4425), .DIN(N3962));
nb1s1 U908 (.Q(N4436), .DIN(N3962));
and2s1 U909 (.Q(N4440), .DIN1(N479), .DIN2(N3956));
and2s1 U910 (.Q(N4445), .DIN1(N490), .DIN2(N3948));
and2s1 U911 (.Q(N4451), .DIN1(N503), .DIN2(N3942));
and2s1 U912 (.Q(N4456), .DIN1(N523), .DIN2(N3933));
and2s1 U913 (.Q(N4462), .DIN1(N534), .DIN2(N3927));
nb1s1 U914 (.Q(N4469), .DIN(N3921));
hi1s1 U915 (.Q(N4477), .DIN(N3921));
nb1s1 U916 (.Q(N4512), .DIN(N3968));
hi1s1 U917 (.Q(N4515), .DIN(N4183));
hi1s1 U918 (.Q(N4516), .DIN(N4184));
hi1s1 U919 (.Q(N4521), .DIN(N4008));
hi1s1 U920 (.Q(N4523), .DIN(N4011));
hi1s1 U921 (.Q(N4524), .DIN(N4198));
hi1s1 U922 (.Q(N4532), .DIN(N3984));
and3s1 U923 (.Q(N4547), .DIN1(N3911), .DIN2(N3169), .DIN3(N3180));
nb1s1 U924 (.Q(N4548), .DIN(N3893));
nb1s1 U925 (.Q(N4551), .DIN(N3887));
nb1s1 U926 (.Q(N4554), .DIN(N3881));
nb1s1 U927 (.Q(N4557), .DIN(N3873));
nb1s1 U928 (.Q(N4560), .DIN(N3867));
nb1s1 U929 (.Q(N4563), .DIN(N3861));
nb1s1 U930 (.Q(N4566), .DIN(N3855));
nb1s1 U931 (.Q(N4569), .DIN(N3849));
nb1s1 U932 (.Q(N4572), .DIN(N3842));
nor2s1 U933 (.Q(N4575), .DIN1(N422), .DIN2(N3873));
nb1s1 U934 (.Q(N4578), .DIN(N3893));
nb1s1 U935 (.Q(N4581), .DIN(N3887));
nb1s1 U936 (.Q(N4584), .DIN(N3881));
nb1s1 U937 (.Q(N4587), .DIN(N3867));
nb1s1 U938 (.Q(N4590), .DIN(N3861));
nb1s1 U939 (.Q(N4593), .DIN(N3855));
nb1s1 U940 (.Q(N4596), .DIN(N3849));
nb1s1 U941 (.Q(N4599), .DIN(N3873));
nb1s1 U942 (.Q(N4602), .DIN(N3842));
nor2s1 U943 (.Q(N4605), .DIN1(N422), .DIN2(N3873));
nor2s1 U944 (.Q(N4608), .DIN1(N374), .DIN2(N3842));
nb1s1 U945 (.Q(N4611), .DIN(N3956));
nb1s1 U946 (.Q(N4614), .DIN(N3948));
nb1s1 U947 (.Q(N4617), .DIN(N3942));
nb1s1 U948 (.Q(N4621), .DIN(N3933));
nb1s1 U949 (.Q(N4624), .DIN(N3927));
nor2s1 U950 (.Q(N4627), .DIN1(N490), .DIN2(N3948));
nb1s1 U951 (.Q(N4630), .DIN(N3956));
nb1s1 U952 (.Q(N4633), .DIN(N3942));
nb1s1 U953 (.Q(N4637), .DIN(N3933));
nb1s1 U954 (.Q(N4640), .DIN(N3927));
nb1s1 U955 (.Q(N4643), .DIN(N3948));
nor2s1 U956 (.Q(N4646), .DIN1(N490), .DIN2(N3948));
nb1s1 U957 (.Q(N4649), .DIN(N3927));
nb1s1 U958 (.Q(N4652), .DIN(N3933));
nb1s1 U959 (.Q(N4655), .DIN(N3921));
nb1s1 U960 (.Q(N4658), .DIN(N3942));
nb1s1 U961 (.Q(N4662), .DIN(N3956));
nb1s1 U962 (.Q(N4665), .DIN(N3948));
nb1s1 U963 (.Q(N4668), .DIN(N3968));
nb1s1 U964 (.Q(N4671), .DIN(N3962));
nb1s1 U965 (.Q(N4674), .DIN(N3873));
nb1s1 U966 (.Q(N4677), .DIN(N3867));
nb1s1 U967 (.Q(N4680), .DIN(N3887));
nb1s1 U968 (.Q(N4683), .DIN(N3881));
nb1s1 U969 (.Q(N4686), .DIN(N3893));
nb1s1 U970 (.Q(N4689), .DIN(N3849));
nb1s1 U971 (.Q(N4692), .DIN(N3842));
nb1s1 U972 (.Q(N4695), .DIN(N3861));
nb1s1 U973 (.Q(N4698), .DIN(N3855));
nnd2s1 U974 (.Q(N4701), .DIN1(N3813), .DIN2(N4223));
nnd2s1 U975 (.Q(N4702), .DIN1(N3810), .DIN2(N4224));
hi1s1 U976 (.Q(N4720), .DIN(N4021));
nnd2s1 U977 (.Q(N4721), .DIN1(N4021), .DIN2(N4263));
hi1s1 U978 (.Q(N4724), .DIN(N4147));
hi1s1 U979 (.Q(N4725), .DIN(N4144));
hi1s1 U980 (.Q(N4726), .DIN(N4159));
hi1s1 U981 (.Q(N4727), .DIN(N4156));
hi1s1 U982 (.Q(N4728), .DIN(N4153));
hi1s1 U983 (.Q(N4729), .DIN(N4097));
hi1s1 U984 (.Q(N4730), .DIN(N4094));
hi1s1 U985 (.Q(N4731), .DIN(N4091));
hi1s1 U986 (.Q(N4732), .DIN(N4088));
hi1s1 U987 (.Q(N4733), .DIN(N4109));
hi1s1 U988 (.Q(N4734), .DIN(N4106));
hi1s1 U989 (.Q(N4735), .DIN(N4103));
hi1s1 U990 (.Q(N4736), .DIN(N4100));
and2s1 U991 (.Q(N4737), .DIN1(N4273), .DIN2(N2877));
and2s1 U992 (.Q(N4738), .DIN1(N4274), .DIN2(N2877));
and2s1 U993 (.Q(N4739), .DIN1(N4276), .DIN2(N2877));
and2s1 U994 (.Q(N4740), .DIN1(N4277), .DIN2(N2877));
and3s1 U995 (.Q(N4741), .DIN1(N4150), .DIN2(N1758), .DIN3(N1755));
hi1s1 U996 (.Q(N4855), .DIN(N4212));
nnd2s1 U997 (.Q(N4856), .DIN1(N4212), .DIN2(N2712));
nnd2s1 U998 (.Q(N4908), .DIN1(N4215), .DIN2(N2718));
hi1s1 U999 (.Q(N4909), .DIN(N4215));
and2s1 U1000 (.Q(N4939), .DIN1(N4515), .DIN2(N4185));
and2s1 U1001 (.Q(N4942), .DIN1(N4516), .DIN2(N4186));
hi1s1 U1002 (.Q(N4947), .DIN(N4219));
and3s1 U1003 (.Q(N4953), .DIN1(N4188), .DIN2(N3775), .DIN3(N3779));
and3s1 U1004 (.Q(N4954), .DIN1(N3771), .DIN2(N4191), .DIN3(N3780));
and3s1 U1005 (.Q(N4955), .DIN1(N4191), .DIN2(N4188), .DIN3(N3038));
and3s1 U1006 (.Q(N4956), .DIN1(N4109), .DIN2(N3097), .DIN3(N3108));
and3s1 U1007 (.Q(N4957), .DIN1(N4106), .DIN2(N3097), .DIN3(N3108));
and3s1 U1008 (.Q(N4958), .DIN1(N4103), .DIN2(N3097), .DIN3(N3108));
and3s1 U1009 (.Q(N4959), .DIN1(N4100), .DIN2(N3097), .DIN3(N3108));
and3s1 U1010 (.Q(N4960), .DIN1(N4159), .DIN2(N3119), .DIN3(N3130));
and3s1 U1011 (.Q(N4961), .DIN1(N4156), .DIN2(N3119), .DIN3(N3130));
hi1s1 U1012 (.Q(N4965), .DIN(N4225));
hi1s1 U1013 (.Q(N4966), .DIN(N4228));
hi1s1 U1014 (.Q(N4967), .DIN(N4231));
hi1s1 U1015 (.Q(N4968), .DIN(N4234));
hi1s1 U1016 (.Q(N4972), .DIN(N4246));
hi1s1 U1017 (.Q(N4973), .DIN(N4249));
hi1s1 U1018 (.Q(N4974), .DIN(N4252));
nnd2s1 U1019 (.Q(N4975), .DIN1(N4252), .DIN2(N4199));
hi1s1 U1020 (.Q(N4976), .DIN(N4206));
hi1s1 U1021 (.Q(N4977), .DIN(N4209));
and3s1 U1022 (.Q(N4978), .DIN1(N3793), .DIN2(N3789), .DIN3(N4206));
and3s1 U1023 (.Q(N4979), .DIN1(N4203), .DIN2(N4200), .DIN3(N4209));
and3s1 U1024 (.Q(N4980), .DIN1(N4097), .DIN2(N3147), .DIN3(N3158));
and3s1 U1025 (.Q(N4981), .DIN1(N4094), .DIN2(N3147), .DIN3(N3158));
and3s1 U1026 (.Q(N4982), .DIN1(N4091), .DIN2(N3147), .DIN3(N3158));
and3s1 U1027 (.Q(N4983), .DIN1(N4088), .DIN2(N3147), .DIN3(N3158));
and3s1 U1028 (.Q(N4984), .DIN1(N4153), .DIN2(N3169), .DIN3(N3180));
and3s1 U1029 (.Q(N4985), .DIN1(N4147), .DIN2(N3169), .DIN3(N3180));
and3s1 U1030 (.Q(N4986), .DIN1(N4144), .DIN2(N3169), .DIN3(N3180));
and3s1 U1031 (.Q(N4987), .DIN1(N4150), .DIN2(N3169), .DIN3(N3180));
nnd2s1 U1032 (.Q(N5049), .DIN1(N4701), .DIN2(N4702));
hi1s1 U1033 (.Q(N5052), .DIN(N4237));
hi1s1 U1034 (.Q(N5053), .DIN(N4240));
hi1s1 U1035 (.Q(N5054), .DIN(N4243));
hi1s1 U1036 (.Q(N5055), .DIN(N4255));
hi1s1 U1037 (.Q(N5056), .DIN(N4258));
nnd2s1 U1038 (.Q(N5057), .DIN1(N3819), .DIN2(N4720));
hi1s1 U1039 (.Q(N5058), .DIN(N4264));
nnd2s1 U1040 (.Q(N5059), .DIN1(N4264), .DIN2(N4267));
and4s1 U1041 (.Q(N5060), .DIN1(N4724), .DIN2(N4725), .DIN3(N4269), .DIN4(N4027));
and4s1 U1042 (.Q(N5061), .DIN1(N4726), .DIN2(N4727), .DIN3(N3827), .DIN4(N4728));
and4s1 U1043 (.Q(N5062), .DIN1(N4729), .DIN2(N4730), .DIN3(N4731), .DIN4(N4732));
and4s1 U1044 (.Q(N5063), .DIN1(N4733), .DIN2(N4734), .DIN3(N4735), .DIN4(N4736));
and2s1 U1045 (.Q(N5065), .DIN1(N4357), .DIN2(N4375));
and3s1 U1046 (.Q(N5066), .DIN1(N4364), .DIN2(N4357), .DIN3(N4379));
and2s1 U1047 (.Q(N5067), .DIN1(N4418), .DIN2(N4436));
and3s1 U1048 (.Q(N5068), .DIN1(N4425), .DIN2(N4418), .DIN3(N4440));
hi1s1 U1049 (.Q(N5069), .DIN(N4548));
nnd2s1 U1050 (.Q(N5070), .DIN1(N4548), .DIN2(N2628));
hi1s1 U1051 (.Q(N5071), .DIN(N4551));
nnd2s1 U1052 (.Q(N5072), .DIN1(N4551), .DIN2(N2629));
hi1s1 U1053 (.Q(N5073), .DIN(N4554));
nnd2s1 U1054 (.Q(N5074), .DIN1(N4554), .DIN2(N2630));
hi1s1 U1055 (.Q(N5075), .DIN(N4557));
nnd2s1 U1056 (.Q(N5076), .DIN1(N4557), .DIN2(N2631));
hi1s1 U1057 (.Q(N5077), .DIN(N4560));
nnd2s1 U1058 (.Q(N5078), .DIN1(N4560), .DIN2(N2632));
hi1s1 U1059 (.Q(N5079), .DIN(N4563));
nnd2s1 U1060 (.Q(N5080), .DIN1(N4563), .DIN2(N2633));
hi1s1 U1061 (.Q(N5081), .DIN(N4566));
nnd2s1 U1062 (.Q(N5082), .DIN1(N4566), .DIN2(N2634));
hi1s1 U1063 (.Q(N5083), .DIN(N4569));
nnd2s1 U1064 (.Q(N5084), .DIN1(N4569), .DIN2(N2635));
hi1s1 U1065 (.Q(N5085), .DIN(N4572));
nnd2s1 U1066 (.Q(N5086), .DIN1(N4572), .DIN2(N2636));
hi1s1 U1067 (.Q(N5087), .DIN(N4575));
nnd2s1 U1068 (.Q(N5088), .DIN1(N4578), .DIN2(N2638));
hi1s1 U1069 (.Q(N5089), .DIN(N4578));
nnd2s1 U1070 (.Q(N5090), .DIN1(N4581), .DIN2(N2639));
hi1s1 U1071 (.Q(N5091), .DIN(N4581));
nnd2s1 U1072 (.Q(N5092), .DIN1(N4584), .DIN2(N2640));
hi1s1 U1073 (.Q(N5093), .DIN(N4584));
nnd2s1 U1074 (.Q(N5094), .DIN1(N4587), .DIN2(N2641));
hi1s1 U1075 (.Q(N5095), .DIN(N4587));
nnd2s1 U1076 (.Q(N5096), .DIN1(N4590), .DIN2(N2642));
hi1s1 U1077 (.Q(N5097), .DIN(N4590));
nnd2s1 U1078 (.Q(N5098), .DIN1(N4593), .DIN2(N2643));
hi1s1 U1079 (.Q(N5099), .DIN(N4593));
nnd2s1 U1080 (.Q(N5100), .DIN1(N4596), .DIN2(N2644));
hi1s1 U1081 (.Q(N5101), .DIN(N4596));
nnd2s1 U1082 (.Q(N5102), .DIN1(N4599), .DIN2(N2645));
hi1s1 U1083 (.Q(N5103), .DIN(N4599));
nnd2s1 U1084 (.Q(N5104), .DIN1(N4602), .DIN2(N2646));
hi1s1 U1085 (.Q(N5105), .DIN(N4602));
hi1s1 U1086 (.Q(N5106), .DIN(N4611));
nnd2s1 U1087 (.Q(N5107), .DIN1(N4611), .DIN2(N2709));
hi1s1 U1088 (.Q(N5108), .DIN(N4614));
nnd2s1 U1089 (.Q(N5109), .DIN1(N4614), .DIN2(N2710));
hi1s1 U1090 (.Q(N5110), .DIN(N4617));
nnd2s1 U1091 (.Q(N5111), .DIN1(N4617), .DIN2(N2711));
nnd2s1 U1092 (.Q(N5112), .DIN1(N1890), .DIN2(N4855));
hi1s1 U1093 (.Q(N5113), .DIN(N4621));
nnd2s1 U1094 (.Q(N5114), .DIN1(N4621), .DIN2(N2713));
hi1s1 U1095 (.Q(N5115), .DIN(N4624));
nnd2s1 U1096 (.Q(N5116), .DIN1(N4624), .DIN2(N2714));
and2s1 U1097 (.Q(N5117), .DIN1(N4364), .DIN2(N4379));
and2s1 U1098 (.Q(N5118), .DIN1(N4364), .DIN2(N4379));
and2s1 U1099 (.Q(N5119), .DIN1(N54), .DIN2(N4405));
hi1s1 U1100 (.Q(N5120), .DIN(N4627));
nnd2s1 U1101 (.Q(N5121), .DIN1(N4630), .DIN2(N2716));
hi1s1 U1102 (.Q(N5122), .DIN(N4630));
nnd2s1 U1103 (.Q(N5123), .DIN1(N4633), .DIN2(N2717));
hi1s1 U1104 (.Q(N5124), .DIN(N4633));
nnd2s1 U1105 (.Q(N5125), .DIN1(N1908), .DIN2(N4909));
nnd2s1 U1106 (.Q(N5126), .DIN1(N4637), .DIN2(N2719));
hi1s1 U1107 (.Q(N5127), .DIN(N4637));
nnd2s1 U1108 (.Q(N5128), .DIN1(N4640), .DIN2(N2720));
hi1s1 U1109 (.Q(N5129), .DIN(N4640));
nnd2s1 U1110 (.Q(N5130), .DIN1(N4643), .DIN2(N2721));
hi1s1 U1111 (.Q(N5131), .DIN(N4643));
and2s1 U1112 (.Q(N5132), .DIN1(N4425), .DIN2(N4440));
and2s1 U1113 (.Q(N5133), .DIN1(N4425), .DIN2(N4440));
hi1s1 U1114 (.Q(N5135), .DIN(N4649));
hi1s1 U1115 (.Q(N5136), .DIN(N4652));
nnd2s1 U1116 (.Q(N5137), .DIN1(N4655), .DIN2(N4521));
hi1s1 U1117 (.Q(N5138), .DIN(N4655));
hi1s1 U1118 (.Q(N5139), .DIN(N4658));
nnd2s1 U1119 (.Q(N5140), .DIN1(N4658), .DIN2(N4947));
hi1s1 U1120 (.Q(N5141), .DIN(N4674));
hi1s1 U1121 (.Q(N5142), .DIN(N4677));
hi1s1 U1122 (.Q(N5143), .DIN(N4680));
hi1s1 U1123 (.Q(N5144), .DIN(N4683));
nnd2s1 U1124 (.Q(N5145), .DIN1(N4686), .DIN2(N4523));
hi1s1 U1125 (.Q(N5146), .DIN(N4686));
nor2s1 U1126 (.Q(N5147), .DIN1(N4953), .DIN2(N4196));
nor2s1 U1127 (.Q(N5148), .DIN1(N4954), .DIN2(N4955));
hi1s1 U1128 (.Q(N5150), .DIN(N4524));
nnd2s1 U1129 (.Q(N5153), .DIN1(N4228), .DIN2(N4965));
nnd2s1 U1130 (.Q(N5154), .DIN1(N4225), .DIN2(N4966));
nnd2s1 U1131 (.Q(N5155), .DIN1(N4234), .DIN2(N4967));
nnd2s1 U1132 (.Q(N5156), .DIN1(N4231), .DIN2(N4968));
hi1s1 U1133 (.Q(N5157), .DIN(N4532));
nnd2s1 U1134 (.Q(N5160), .DIN1(N4249), .DIN2(N4972));
nnd2s1 U1135 (.Q(N5161), .DIN1(N4246), .DIN2(N4973));
nnd2s1 U1136 (.Q(N5162), .DIN1(N3816), .DIN2(N4974));
and3s1 U1137 (.Q(N5163), .DIN1(N4200), .DIN2(N3793), .DIN3(N4976));
and3s1 U1138 (.Q(N5164), .DIN1(N3789), .DIN2(N4203), .DIN3(N4977));
and3s1 U1139 (.Q(N5165), .DIN1(N4942), .DIN2(N3147), .DIN3(N3158));
hi1s1 U1140 (.Q(N5166), .DIN(N4512));
nb1s1 U1141 (.Q(N5169), .DIN(N4290));
hi1s1 U1142 (.Q(N5172), .DIN(N4605));
nb1s1 U1143 (.Q(N5173), .DIN(N4325));
hi1s1 U1144 (.Q(N5176), .DIN(N4608));
nb1s1 U1145 (.Q(N5177), .DIN(N4349));
nb1s1 U1146 (.Q(N5180), .DIN(N4405));
nb1s1 U1147 (.Q(N5183), .DIN(N4357));
nb1s1 U1148 (.Q(N5186), .DIN(N4357));
nb1s1 U1149 (.Q(N5189), .DIN(N4364));
nb1s1 U1150 (.Q(N5192), .DIN(N4364));
nb1s1 U1151 (.Q(N5195), .DIN(N4385));
hi1s1 U1152 (.Q(N5198), .DIN(N4646));
nb1s1 U1153 (.Q(N5199), .DIN(N4418));
nb1s1 U1154 (.Q(N5202), .DIN(N4425));
nb1s1 U1155 (.Q(N5205), .DIN(N4445));
nb1s1 U1156 (.Q(N5208), .DIN(N4418));
nb1s1 U1157 (.Q(N5211), .DIN(N4425));
nb1s1 U1158 (.Q(N5214), .DIN(N4477));
nb1s1 U1159 (.Q(N5217), .DIN(N4469));
nb1s1 U1160 (.Q(N5220), .DIN(N4477));
hi1s1 U1161 (.Q(N5223), .DIN(N4662));
hi1s1 U1162 (.Q(N5224), .DIN(N4665));
hi1s1 U1163 (.Q(N5225), .DIN(N4668));
hi1s1 U1164 (.Q(N5226), .DIN(N4671));
hi1s1 U1165 (.Q(N5227), .DIN(N4689));
hi1s1 U1166 (.Q(N5228), .DIN(N4692));
hi1s1 U1167 (.Q(N5229), .DIN(N4695));
hi1s1 U1168 (.Q(N5230), .DIN(N4698));
nnd2s1 U1169 (.Q(N5232), .DIN1(N4240), .DIN2(N5052));
nnd2s1 U1170 (.Q(N5233), .DIN1(N4237), .DIN2(N5053));
nnd2s1 U1171 (.Q(N5234), .DIN1(N4258), .DIN2(N5055));
nnd2s1 U1172 (.Q(N5235), .DIN1(N4255), .DIN2(N5056));
nnd2s1 U1173 (.Q(N5236), .DIN1(N4721), .DIN2(N5057));
nnd2s1 U1174 (.Q(N5239), .DIN1(N3824), .DIN2(N5058));
and3s1 U1175 (.Q(N5240), .DIN1(N5060), .DIN2(N5061), .DIN3(N4270));
hi1s1 U1176 (.Q(N5241), .DIN(N4939));
nnd2s1 U1177 (.Q(N5242), .DIN1(N1824), .DIN2(N5069));
nnd2s1 U1178 (.Q(N5243), .DIN1(N1827), .DIN2(N5071));
nnd2s1 U1179 (.Q(N5244), .DIN1(N1830), .DIN2(N5073));
nnd2s1 U1180 (.Q(N5245), .DIN1(N1833), .DIN2(N5075));
nnd2s1 U1181 (.Q(N5246), .DIN1(N1836), .DIN2(N5077));
nnd2s1 U1182 (.Q(N5247), .DIN1(N1839), .DIN2(N5079));
nnd2s1 U1183 (.Q(N5248), .DIN1(N1842), .DIN2(N5081));
nnd2s1 U1184 (.Q(N5249), .DIN1(N1845), .DIN2(N5083));
nnd2s1 U1185 (.Q(N5250), .DIN1(N1848), .DIN2(N5085));
nnd2s1 U1186 (.Q(N5252), .DIN1(N1854), .DIN2(N5089));
nnd2s1 U1187 (.Q(N5253), .DIN1(N1857), .DIN2(N5091));
nnd2s1 U1188 (.Q(N5254), .DIN1(N1860), .DIN2(N5093));
nnd2s1 U1189 (.Q(N5255), .DIN1(N1863), .DIN2(N5095));
nnd2s1 U1190 (.Q(N5256), .DIN1(N1866), .DIN2(N5097));
nnd2s1 U1191 (.Q(N5257), .DIN1(N1869), .DIN2(N5099));
nnd2s1 U1192 (.Q(N5258), .DIN1(N1872), .DIN2(N5101));
nnd2s1 U1193 (.Q(N5259), .DIN1(N1875), .DIN2(N5103));
nnd2s1 U1194 (.Q(N5260), .DIN1(N1878), .DIN2(N5105));
nnd2s1 U1195 (.Q(N5261), .DIN1(N1881), .DIN2(N5106));
nnd2s1 U1196 (.Q(N5262), .DIN1(N1884), .DIN2(N5108));
nnd2s1 U1197 (.Q(N5263), .DIN1(N1887), .DIN2(N5110));
nnd2s1 U1198 (.Q(N5264), .DIN1(N5112), .DIN2(N4856));
nnd2s1 U1199 (.Q(N5274), .DIN1(N1893), .DIN2(N5113));
nnd2s1 U1200 (.Q(N5275), .DIN1(N1896), .DIN2(N5115));
nnd2s1 U1201 (.Q(N5282), .DIN1(N1902), .DIN2(N5122));
nnd2s1 U1202 (.Q(N5283), .DIN1(N1905), .DIN2(N5124));
nnd2s1 U1203 (.Q(N5284), .DIN1(N4908), .DIN2(N5125));
nnd2s1 U1204 (.Q(N5298), .DIN1(N1911), .DIN2(N5127));
nnd2s1 U1205 (.Q(N5299), .DIN1(N1914), .DIN2(N5129));
nnd2s1 U1206 (.Q(N5300), .DIN1(N1917), .DIN2(N5131));
nnd2s1 U1207 (.Q(N5303), .DIN1(N4652), .DIN2(N5135));
nnd2s1 U1208 (.Q(N5304), .DIN1(N4649), .DIN2(N5136));
nnd2s1 U1209 (.Q(N5305), .DIN1(N4008), .DIN2(N5138));
nnd2s1 U1210 (.Q(N5306), .DIN1(N4219), .DIN2(N5139));
nnd2s1 U1211 (.Q(N5307), .DIN1(N4677), .DIN2(N5141));
nnd2s1 U1212 (.Q(N5308), .DIN1(N4674), .DIN2(N5142));
nnd2s1 U1213 (.Q(N5309), .DIN1(N4683), .DIN2(N5143));
nnd2s1 U1214 (.Q(N5310), .DIN1(N4680), .DIN2(N5144));
nnd2s1 U1215 (.Q(N5311), .DIN1(N4011), .DIN2(N5146));
hi1s1 U1216 (.Q(N5312), .DIN(N5049));
nnd2s1 U1217 (.Q(N5315), .DIN1(N5153), .DIN2(N5154));
nnd2s1 U1218 (.Q(N5319), .DIN1(N5155), .DIN2(N5156));
nnd2s1 U1219 (.Q(N5324), .DIN1(N5160), .DIN2(N5161));
nnd2s1 U1220 (.Q(N5328), .DIN1(N5162), .DIN2(N4975));
nor2s1 U1221 (.Q(N5331), .DIN1(N5163), .DIN2(N4978));
nor2s1 U1222 (.Q(N5332), .DIN1(N5164), .DIN2(N4979));
or2s1 U1223 (.Q(N5346), .DIN1(N4412), .DIN2(N5119));
nnd2s1 U1224 (.Q(N5363), .DIN1(N4665), .DIN2(N5223));
nnd2s1 U1225 (.Q(N5364), .DIN1(N4662), .DIN2(N5224));
nnd2s1 U1226 (.Q(N5365), .DIN1(N4671), .DIN2(N5225));
nnd2s1 U1227 (.Q(N5366), .DIN1(N4668), .DIN2(N5226));
nnd2s1 U1228 (.Q(N5367), .DIN1(N4692), .DIN2(N5227));
nnd2s1 U1229 (.Q(N5368), .DIN1(N4689), .DIN2(N5228));
nnd2s1 U1230 (.Q(N5369), .DIN1(N4698), .DIN2(N5229));
nnd2s1 U1231 (.Q(N5370), .DIN1(N4695), .DIN2(N5230));
nnd2s1 U1232 (.Q(N5371), .DIN1(N5148), .DIN2(N5147));
nb1s1 U1233 (.Q(N5374), .DIN(N4939));
nnd2s1 U1234 (.Q(N5377), .DIN1(N5232), .DIN2(N5233));
nnd2s1 U1235 (.Q(N5382), .DIN1(N5234), .DIN2(N5235));
nnd2s1 U1236 (.Q(N5385), .DIN1(N5239), .DIN2(N5059));
and3s1 U1237 (.Q(N5388), .DIN1(N5062), .DIN2(N5063), .DIN3(N5241));
nnd2s1 U1238 (.Q(N5389), .DIN1(N5242), .DIN2(N5070));
nnd2s1 U1239 (.Q(N5396), .DIN1(N5243), .DIN2(N5072));
nnd2s1 U1240 (.Q(N5407), .DIN1(N5244), .DIN2(N5074));
nnd2s1 U1241 (.Q(N5418), .DIN1(N5245), .DIN2(N5076));
nnd2s1 U1242 (.Q(N5424), .DIN1(N5246), .DIN2(N5078));
nnd2s1 U1243 (.Q(N5431), .DIN1(N5247), .DIN2(N5080));
nnd2s1 U1244 (.Q(N5441), .DIN1(N5248), .DIN2(N5082));
nnd2s1 U1245 (.Q(N5452), .DIN1(N5249), .DIN2(N5084));
nnd2s1 U1246 (.Q(N5462), .DIN1(N5250), .DIN2(N5086));
hi1s1 U1247 (.Q(N5469), .DIN(N5169));
nnd2s1 U1248 (.Q(N5470), .DIN1(N5088), .DIN2(N5252));
nnd2s1 U1249 (.Q(N5477), .DIN1(N5090), .DIN2(N5253));
nnd2s1 U1250 (.Q(N5488), .DIN1(N5092), .DIN2(N5254));
nnd2s1 U1251 (.Q(N5498), .DIN1(N5094), .DIN2(N5255));
nnd2s1 U1252 (.Q(N5506), .DIN1(N5096), .DIN2(N5256));
nnd2s1 U1253 (.Q(N5520), .DIN1(N5098), .DIN2(N5257));
nnd2s1 U1254 (.Q(N5536), .DIN1(N5100), .DIN2(N5258));
nnd2s1 U1255 (.Q(N5549), .DIN1(N5102), .DIN2(N5259));
nnd2s1 U1256 (.Q(N5555), .DIN1(N5104), .DIN2(N5260));
nnd2s1 U1257 (.Q(N5562), .DIN1(N5261), .DIN2(N5107));
nnd2s1 U1258 (.Q(N5573), .DIN1(N5262), .DIN2(N5109));
nnd2s1 U1259 (.Q(N5579), .DIN1(N5263), .DIN2(N5111));
nnd2s1 U1260 (.Q(N5595), .DIN1(N5274), .DIN2(N5114));
nnd2s1 U1261 (.Q(N5606), .DIN1(N5275), .DIN2(N5116));
nnd2s1 U1262 (.Q(N5616), .DIN1(N5180), .DIN2(N2715));
hi1s1 U1263 (.Q(N5617), .DIN(N5180));
hi1s1 U1264 (.Q(N5618), .DIN(N5183));
hi1s1 U1265 (.Q(N5619), .DIN(N5186));
hi1s1 U1266 (.Q(N5620), .DIN(N5189));
hi1s1 U1267 (.Q(N5621), .DIN(N5192));
hi1s1 U1268 (.Q(N5622), .DIN(N5195));
nnd2s1 U1269 (.Q(N5624), .DIN1(N5121), .DIN2(N5282));
nnd2s1 U1270 (.Q(N5634), .DIN1(N5123), .DIN2(N5283));
nnd2s1 U1271 (.Q(N5655), .DIN1(N5126), .DIN2(N5298));
nnd2s1 U1272 (.Q(N5671), .DIN1(N5128), .DIN2(N5299));
nnd2s1 U1273 (.Q(N5684), .DIN1(N5130), .DIN2(N5300));
hi1s1 U1274 (.Q(N5690), .DIN(N5202));
hi1s1 U1275 (.Q(N5691), .DIN(N5211));
nnd2s1 U1276 (.Q(N5692), .DIN1(N5303), .DIN2(N5304));
nnd2s1 U1277 (.Q(N5696), .DIN1(N5137), .DIN2(N5305));
nnd2s1 U1278 (.Q(N5700), .DIN1(N5306), .DIN2(N5140));
nnd2s1 U1279 (.Q(N5703), .DIN1(N5307), .DIN2(N5308));
nnd2s1 U1280 (.Q(N5707), .DIN1(N5309), .DIN2(N5310));
nnd2s1 U1281 (.Q(N5711), .DIN1(N5145), .DIN2(N5311));
and2s1 U1282 (.Q(N5726), .DIN1(N5166), .DIN2(N4512));
hi1s1 U1283 (.Q(N5727), .DIN(N5173));
hi1s1 U1284 (.Q(N5728), .DIN(N5177));
hi1s1 U1285 (.Q(N5730), .DIN(N5199));
hi1s1 U1286 (.Q(N5731), .DIN(N5205));
hi1s1 U1287 (.Q(N5732), .DIN(N5208));
hi1s1 U1288 (.Q(N5733), .DIN(N5214));
hi1s1 U1289 (.Q(N5734), .DIN(N5217));
hi1s1 U1290 (.Q(N5735), .DIN(N5220));
nnd2s1 U1291 (.Q(N5736), .DIN1(N5365), .DIN2(N5366));
nnd2s1 U1292 (.Q(N5739), .DIN1(N5363), .DIN2(N5364));
nnd2s1 U1293 (.Q(N5742), .DIN1(N5369), .DIN2(N5370));
nnd2s1 U1294 (.Q(N5745), .DIN1(N5367), .DIN2(N5368));
hi1s1 U1295 (.Q(N5755), .DIN(N5236));
nnd2s1 U1296 (.Q(N5756), .DIN1(N5332), .DIN2(N5331));
and2s1 U1297 (.Q(N5954), .DIN1(N5264), .DIN2(N4396));
nnd2s1 U1298 (.Q(N5955), .DIN1(N1899), .DIN2(N5617));
hi1s1 U1299 (.Q(N5956), .DIN(N5346));
and2s1 U1300 (.Q(N6005), .DIN1(N5284), .DIN2(N4456));
and2s1 U1301 (.Q(N6006), .DIN1(N5284), .DIN2(N4456));
hi1s1 U1302 (.Q(N6023), .DIN(N5371));
nnd2s1 U1303 (.Q(N6024), .DIN1(N5371), .DIN2(N5312));
hi1s1 U1304 (.Q(N6025), .DIN(N5315));
hi1s1 U1305 (.Q(N6028), .DIN(N5324));
nb1s1 U1306 (.Q(N6031), .DIN(N5319));
nb1s1 U1307 (.Q(N6034), .DIN(N5319));
nb1s1 U1308 (.Q(N6037), .DIN(N5328));
nb1s1 U1309 (.Q(N6040), .DIN(N5328));
hi1s1 U1310 (.Q(N6044), .DIN(N5385));
or2s1 U1311 (.Q(N6045), .DIN1(N5166), .DIN2(N5726));
nb1s1 U1312 (.Q(N6048), .DIN(N5264));
nb1s1 U1313 (.Q(N6051), .DIN(N5284));
nb1s1 U1314 (.Q(N6054), .DIN(N5284));
hi1s1 U1315 (.Q(N6065), .DIN(N5374));
nnd2s1 U1316 (.Q(N6066), .DIN1(N5374), .DIN2(N5054));
hi1s1 U1317 (.Q(N6067), .DIN(N5377));
hi1s1 U1318 (.Q(N6068), .DIN(N5382));
nnd2s1 U1319 (.Q(N6069), .DIN1(N5382), .DIN2(N5755));
and2s1 U1320 (.Q(N6071), .DIN1(N5470), .DIN2(N4316));
and3s1 U1321 (.Q(N6072), .DIN1(N5477), .DIN2(N5470), .DIN3(N4320));
and4s1 U1322 (.Q(N6073), .DIN1(N5488), .DIN2(N5470), .DIN3(N4325), .DIN4(N5477));
and4s1 U1323 (.Q(N6074), .DIN1(N5562), .DIN2(N4357), .DIN3(N4385), .DIN4(N4364));
and2s1 U1324 (.Q(N6075), .DIN1(N5389), .DIN2(N4280));
and3s1 U1325 (.Q(N6076), .DIN1(N5396), .DIN2(N5389), .DIN3(N4284));
and4s1 U1326 (.Q(N6077), .DIN1(N5407), .DIN2(N5389), .DIN3(N4290), .DIN4(N5396));
and4s1 U1327 (.Q(N6078), .DIN1(N5624), .DIN2(N4418), .DIN3(N4445), .DIN4(N4425));
hi1s1 U1328 (.Q(N6079), .DIN(N5418));
and4s1 U1329 (.Q(N6080), .DIN1(N5396), .DIN2(N5418), .DIN3(N5407), .DIN4(N5389));
and2s1 U1330 (.Q(N6083), .DIN1(N5396), .DIN2(N4284));
and3s1 U1331 (.Q(N6084), .DIN1(N5407), .DIN2(N4290), .DIN3(N5396));
and3s1 U1332 (.Q(N6085), .DIN1(N5418), .DIN2(N5407), .DIN3(N5396));
and2s1 U1333 (.Q(N6086), .DIN1(N5396), .DIN2(N4284));
and3s1 U1334 (.Q(N6087), .DIN1(N4290), .DIN2(N5407), .DIN3(N5396));
and2s1 U1335 (.Q(N6088), .DIN1(N5407), .DIN2(N4290));
and2s1 U1336 (.Q(N6089), .DIN1(N5418), .DIN2(N5407));
and2s1 U1337 (.Q(N6090), .DIN1(N5407), .DIN2(N4290));
and5s1 U1338 (.Q(N6091), .DIN1(N5431), .DIN2(N5462), .DIN3(N5441), .DIN4(N5424), .DIN5(N5452));
and2s1 U1339 (.Q(N6094), .DIN1(N5424), .DIN2(N4298));
and3s1 U1340 (.Q(N6095), .DIN1(N5431), .DIN2(N5424), .DIN3(N4301));
and4s1 U1341 (.Q(N6096), .DIN1(N5441), .DIN2(N5424), .DIN3(N4305), .DIN4(N5431));
and5s1 U1342 (.Q(N6097), .DIN1(N5452), .DIN2(N5441), .DIN3(N5424), .DIN4(N4310), .DIN5(N5431));
and2s1 U1343 (.Q(N6098), .DIN1(N5431), .DIN2(N4301));
and3s1 U1344 (.Q(N6099), .DIN1(N5441), .DIN2(N4305), .DIN3(N5431));
and4s1 U1345 (.Q(N6100), .DIN1(N5452), .DIN2(N5441), .DIN3(N4310), .DIN4(N5431));
and5s1 U1346 (.Q(N6101), .DIN1(N4), .DIN2(N5462), .DIN3(N5441), .DIN4(N5452), .DIN5(N5431));
and2s1 U1347 (.Q(N6102), .DIN1(N4305), .DIN2(N5441));
and3s1 U1348 (.Q(N6103), .DIN1(N5452), .DIN2(N5441), .DIN3(N4310));
and4s1 U1349 (.Q(N6104), .DIN1(N4), .DIN2(N5462), .DIN3(N5441), .DIN4(N5452));
and2s1 U1350 (.Q(N6105), .DIN1(N5452), .DIN2(N4310));
and3s1 U1351 (.Q(N6106), .DIN1(N4), .DIN2(N5462), .DIN3(N5452));
and2s1 U1352 (.Q(N6107), .DIN1(N4), .DIN2(N5462));
and4s1 U1353 (.Q(N6108), .DIN1(N5549), .DIN2(N5488), .DIN3(N5477), .DIN4(N5470));
and2s1 U1354 (.Q(N6111), .DIN1(N5477), .DIN2(N4320));
and3s1 U1355 (.Q(N6112), .DIN1(N5488), .DIN2(N4325), .DIN3(N5477));
and3s1 U1356 (.Q(N6113), .DIN1(N5549), .DIN2(N5488), .DIN3(N5477));
and2s1 U1357 (.Q(N6114), .DIN1(N5477), .DIN2(N4320));
and3s1 U1358 (.Q(N6115), .DIN1(N5488), .DIN2(N4325), .DIN3(N5477));
and2s1 U1359 (.Q(N6116), .DIN1(N5488), .DIN2(N4325));
and5s1 U1360 (.Q(N6117), .DIN1(N5555), .DIN2(N5536), .DIN3(N5520), .DIN4(N5506), .DIN5(N5498));
and2s1 U1361 (.Q(N6120), .DIN1(N5498), .DIN2(N4332));
and3s1 U1362 (.Q(N6121), .DIN1(N5506), .DIN2(N5498), .DIN3(N4336));
and4s1 U1363 (.Q(N6122), .DIN1(N5520), .DIN2(N5498), .DIN3(N4342), .DIN4(N5506));
and5s1 U1364 (.Q(N6123), .DIN1(N5536), .DIN2(N5520), .DIN3(N5498), .DIN4(N4349), .DIN5(N5506));
and2s1 U1365 (.Q(N6124), .DIN1(N5506), .DIN2(N4336));
and3s1 U1366 (.Q(N6125), .DIN1(N5520), .DIN2(N4342), .DIN3(N5506));
and4s1 U1367 (.Q(N6126), .DIN1(N5536), .DIN2(N5520), .DIN3(N4349), .DIN4(N5506));
and4s1 U1368 (.Q(N6127), .DIN1(N5555), .DIN2(N5520), .DIN3(N5506), .DIN4(N5536));
and2s1 U1369 (.Q(N6128), .DIN1(N5506), .DIN2(N4336));
and3s1 U1370 (.Q(N6129), .DIN1(N5520), .DIN2(N4342), .DIN3(N5506));
and4s1 U1371 (.Q(N6130), .DIN1(N5536), .DIN2(N5520), .DIN3(N4349), .DIN4(N5506));
and2s1 U1372 (.Q(N6131), .DIN1(N5520), .DIN2(N4342));
and3s1 U1373 (.Q(N6132), .DIN1(N5536), .DIN2(N5520), .DIN3(N4349));
and3s1 U1374 (.Q(N6133), .DIN1(N5555), .DIN2(N5520), .DIN3(N5536));
and2s1 U1375 (.Q(N6134), .DIN1(N5520), .DIN2(N4342));
and3s1 U1376 (.Q(N6135), .DIN1(N5536), .DIN2(N5520), .DIN3(N4349));
and2s1 U1377 (.Q(N6136), .DIN1(N5536), .DIN2(N4349));
and2s1 U1378 (.Q(N6137), .DIN1(N5549), .DIN2(N5488));
and2s1 U1379 (.Q(N6138), .DIN1(N5555), .DIN2(N5536));
hi1s1 U1380 (.Q(N6139), .DIN(N5573));
and4s1 U1381 (.Q(N6140), .DIN1(N4364), .DIN2(N5573), .DIN3(N5562), .DIN4(N4357));
and3s1 U1382 (.Q(N6143), .DIN1(N5562), .DIN2(N4385), .DIN3(N4364));
and3s1 U1383 (.Q(N6144), .DIN1(N5573), .DIN2(N5562), .DIN3(N4364));
and3s1 U1384 (.Q(N6145), .DIN1(N4385), .DIN2(N5562), .DIN3(N4364));
and2s1 U1385 (.Q(N6146), .DIN1(N5562), .DIN2(N4385));
and2s1 U1386 (.Q(N6147), .DIN1(N5573), .DIN2(N5562));
and2s1 U1387 (.Q(N6148), .DIN1(N5562), .DIN2(N4385));
and5s1 U1388 (.Q(N6149), .DIN1(N5264), .DIN2(N4405), .DIN3(N5595), .DIN4(N5579), .DIN5(N5606));
and2s1 U1389 (.Q(N6152), .DIN1(N5579), .DIN2(N4067));
and3s1 U1390 (.Q(N6153), .DIN1(N5264), .DIN2(N5579), .DIN3(N4396));
and4s1 U1391 (.Q(N6154), .DIN1(N5595), .DIN2(N5579), .DIN3(N4400), .DIN4(N5264));
and5s1 U1392 (.Q(N6155), .DIN1(N5606), .DIN2(N5595), .DIN3(N5579), .DIN4(N4412), .DIN5(N5264));
and3s1 U1393 (.Q(N6156), .DIN1(N5595), .DIN2(N4400), .DIN3(N5264));
and4s1 U1394 (.Q(N6157), .DIN1(N5606), .DIN2(N5595), .DIN3(N4412), .DIN4(N5264));
and5s1 U1395 (.Q(N6158), .DIN1(N54), .DIN2(N4405), .DIN3(N5595), .DIN4(N5606), .DIN5(N5264));
and2s1 U1396 (.Q(N6159), .DIN1(N4400), .DIN2(N5595));
and3s1 U1397 (.Q(N6160), .DIN1(N5606), .DIN2(N5595), .DIN3(N4412));
and4s1 U1398 (.Q(N6161), .DIN1(N54), .DIN2(N4405), .DIN3(N5595), .DIN4(N5606));
and2s1 U1399 (.Q(N6162), .DIN1(N5606), .DIN2(N4412));
and3s1 U1400 (.Q(N6163), .DIN1(N54), .DIN2(N4405), .DIN3(N5606));
nnd2s1 U1401 (.Q(N6164), .DIN1(N5616), .DIN2(N5955));
and4s1 U1402 (.Q(N6168), .DIN1(N5684), .DIN2(N5624), .DIN3(N4425), .DIN4(N4418));
and3s1 U1403 (.Q(N6171), .DIN1(N5624), .DIN2(N4445), .DIN3(N4425));
and3s1 U1404 (.Q(N6172), .DIN1(N5684), .DIN2(N5624), .DIN3(N4425));
and3s1 U1405 (.Q(N6173), .DIN1(N5624), .DIN2(N4445), .DIN3(N4425));
and2s1 U1406 (.Q(N6174), .DIN1(N5624), .DIN2(N4445));
and5s1 U1407 (.Q(N6175), .DIN1(N4477), .DIN2(N5671), .DIN3(N5655), .DIN4(N5284), .DIN5(N5634));
and2s1 U1408 (.Q(N6178), .DIN1(N5634), .DIN2(N4080));
and3s1 U1409 (.Q(N6179), .DIN1(N5284), .DIN2(N5634), .DIN3(N4456));
and4s1 U1410 (.Q(N6180), .DIN1(N5655), .DIN2(N5634), .DIN3(N4462), .DIN4(N5284));
and5s1 U1411 (.Q(N6181), .DIN1(N5671), .DIN2(N5655), .DIN3(N5634), .DIN4(N4469), .DIN5(N5284));
and3s1 U1412 (.Q(N6182), .DIN1(N5655), .DIN2(N4462), .DIN3(N5284));
and4s1 U1413 (.Q(N6183), .DIN1(N5671), .DIN2(N5655), .DIN3(N4469), .DIN4(N5284));
and4s1 U1414 (.Q(N6184), .DIN1(N4477), .DIN2(N5655), .DIN3(N5284), .DIN4(N5671));
and3s1 U1415 (.Q(N6185), .DIN1(N5655), .DIN2(N4462), .DIN3(N5284));
and4s1 U1416 (.Q(N6186), .DIN1(N5671), .DIN2(N5655), .DIN3(N4469), .DIN4(N5284));
and2s1 U1417 (.Q(N6187), .DIN1(N5655), .DIN2(N4462));
and3s1 U1418 (.Q(N6188), .DIN1(N5671), .DIN2(N5655), .DIN3(N4469));
and3s1 U1419 (.Q(N6189), .DIN1(N4477), .DIN2(N5655), .DIN3(N5671));
and2s1 U1420 (.Q(N6190), .DIN1(N5655), .DIN2(N4462));
and3s1 U1421 (.Q(N6191), .DIN1(N5671), .DIN2(N5655), .DIN3(N4469));
and2s1 U1422 (.Q(N6192), .DIN1(N5671), .DIN2(N4469));
and2s1 U1423 (.Q(N6193), .DIN1(N5684), .DIN2(N5624));
and2s1 U1424 (.Q(N6194), .DIN1(N4477), .DIN2(N5671));
hi1s1 U1425 (.Q(N6197), .DIN(N5692));
hi1s1 U1426 (.Q(N6200), .DIN(N5696));
hi1s1 U1427 (.Q(N6203), .DIN(N5703));
hi1s1 U1428 (.Q(N6206), .DIN(N5707));
nb1s1 U1429 (.Q(N6209), .DIN(N5700));
nb1s1 U1430 (.Q(N6212), .DIN(N5700));
nb1s1 U1431 (.Q(N6215), .DIN(N5711));
nb1s1 U1432 (.Q(N6218), .DIN(N5711));
nnd2s1 U1433 (.Q(N6221), .DIN1(N5049), .DIN2(N6023));
hi1s1 U1434 (.Q(N6234), .DIN(N5756));
nnd2s1 U1435 (.Q(N6235), .DIN1(N5756), .DIN2(N6044));
nb1s1 U1436 (.Q(N6238), .DIN(N5462));
nb1s1 U1437 (.Q(N6241), .DIN(N5389));
nb1s1 U1438 (.Q(N6244), .DIN(N5389));
nb1s1 U1439 (.Q(N6247), .DIN(N5396));
nb1s1 U1440 (.Q(N6250), .DIN(N5396));
nb1s1 U1441 (.Q(N6253), .DIN(N5407));
nb1s1 U1442 (.Q(N6256), .DIN(N5407));
nb1s1 U1443 (.Q(N6259), .DIN(N5424));
nb1s1 U1444 (.Q(N6262), .DIN(N5431));
nb1s1 U1445 (.Q(N6265), .DIN(N5441));
nb1s1 U1446 (.Q(N6268), .DIN(N5452));
nb1s1 U1447 (.Q(N6271), .DIN(N5549));
nb1s1 U1448 (.Q(N6274), .DIN(N5488));
nb1s1 U1449 (.Q(N6277), .DIN(N5470));
nb1s1 U1450 (.Q(N6280), .DIN(N5477));
nb1s1 U1451 (.Q(N6283), .DIN(N5549));
nb1s1 U1452 (.Q(N6286), .DIN(N5488));
nb1s1 U1453 (.Q(N6289), .DIN(N5470));
nb1s1 U1454 (.Q(N6292), .DIN(N5477));
nb1s1 U1455 (.Q(N6295), .DIN(N5555));
nb1s1 U1456 (.Q(N6298), .DIN(N5536));
nb1s1 U1457 (.Q(N6301), .DIN(N5498));
nb1s1 U1458 (.Q(N6304), .DIN(N5520));
nb1s1 U1459 (.Q(N6307), .DIN(N5506));
nb1s1 U1460 (.Q(N6310), .DIN(N5506));
nb1s1 U1461 (.Q(N6313), .DIN(N5555));
nb1s1 U1462 (.Q(N6316), .DIN(N5536));
nb1s1 U1463 (.Q(N6319), .DIN(N5498));
nb1s1 U1464 (.Q(N6322), .DIN(N5520));
nb1s1 U1465 (.Q(N6325), .DIN(N5562));
nb1s1 U1466 (.Q(N6328), .DIN(N5562));
nb1s1 U1467 (.Q(N6331), .DIN(N5579));
nb1s1 U1468 (.Q(N6335), .DIN(N5595));
nb1s1 U1469 (.Q(N6338), .DIN(N5606));
nb1s1 U1470 (.Q(N6341), .DIN(N5684));
nb1s1 U1471 (.Q(N6344), .DIN(N5624));
nb1s1 U1472 (.Q(N6347), .DIN(N5684));
nb1s1 U1473 (.Q(N6350), .DIN(N5624));
nb1s1 U1474 (.Q(N6353), .DIN(N5671));
nb1s1 U1475 (.Q(N6356), .DIN(N5634));
nb1s1 U1476 (.Q(N6359), .DIN(N5655));
nb1s1 U1477 (.Q(N6364), .DIN(N5671));
nb1s1 U1478 (.Q(N6367), .DIN(N5634));
nb1s1 U1479 (.Q(N6370), .DIN(N5655));
hi1s1 U1480 (.Q(N6373), .DIN(N5736));
hi1s1 U1481 (.Q(N6374), .DIN(N5739));
hi1s1 U1482 (.Q(N6375), .DIN(N5742));
hi1s1 U1483 (.Q(N6376), .DIN(N5745));
nnd2s1 U1484 (.Q(N6377), .DIN1(N4243), .DIN2(N6065));
nnd2s1 U1485 (.Q(N6378), .DIN1(N5236), .DIN2(N6068));
or4s1 U1486 (.Q(N6382), .DIN1(N4268), .DIN2(N6071), .DIN3(N6072), .DIN4(N6073));
or4s1 U1487 (.Q(N6386), .DIN1(N3968), .DIN2(N5065), .DIN3(N5066), .DIN4(N6074));
or4s1 U1488 (.Q(N6388), .DIN1(N4271), .DIN2(N6075), .DIN3(N6076), .DIN4(N6077));
or4s1 U1489 (.Q(N6392), .DIN1(N3968), .DIN2(N5067), .DIN3(N5068), .DIN4(N6078));
or5s1 U1490 (.Q(N6397), .DIN1(N4297), .DIN2(N6094), .DIN3(N6095), .DIN4(N6096), .DIN5(N6097));
or2s1 U1491 (.Q(N6411), .DIN1(N4320), .DIN2(N6116));
or5s1 U1492 (.Q(N6415), .DIN1(N4331), .DIN2(N6120), .DIN3(N6121), .DIN4(N6122), .DIN5(N6123));
or2s1 U1493 (.Q(N6419), .DIN1(N4342), .DIN2(N6136));
or5s1 U1494 (.Q(N6427), .DIN1(N4392), .DIN2(N6152), .DIN3(N6153), .DIN4(N6154), .DIN5(N6155));
hi1s1 U1495 (.Q(N6434), .DIN(N6048));
or2s1 U1496 (.Q(N6437), .DIN1(N4440), .DIN2(N6174));
or5s1 U1497 (.Q(N6441), .DIN1(N4451), .DIN2(N6178), .DIN3(N6179), .DIN4(N6180), .DIN5(N6181));
or2s1 U1498 (.Q(N6445), .DIN1(N4462), .DIN2(N6192));
hi1s1 U1499 (.Q(N6448), .DIN(N6051));
hi1s1 U1500 (.Q(N6449), .DIN(N6054));
nnd2s1 U1501 (.Q(N6466), .DIN1(N6221), .DIN2(N6024));
hi1s1 U1502 (.Q(N6469), .DIN(N6031));
hi1s1 U1503 (.Q(N6470), .DIN(N6034));
hi1s1 U1504 (.Q(N6471), .DIN(N6037));
hi1s1 U1505 (.Q(N6472), .DIN(N6040));
and3s1 U1506 (.Q(N6473), .DIN1(N5315), .DIN2(N4524), .DIN3(N6031));
and3s1 U1507 (.Q(N6474), .DIN1(N6025), .DIN2(N5150), .DIN3(N6034));
and3s1 U1508 (.Q(N6475), .DIN1(N5324), .DIN2(N4532), .DIN3(N6037));
and3s1 U1509 (.Q(N6476), .DIN1(N6028), .DIN2(N5157), .DIN3(N6040));
nnd2s1 U1510 (.Q(N6477), .DIN1(N5385), .DIN2(N6234));
nnd2s1 U1511 (.Q(N6478), .DIN1(N6045), .DIN2(N132));
or4s1 U1512 (.Q(N6482), .DIN1(N4280), .DIN2(N6083), .DIN3(N6084), .DIN4(N6085));
nor3s1 U1513 (.Q(N6486), .DIN1(N4280), .DIN2(N6086), .DIN3(N6087));
or3s1 U1514 (.Q(N6490), .DIN1(N4284), .DIN2(N6088), .DIN3(N6089));
nor2s1 U1515 (.Q(N6494), .DIN1(N4284), .DIN2(N6090));
or5s1 U1516 (.Q(N6500), .DIN1(N4298), .DIN2(N6098), .DIN3(N6099), .DIN4(N6100), .DIN5(N6101));
or4s1 U1517 (.Q(N6504), .DIN1(N4301), .DIN2(N6102), .DIN3(N6103), .DIN4(N6104));
or3s1 U1518 (.Q(N6508), .DIN1(N4305), .DIN2(N6105), .DIN3(N6106));
or2s1 U1519 (.Q(N6512), .DIN1(N4310), .DIN2(N6107));
or4s1 U1520 (.Q(N6516), .DIN1(N4316), .DIN2(N6111), .DIN3(N6112), .DIN4(N6113));
nor3s1 U1521 (.Q(N6526), .DIN1(N4316), .DIN2(N6114), .DIN3(N6115));
or4s1 U1522 (.Q(N6536), .DIN1(N4336), .DIN2(N6131), .DIN3(N6132), .DIN4(N6133));
or5s1 U1523 (.Q(N6539), .DIN1(N4332), .DIN2(N6124), .DIN3(N6125), .DIN4(N6126), .DIN5(N6127));
nor3s1 U1524 (.Q(N6553), .DIN1(N4336), .DIN2(N6134), .DIN3(N6135));
nor4s1 U1525 (.Q(N6556), .DIN1(N4332), .DIN2(N6128), .DIN3(N6129), .DIN4(N6130));
or4s1 U1526 (.Q(N6566), .DIN1(N4375), .DIN2(N5117), .DIN3(N6143), .DIN4(N6144));
nor3s1 U1527 (.Q(N6569), .DIN1(N4375), .DIN2(N5118), .DIN3(N6145));
or3s1 U1528 (.Q(N6572), .DIN1(N4379), .DIN2(N6146), .DIN3(N6147));
nor2s1 U1529 (.Q(N6575), .DIN1(N4379), .DIN2(N6148));
or5s1 U1530 (.Q(N6580), .DIN1(N4067), .DIN2(N5954), .DIN3(N6156), .DIN4(N6157), .DIN5(N6158));
or4s1 U1531 (.Q(N6584), .DIN1(N4396), .DIN2(N6159), .DIN3(N6160), .DIN4(N6161));
or3s1 U1532 (.Q(N6587), .DIN1(N4400), .DIN2(N6162), .DIN3(N6163));
or4s1 U1533 (.Q(N6592), .DIN1(N4436), .DIN2(N5132), .DIN3(N6171), .DIN4(N6172));
nor3s1 U1534 (.Q(N6599), .DIN1(N4436), .DIN2(N5133), .DIN3(N6173));
or4s1 U1535 (.Q(N6606), .DIN1(N4456), .DIN2(N6187), .DIN3(N6188), .DIN4(N6189));
or5s1 U1536 (.Q(N6609), .DIN1(N4080), .DIN2(N6005), .DIN3(N6182), .DIN4(N6183), .DIN5(N6184));
nor3s1 U1537 (.Q(N6619), .DIN1(N4456), .DIN2(N6190), .DIN3(N6191));
nor4s1 U1538 (.Q(N6622), .DIN1(N4080), .DIN2(N6006), .DIN3(N6185), .DIN4(N6186));
nnd2s1 U1539 (.Q(N6630), .DIN1(N5739), .DIN2(N6373));
nnd2s1 U1540 (.Q(N6631), .DIN1(N5736), .DIN2(N6374));
nnd2s1 U1541 (.Q(N6632), .DIN1(N5745), .DIN2(N6375));
nnd2s1 U1542 (.Q(N6633), .DIN1(N5742), .DIN2(N6376));
nnd2s1 U1543 (.Q(N6634), .DIN1(N6377), .DIN2(N6066));
nnd2s1 U1544 (.Q(N6637), .DIN1(N6069), .DIN2(N6378));
hi1s1 U1545 (.Q(N6640), .DIN(N6164));
and2s1 U1546 (.Q(N6641), .DIN1(N6108), .DIN2(N6117));
and2s1 U1547 (.Q(N6643), .DIN1(N6140), .DIN2(N6149));
and2s1 U1548 (.Q(N6646), .DIN1(N6168), .DIN2(N6175));
and2s1 U1549 (.Q(N6648), .DIN1(N6080), .DIN2(N6091));
nnd2s1 U1550 (.Q(N6650), .DIN1(N6238), .DIN2(N2637));
hi1s1 U1551 (.Q(N6651), .DIN(N6238));
hi1s1 U1552 (.Q(N6653), .DIN(N6241));
hi1s1 U1553 (.Q(N6655), .DIN(N6244));
hi1s1 U1554 (.Q(N6657), .DIN(N6247));
hi1s1 U1555 (.Q(N6659), .DIN(N6250));
nnd2s1 U1556 (.Q(N6660), .DIN1(N6253), .DIN2(N5087));
hi1s1 U1557 (.Q(N6661), .DIN(N6253));
nnd2s1 U1558 (.Q(N6662), .DIN1(N6256), .DIN2(N5469));
hi1s1 U1559 (.Q(N6663), .DIN(N6256));
and2s1 U1560 (.Q(N6664), .DIN1(N6091), .DIN2(N4));
hi1s1 U1561 (.Q(N6666), .DIN(N6259));
hi1s1 U1562 (.Q(N6668), .DIN(N6262));
hi1s1 U1563 (.Q(N6670), .DIN(N6265));
hi1s1 U1564 (.Q(N6672), .DIN(N6268));
hi1s1 U1565 (.Q(N6675), .DIN(N6117));
hi1s1 U1566 (.Q(N6680), .DIN(N6280));
hi1s1 U1567 (.Q(N6681), .DIN(N6292));
hi1s1 U1568 (.Q(N6682), .DIN(N6307));
hi1s1 U1569 (.Q(N6683), .DIN(N6310));
nnd2s1 U1570 (.Q(N6689), .DIN1(N6325), .DIN2(N5120));
hi1s1 U1571 (.Q(N6690), .DIN(N6325));
nnd2s1 U1572 (.Q(N6691), .DIN1(N6328), .DIN2(N5622));
hi1s1 U1573 (.Q(N6692), .DIN(N6328));
and2s1 U1574 (.Q(N6693), .DIN1(N6149), .DIN2(N54));
hi1s1 U1575 (.Q(N6695), .DIN(N6331));
hi1s1 U1576 (.Q(N6698), .DIN(N6335));
nnd2s1 U1577 (.Q(N6699), .DIN1(N6338), .DIN2(N5956));
hi1s1 U1578 (.Q(N6700), .DIN(N6338));
hi1s1 U1579 (.Q(N6703), .DIN(N6175));
hi1s1 U1580 (.Q(N6708), .DIN(N6209));
hi1s1 U1581 (.Q(N6709), .DIN(N6212));
hi1s1 U1582 (.Q(N6710), .DIN(N6215));
hi1s1 U1583 (.Q(N6711), .DIN(N6218));
and3s1 U1584 (.Q(N6712), .DIN1(N5696), .DIN2(N5692), .DIN3(N6209));
and3s1 U1585 (.Q(N6713), .DIN1(N6200), .DIN2(N6197), .DIN3(N6212));
and3s1 U1586 (.Q(N6714), .DIN1(N5707), .DIN2(N5703), .DIN3(N6215));
and3s1 U1587 (.Q(N6715), .DIN1(N6206), .DIN2(N6203), .DIN3(N6218));
nb1s1 U1588 (.Q(N6716), .DIN(N6466));
and3s1 U1589 (.Q(N6718), .DIN1(N6164), .DIN2(N1777), .DIN3(N3130));
and3s1 U1590 (.Q(N6719), .DIN1(N5150), .DIN2(N5315), .DIN3(N6469));
and3s1 U1591 (.Q(N6720), .DIN1(N4524), .DIN2(N6025), .DIN3(N6470));
and3s1 U1592 (.Q(N6721), .DIN1(N5157), .DIN2(N5324), .DIN3(N6471));
and3s1 U1593 (.Q(N6722), .DIN1(N4532), .DIN2(N6028), .DIN3(N6472));
nnd2s1 U1594 (.Q(N6724), .DIN1(N6477), .DIN2(N6235));
hi1s1 U1595 (.Q(N6739), .DIN(N6271));
hi1s1 U1596 (.Q(N6740), .DIN(N6274));
hi1s1 U1597 (.Q(N6741), .DIN(N6277));
hi1s1 U1598 (.Q(N6744), .DIN(N6283));
hi1s1 U1599 (.Q(N6745), .DIN(N6286));
hi1s1 U1600 (.Q(N6746), .DIN(N6289));
hi1s1 U1601 (.Q(N6751), .DIN(N6295));
hi1s1 U1602 (.Q(N6752), .DIN(N6298));
hi1s1 U1603 (.Q(N6753), .DIN(N6301));
hi1s1 U1604 (.Q(N6754), .DIN(N6304));
hi1s1 U1605 (.Q(N6755), .DIN(N6322));
hi1s1 U1606 (.Q(N6760), .DIN(N6313));
hi1s1 U1607 (.Q(N6761), .DIN(N6316));
hi1s1 U1608 (.Q(N6762), .DIN(N6319));
hi1s1 U1609 (.Q(N6772), .DIN(N6341));
hi1s1 U1610 (.Q(N6773), .DIN(N6344));
hi1s1 U1611 (.Q(N6776), .DIN(N6347));
hi1s1 U1612 (.Q(N6777), .DIN(N6350));
hi1s1 U1613 (.Q(N6782), .DIN(N6353));
hi1s1 U1614 (.Q(N6783), .DIN(N6356));
hi1s1 U1615 (.Q(N6784), .DIN(N6359));
hi1s1 U1616 (.Q(N6785), .DIN(N6370));
hi1s1 U1617 (.Q(N6790), .DIN(N6364));
hi1s1 U1618 (.Q(N6791), .DIN(N6367));
nnd2s1 U1619 (.Q(N6792), .DIN1(N6630), .DIN2(N6631));
nnd2s1 U1620 (.Q(N6795), .DIN1(N6632), .DIN2(N6633));
and2s1 U1621 (.Q(N6801), .DIN1(N6108), .DIN2(N6415));
and2s1 U1622 (.Q(N6802), .DIN1(N6427), .DIN2(N6140));
and2s1 U1623 (.Q(N6803), .DIN1(N6397), .DIN2(N6080));
and2s1 U1624 (.Q(N6804), .DIN1(N6168), .DIN2(N6441));
hi1s1 U1625 (.Q(N6805), .DIN(N6466));
nnd2s1 U1626 (.Q(N6806), .DIN1(N1851), .DIN2(N6651));
hi1s1 U1627 (.Q(N6807), .DIN(N6482));
nnd2s1 U1628 (.Q(N6808), .DIN1(N6482), .DIN2(N6653));
hi1s1 U1629 (.Q(N6809), .DIN(N6486));
nnd2s1 U1630 (.Q(N6810), .DIN1(N6486), .DIN2(N6655));
hi1s1 U1631 (.Q(N6811), .DIN(N6490));
nnd2s1 U1632 (.Q(N6812), .DIN1(N6490), .DIN2(N6657));
hi1s1 U1633 (.Q(N6813), .DIN(N6494));
nnd2s1 U1634 (.Q(N6814), .DIN1(N6494), .DIN2(N6659));
nnd2s1 U1635 (.Q(N6815), .DIN1(N4575), .DIN2(N6661));
nnd2s1 U1636 (.Q(N6816), .DIN1(N5169), .DIN2(N6663));
or2s1 U1637 (.Q(N6817), .DIN1(N6397), .DIN2(N6664));
hi1s1 U1638 (.Q(N6823), .DIN(N6500));
nnd2s1 U1639 (.Q(N6824), .DIN1(N6500), .DIN2(N6666));
hi1s1 U1640 (.Q(N6825), .DIN(N6504));
nnd2s1 U1641 (.Q(N6826), .DIN1(N6504), .DIN2(N6668));
hi1s1 U1642 (.Q(N6827), .DIN(N6508));
nnd2s1 U1643 (.Q(N6828), .DIN1(N6508), .DIN2(N6670));
hi1s1 U1644 (.Q(N6829), .DIN(N6512));
nnd2s1 U1645 (.Q(N6830), .DIN1(N6512), .DIN2(N6672));
hi1s1 U1646 (.Q(N6831), .DIN(N6415));
hi1s1 U1647 (.Q(N6834), .DIN(N6566));
nnd2s1 U1648 (.Q(N6835), .DIN1(N6566), .DIN2(N5618));
hi1s1 U1649 (.Q(N6836), .DIN(N6569));
nnd2s1 U1650 (.Q(N6837), .DIN1(N6569), .DIN2(N5619));
hi1s1 U1651 (.Q(N6838), .DIN(N6572));
nnd2s1 U1652 (.Q(N6839), .DIN1(N6572), .DIN2(N5620));
hi1s1 U1653 (.Q(N6840), .DIN(N6575));
nnd2s1 U1654 (.Q(N6841), .DIN1(N6575), .DIN2(N5621));
nnd2s1 U1655 (.Q(N6842), .DIN1(N4627), .DIN2(N6690));
nnd2s1 U1656 (.Q(N6843), .DIN1(N5195), .DIN2(N6692));
or2s1 U1657 (.Q(N6844), .DIN1(N6427), .DIN2(N6693));
hi1s1 U1658 (.Q(N6850), .DIN(N6580));
nnd2s1 U1659 (.Q(N6851), .DIN1(N6580), .DIN2(N6695));
hi1s1 U1660 (.Q(N6852), .DIN(N6584));
nnd2s1 U1661 (.Q(N6853), .DIN1(N6584), .DIN2(N6434));
hi1s1 U1662 (.Q(N6854), .DIN(N6587));
nnd2s1 U1663 (.Q(N6855), .DIN1(N6587), .DIN2(N6698));
nnd2s1 U1664 (.Q(N6856), .DIN1(N5346), .DIN2(N6700));
hi1s1 U1665 (.Q(N6857), .DIN(N6441));
and3s1 U1666 (.Q(N6860), .DIN1(N6197), .DIN2(N5696), .DIN3(N6708));
and3s1 U1667 (.Q(N6861), .DIN1(N5692), .DIN2(N6200), .DIN3(N6709));
and3s1 U1668 (.Q(N6862), .DIN1(N6203), .DIN2(N5707), .DIN3(N6710));
and3s1 U1669 (.Q(N6863), .DIN1(N5703), .DIN2(N6206), .DIN3(N6711));
or3s1 U1670 (.Q(N6866), .DIN1(N4197), .DIN2(N6718), .DIN3(N3785));
nor2s1 U1671 (.Q(N6872), .DIN1(N6719), .DIN2(N6473));
nor2s1 U1672 (.Q(N6873), .DIN1(N6720), .DIN2(N6474));
nor2s1 U1673 (.Q(N6874), .DIN1(N6721), .DIN2(N6475));
nor2s1 U1674 (.Q(N6875), .DIN1(N6722), .DIN2(N6476));
hi1s1 U1675 (.Q(N6876), .DIN(N6637));
nb1s1 U1676 (.Q(N6877), .DIN(N6724));
and2s1 U1677 (.Q(N6879), .DIN1(N6045), .DIN2(N6478));
and2s1 U1678 (.Q(N6880), .DIN1(N6478), .DIN2(N132));
or2s1 U1679 (.Q(N6881), .DIN1(N6411), .DIN2(N6137));
hi1s1 U1680 (.Q(N6884), .DIN(N6516));
hi1s1 U1681 (.Q(N6885), .DIN(N6411));
hi1s1 U1682 (.Q(N6888), .DIN(N6526));
hi1s1 U1683 (.Q(N6889), .DIN(N6536));
nnd2s1 U1684 (.Q(N6890), .DIN1(N6536), .DIN2(N5176));
or2s1 U1685 (.Q(N6891), .DIN1(N6419), .DIN2(N6138));
hi1s1 U1686 (.Q(N6894), .DIN(N6539));
hi1s1 U1687 (.Q(N6895), .DIN(N6553));
nnd2s1 U1688 (.Q(N6896), .DIN1(N6553), .DIN2(N5728));
hi1s1 U1689 (.Q(N6897), .DIN(N6419));
hi1s1 U1690 (.Q(N6900), .DIN(N6556));
or2s1 U1691 (.Q(N6901), .DIN1(N6437), .DIN2(N6193));
hi1s1 U1692 (.Q(N6904), .DIN(N6592));
hi1s1 U1693 (.Q(N6905), .DIN(N6437));
hi1s1 U1694 (.Q(N6908), .DIN(N6599));
or2s1 U1695 (.Q(N6909), .DIN1(N6445), .DIN2(N6194));
hi1s1 U1696 (.Q(N6912), .DIN(N6606));
hi1s1 U1697 (.Q(N6913), .DIN(N6609));
hi1s1 U1698 (.Q(N6914), .DIN(N6619));
nnd2s1 U1699 (.Q(N6915), .DIN1(N6619), .DIN2(N5734));
hi1s1 U1700 (.Q(N6916), .DIN(N6445));
hi1s1 U1701 (.Q(N6919), .DIN(N6622));
hi1s1 U1702 (.Q(N6922), .DIN(N6634));
nnd2s1 U1703 (.Q(N6923), .DIN1(N6634), .DIN2(N6067));
or2s1 U1704 (.Q(N6924), .DIN1(N6382), .DIN2(N6801));
or2s1 U1705 (.Q(N6925), .DIN1(N6386), .DIN2(N6802));
or2s1 U1706 (.Q(N6926), .DIN1(N6388), .DIN2(N6803));
or2s1 U1707 (.Q(N6927), .DIN1(N6392), .DIN2(N6804));
hi1s1 U1708 (.Q(N6930), .DIN(N6724));
nnd2s1 U1709 (.Q(N6932), .DIN1(N6650), .DIN2(N6806));
nnd2s1 U1710 (.Q(N6935), .DIN1(N6241), .DIN2(N6807));
nnd2s1 U1711 (.Q(N6936), .DIN1(N6244), .DIN2(N6809));
nnd2s1 U1712 (.Q(N6937), .DIN1(N6247), .DIN2(N6811));
nnd2s1 U1713 (.Q(N6938), .DIN1(N6250), .DIN2(N6813));
nnd2s1 U1714 (.Q(N6939), .DIN1(N6660), .DIN2(N6815));
nnd2s1 U1715 (.Q(N6940), .DIN1(N6662), .DIN2(N6816));
nnd2s1 U1716 (.Q(N6946), .DIN1(N6259), .DIN2(N6823));
nnd2s1 U1717 (.Q(N6947), .DIN1(N6262), .DIN2(N6825));
nnd2s1 U1718 (.Q(N6948), .DIN1(N6265), .DIN2(N6827));
nnd2s1 U1719 (.Q(N6949), .DIN1(N6268), .DIN2(N6829));
nnd2s1 U1720 (.Q(N6953), .DIN1(N5183), .DIN2(N6834));
nnd2s1 U1721 (.Q(N6954), .DIN1(N5186), .DIN2(N6836));
nnd2s1 U1722 (.Q(N6955), .DIN1(N5189), .DIN2(N6838));
nnd2s1 U1723 (.Q(N6956), .DIN1(N5192), .DIN2(N6840));
nnd2s1 U1724 (.Q(N6957), .DIN1(N6689), .DIN2(N6842));
nnd2s1 U1725 (.Q(N6958), .DIN1(N6691), .DIN2(N6843));
nnd2s1 U1726 (.Q(N6964), .DIN1(N6331), .DIN2(N6850));
nnd2s1 U1727 (.Q(N6965), .DIN1(N6048), .DIN2(N6852));
nnd2s1 U1728 (.Q(N6966), .DIN1(N6335), .DIN2(N6854));
nnd2s1 U1729 (.Q(N6967), .DIN1(N6699), .DIN2(N6856));
nor2s1 U1730 (.Q(N6973), .DIN1(N6860), .DIN2(N6712));
nor2s1 U1731 (.Q(N6974), .DIN1(N6861), .DIN2(N6713));
nor2s1 U1732 (.Q(N6975), .DIN1(N6862), .DIN2(N6714));
nor2s1 U1733 (.Q(N6976), .DIN1(N6863), .DIN2(N6715));
hi1s1 U1734 (.Q(N6977), .DIN(N6792));
hi1s1 U1735 (.Q(N6978), .DIN(N6795));
or2s1 U1736 (.Q(N6979), .DIN1(N6879), .DIN2(N6880));
nnd2s1 U1737 (.Q(N6987), .DIN1(N4608), .DIN2(N6889));
nnd2s1 U1738 (.Q(N6990), .DIN1(N5177), .DIN2(N6895));
nnd2s1 U1739 (.Q(N6999), .DIN1(N5217), .DIN2(N6914));
nnd2s1 U1740 (.Q(N7002), .DIN1(N5377), .DIN2(N6922));
nnd2s1 U1741 (.Q(N7003), .DIN1(N6873), .DIN2(N6872));
nnd2s1 U1742 (.Q(N7006), .DIN1(N6875), .DIN2(N6874));
and3s1 U1743 (.Q(N7011), .DIN1(N6866), .DIN2(N2681), .DIN3(N2692));
and3s1 U1744 (.Q(N7012), .DIN1(N6866), .DIN2(N2756), .DIN3(N2767));
and3s1 U1745 (.Q(N7013), .DIN1(N6866), .DIN2(N2779), .DIN3(N2790));
hi1s1 U1746 (.Q(N7015), .DIN(N6866));
and3s1 U1747 (.Q(N7016), .DIN1(N6866), .DIN2(N2801), .DIN3(N2812));
nnd2s1 U1748 (.Q(N7018), .DIN1(N6935), .DIN2(N6808));
nnd2s1 U1749 (.Q(N7019), .DIN1(N6936), .DIN2(N6810));
nnd2s1 U1750 (.Q(N7020), .DIN1(N6937), .DIN2(N6812));
nnd2s1 U1751 (.Q(N7021), .DIN1(N6938), .DIN2(N6814));
hi1s1 U1752 (.Q(N7022), .DIN(N6939));
hi1s1 U1753 (.Q(N7023), .DIN(N6817));
nnd2s1 U1754 (.Q(N7028), .DIN1(N6946), .DIN2(N6824));
nnd2s1 U1755 (.Q(N7031), .DIN1(N6947), .DIN2(N6826));
nnd2s1 U1756 (.Q(N7034), .DIN1(N6948), .DIN2(N6828));
nnd2s1 U1757 (.Q(N7037), .DIN1(N6949), .DIN2(N6830));
and2s1 U1758 (.Q(N7040), .DIN1(N6817), .DIN2(N6079));
and2s1 U1759 (.Q(N7041), .DIN1(N6831), .DIN2(N6675));
nnd2s1 U1760 (.Q(N7044), .DIN1(N6953), .DIN2(N6835));
nnd2s1 U1761 (.Q(N7045), .DIN1(N6954), .DIN2(N6837));
nnd2s1 U1762 (.Q(N7046), .DIN1(N6955), .DIN2(N6839));
nnd2s1 U1763 (.Q(N7047), .DIN1(N6956), .DIN2(N6841));
hi1s1 U1764 (.Q(N7048), .DIN(N6957));
hi1s1 U1765 (.Q(N7049), .DIN(N6844));
nnd2s1 U1766 (.Q(N7054), .DIN1(N6964), .DIN2(N6851));
nnd2s1 U1767 (.Q(N7057), .DIN1(N6965), .DIN2(N6853));
nnd2s1 U1768 (.Q(N7060), .DIN1(N6966), .DIN2(N6855));
and2s1 U1769 (.Q(N7064), .DIN1(N6844), .DIN2(N6139));
and2s1 U1770 (.Q(N7065), .DIN1(N6857), .DIN2(N6703));
hi1s1 U1771 (.Q(N7072), .DIN(N6881));
nnd2s1 U1772 (.Q(N7073), .DIN1(N6881), .DIN2(N5172));
hi1s1 U1773 (.Q(N7074), .DIN(N6885));
nnd2s1 U1774 (.Q(N7075), .DIN1(N6885), .DIN2(N5727));
nnd2s1 U1775 (.Q(N7076), .DIN1(N6890), .DIN2(N6987));
hi1s1 U1776 (.Q(N7079), .DIN(N6891));
nnd2s1 U1777 (.Q(N7080), .DIN1(N6896), .DIN2(N6990));
hi1s1 U1778 (.Q(N7083), .DIN(N6897));
hi1s1 U1779 (.Q(N7084), .DIN(N6901));
nnd2s1 U1780 (.Q(N7085), .DIN1(N6901), .DIN2(N5198));
hi1s1 U1781 (.Q(N7086), .DIN(N6905));
nnd2s1 U1782 (.Q(N7087), .DIN1(N6905), .DIN2(N5731));
hi1s1 U1783 (.Q(N7088), .DIN(N6909));
nnd2s1 U1784 (.Q(N7089), .DIN1(N6909), .DIN2(N6912));
nnd2s1 U1785 (.Q(N7090), .DIN1(N6915), .DIN2(N6999));
hi1s1 U1786 (.Q(N7093), .DIN(N6916));
nnd2s1 U1787 (.Q(N7094), .DIN1(N6974), .DIN2(N6973));
nnd2s1 U1788 (.Q(N7097), .DIN1(N6976), .DIN2(N6975));
nnd2s1 U1789 (.Q(N7101), .DIN1(N7002), .DIN2(N6923));
hi1s1 U1790 (.Q(N7105), .DIN(N6932));
hi1s1 U1791 (.Q(N7110), .DIN(N6967));
and3s1 U1792 (.Q(N7114), .DIN1(N6979), .DIN2(N603), .DIN3(N1755));
hi1s1 U1793 (.Q(N7115), .DIN(N7019));
hi1s1 U1794 (.Q(N7116), .DIN(N7021));
and2s1 U1795 (.Q(N7125), .DIN1(N6817), .DIN2(N7018));
and2s1 U1796 (.Q(N7126), .DIN1(N6817), .DIN2(N7020));
and2s1 U1797 (.Q(N7127), .DIN1(N6817), .DIN2(N7022));
hi1s1 U1798 (.Q(N7130), .DIN(N7045));
hi1s1 U1799 (.Q(N7131), .DIN(N7047));
and2s1 U1800 (.Q(N7139), .DIN1(N6844), .DIN2(N7044));
and2s1 U1801 (.Q(N7140), .DIN1(N6844), .DIN2(N7046));
and2s1 U1802 (.Q(N7141), .DIN1(N6844), .DIN2(N7048));
and3s1 U1803 (.Q(N7146), .DIN1(N6932), .DIN2(N1761), .DIN3(N3108));
and3s1 U1804 (.Q(N7147), .DIN1(N6967), .DIN2(N1777), .DIN3(N3130));
hi1s1 U1805 (.Q(N7149), .DIN(N7003));
hi1s1 U1806 (.Q(N7150), .DIN(N7006));
nnd2s1 U1807 (.Q(N7151), .DIN1(N7006), .DIN2(N6876));
nnd2s1 U1808 (.Q(N7152), .DIN1(N4605), .DIN2(N7072));
nnd2s1 U1809 (.Q(N7153), .DIN1(N5173), .DIN2(N7074));
nnd2s1 U1810 (.Q(N7158), .DIN1(N4646), .DIN2(N7084));
nnd2s1 U1811 (.Q(N7159), .DIN1(N5205), .DIN2(N7086));
nnd2s1 U1812 (.Q(N7160), .DIN1(N6606), .DIN2(N7088));
hi1s1 U1813 (.Q(N7166), .DIN(N7037));
hi1s1 U1814 (.Q(N7167), .DIN(N7034));
hi1s1 U1815 (.Q(N7168), .DIN(N7031));
hi1s1 U1816 (.Q(N7169), .DIN(N7028));
hi1s1 U1817 (.Q(N7170), .DIN(N7060));
hi1s1 U1818 (.Q(N7171), .DIN(N7057));
hi1s1 U1819 (.Q(N7172), .DIN(N7054));
and2s1 U1820 (.Q(N7173), .DIN1(N7115), .DIN2(N7023));
and2s1 U1821 (.Q(N7174), .DIN1(N7116), .DIN2(N7023));
and2s1 U1822 (.Q(N7175), .DIN1(N6940), .DIN2(N7023));
and2s1 U1823 (.Q(N7176), .DIN1(N5418), .DIN2(N7023));
hi1s1 U1824 (.Q(N7177), .DIN(N7041));
and2s1 U1825 (.Q(N7178), .DIN1(N7130), .DIN2(N7049));
and2s1 U1826 (.Q(N7179), .DIN1(N7131), .DIN2(N7049));
and2s1 U1827 (.Q(N7180), .DIN1(N6958), .DIN2(N7049));
and2s1 U1828 (.Q(N7181), .DIN1(N5573), .DIN2(N7049));
hi1s1 U1829 (.Q(N7182), .DIN(N7065));
hi1s1 U1830 (.Q(N7183), .DIN(N7094));
nnd2s1 U1831 (.Q(N7184), .DIN1(N7094), .DIN2(N6977));
hi1s1 U1832 (.Q(N7185), .DIN(N7097));
nnd2s1 U1833 (.Q(N7186), .DIN1(N7097), .DIN2(N6978));
and3s1 U1834 (.Q(N7187), .DIN1(N7037), .DIN2(N1761), .DIN3(N3108));
and3s1 U1835 (.Q(N7188), .DIN1(N7034), .DIN2(N1761), .DIN3(N3108));
and3s1 U1836 (.Q(N7189), .DIN1(N7031), .DIN2(N1761), .DIN3(N3108));
or3s1 U1837 (.Q(N7190), .DIN1(N4956), .DIN2(N7146), .DIN3(N3781));
and3s1 U1838 (.Q(N7196), .DIN1(N7060), .DIN2(N1777), .DIN3(N3130));
and3s1 U1839 (.Q(N7197), .DIN1(N7057), .DIN2(N1777), .DIN3(N3130));
or3s1 U1840 (.Q(N7198), .DIN1(N4960), .DIN2(N7147), .DIN3(N3786));
nnd2s1 U1841 (.Q(N7204), .DIN1(N7101), .DIN2(N7149));
hi1s1 U1842 (.Q(N7205), .DIN(N7101));
nnd2s1 U1843 (.Q(N7206), .DIN1(N6637), .DIN2(N7150));
and3s1 U1844 (.Q(N7207), .DIN1(N7028), .DIN2(N1793), .DIN3(N3158));
and3s1 U1845 (.Q(N7208), .DIN1(N7054), .DIN2(N1807), .DIN3(N3180));
nnd2s1 U1846 (.Q(N7209), .DIN1(N7073), .DIN2(N7152));
nnd2s1 U1847 (.Q(N7212), .DIN1(N7075), .DIN2(N7153));
hi1s1 U1848 (.Q(N7215), .DIN(N7076));
nnd2s1 U1849 (.Q(N7216), .DIN1(N7076), .DIN2(N7079));
hi1s1 U1850 (.Q(N7217), .DIN(N7080));
nnd2s1 U1851 (.Q(N7218), .DIN1(N7080), .DIN2(N7083));
nnd2s1 U1852 (.Q(N7219), .DIN1(N7085), .DIN2(N7158));
nnd2s1 U1853 (.Q(N7222), .DIN1(N7087), .DIN2(N7159));
nnd2s1 U1854 (.Q(N7225), .DIN1(N7089), .DIN2(N7160));
hi1s1 U1855 (.Q(N7228), .DIN(N7090));
nnd2s1 U1856 (.Q(N7229), .DIN1(N7090), .DIN2(N7093));
or2s1 U1857 (.Q(N7236), .DIN1(N7173), .DIN2(N7125));
or2s1 U1858 (.Q(N7239), .DIN1(N7174), .DIN2(N7126));
or2s1 U1859 (.Q(N7242), .DIN1(N7175), .DIN2(N7127));
or2s1 U1860 (.Q(N7245), .DIN1(N7176), .DIN2(N7040));
or2s1 U1861 (.Q(N7250), .DIN1(N7178), .DIN2(N7139));
or2s1 U1862 (.Q(N7257), .DIN1(N7179), .DIN2(N7140));
or2s1 U1863 (.Q(N7260), .DIN1(N7180), .DIN2(N7141));
or2s1 U1864 (.Q(N7263), .DIN1(N7181), .DIN2(N7064));
nnd2s1 U1865 (.Q(N7268), .DIN1(N6792), .DIN2(N7183));
nnd2s1 U1866 (.Q(N7269), .DIN1(N6795), .DIN2(N7185));
or3s1 U1867 (.Q(N7270), .DIN1(N4957), .DIN2(N7187), .DIN3(N3782));
or3s1 U1868 (.Q(N7276), .DIN1(N4958), .DIN2(N7188), .DIN3(N3783));
or3s1 U1869 (.Q(N7282), .DIN1(N4959), .DIN2(N7189), .DIN3(N3784));
or3s1 U1870 (.Q(N7288), .DIN1(N4961), .DIN2(N7196), .DIN3(N3787));
or3s1 U1871 (.Q(N7294), .DIN1(N3998), .DIN2(N7197), .DIN3(N3788));
nnd2s1 U1872 (.Q(N7300), .DIN1(N7003), .DIN2(N7205));
nnd2s1 U1873 (.Q(N7301), .DIN1(N7206), .DIN2(N7151));
or3s1 U1874 (.Q(N7304), .DIN1(N4980), .DIN2(N7207), .DIN3(N3800));
or3s1 U1875 (.Q(N7310), .DIN1(N4984), .DIN2(N7208), .DIN3(N3805));
nnd2s1 U1876 (.Q(N7320), .DIN1(N6891), .DIN2(N7215));
nnd2s1 U1877 (.Q(N7321), .DIN1(N6897), .DIN2(N7217));
nnd2s1 U1878 (.Q(N7328), .DIN1(N6916), .DIN2(N7228));
and3s1 U1879 (.Q(N7338), .DIN1(N7190), .DIN2(N1185), .DIN3(N2692));
and3s1 U1880 (.Q(N7339), .DIN1(N7198), .DIN2(N2681), .DIN3(N2692));
and3s1 U1881 (.Q(N7340), .DIN1(N7190), .DIN2(N1247), .DIN3(N2767));
and3s1 U1882 (.Q(N7341), .DIN1(N7198), .DIN2(N2756), .DIN3(N2767));
and3s1 U1883 (.Q(N7342), .DIN1(N7190), .DIN2(N1327), .DIN3(N2790));
and3s1 U1884 (.Q(N7349), .DIN1(N7198), .DIN2(N2779), .DIN3(N2790));
and3s1 U1885 (.Q(N7357), .DIN1(N7198), .DIN2(N2801), .DIN3(N2812));
hi1s1 U1886 (.Q(N7363), .DIN(N7198));
and3s1 U1887 (.Q(N7364), .DIN1(N7190), .DIN2(N1351), .DIN3(N2812));
hi1s1 U1888 (.Q(N7365), .DIN(N7190));
nnd2s1 U1889 (.Q(N7394), .DIN1(N7268), .DIN2(N7184));
nnd2s1 U1890 (.Q(N7397), .DIN1(N7269), .DIN2(N7186));
nnd2s1 U1891 (.Q(N7402), .DIN1(N7204), .DIN2(N7300));
hi1s1 U1892 (.Q(N7405), .DIN(N7209));
nnd2s1 U1893 (.Q(N7406), .DIN1(N7209), .DIN2(N6884));
hi1s1 U1894 (.Q(N7407), .DIN(N7212));
nnd2s1 U1895 (.Q(N7408), .DIN1(N7212), .DIN2(N6888));
nnd2s1 U1896 (.Q(N7409), .DIN1(N7320), .DIN2(N7216));
nnd2s1 U1897 (.Q(N7412), .DIN1(N7321), .DIN2(N7218));
hi1s1 U1898 (.Q(N7415), .DIN(N7219));
nnd2s1 U1899 (.Q(N7416), .DIN1(N7219), .DIN2(N6904));
hi1s1 U1900 (.Q(N7417), .DIN(N7222));
nnd2s1 U1901 (.Q(N7418), .DIN1(N7222), .DIN2(N6908));
hi1s1 U1902 (.Q(N7419), .DIN(N7225));
nnd2s1 U1903 (.Q(N7420), .DIN1(N7225), .DIN2(N6913));
nnd2s1 U1904 (.Q(N7421), .DIN1(N7328), .DIN2(N7229));
hi1s1 U1905 (.Q(N7424), .DIN(N7245));
hi1s1 U1906 (.Q(N7425), .DIN(N7242));
hi1s1 U1907 (.Q(N7426), .DIN(N7239));
hi1s1 U1908 (.Q(N7427), .DIN(N7236));
hi1s1 U1909 (.Q(N7428), .DIN(N7263));
hi1s1 U1910 (.Q(N7429), .DIN(N7260));
hi1s1 U1911 (.Q(N7430), .DIN(N7257));
hi1s1 U1912 (.Q(N7431), .DIN(N7250));
hi1s1 U1913 (.Q(N7432), .DIN(N7250));
and3s1 U1914 (.Q(N7433), .DIN1(N7310), .DIN2(N2653), .DIN3(N2664));
and3s1 U1915 (.Q(N7434), .DIN1(N7304), .DIN2(N1161), .DIN3(N2664));
or4s1 U1916 (.Q(N7435), .DIN1(N7011), .DIN2(N7338), .DIN3(N3621), .DIN4(N2591));
and3s1 U1917 (.Q(N7436), .DIN1(N7270), .DIN2(N1185), .DIN3(N2692));
and3s1 U1918 (.Q(N7437), .DIN1(N7288), .DIN2(N2681), .DIN3(N2692));
and3s1 U1919 (.Q(N7438), .DIN1(N7276), .DIN2(N1185), .DIN3(N2692));
and3s1 U1920 (.Q(N7439), .DIN1(N7294), .DIN2(N2681), .DIN3(N2692));
and3s1 U1921 (.Q(N7440), .DIN1(N7282), .DIN2(N1185), .DIN3(N2692));
and3s1 U1922 (.Q(N7441), .DIN1(N7310), .DIN2(N2728), .DIN3(N2739));
and3s1 U1923 (.Q(N7442), .DIN1(N7304), .DIN2(N1223), .DIN3(N2739));
or4s1 U1924 (.Q(N7443), .DIN1(N7012), .DIN2(N7340), .DIN3(N3632), .DIN4(N2600));
and3s1 U1925 (.Q(N7444), .DIN1(N7270), .DIN2(N1247), .DIN3(N2767));
and3s1 U1926 (.Q(N7445), .DIN1(N7288), .DIN2(N2756), .DIN3(N2767));
and3s1 U1927 (.Q(N7446), .DIN1(N7276), .DIN2(N1247), .DIN3(N2767));
and3s1 U1928 (.Q(N7447), .DIN1(N7294), .DIN2(N2756), .DIN3(N2767));
and3s1 U1929 (.Q(N7448), .DIN1(N7282), .DIN2(N1247), .DIN3(N2767));
or4s1 U1930 (.Q(N7449), .DIN1(N7013), .DIN2(N7342), .DIN3(N3641), .DIN4(N2605));
and3s1 U1931 (.Q(N7450), .DIN1(N7310), .DIN2(N3041), .DIN3(N3052));
and3s1 U1932 (.Q(N7451), .DIN1(N7304), .DIN2(N1697), .DIN3(N3052));
and3s1 U1933 (.Q(N7452), .DIN1(N7294), .DIN2(N2779), .DIN3(N2790));
and3s1 U1934 (.Q(N7453), .DIN1(N7282), .DIN2(N1327), .DIN3(N2790));
and3s1 U1935 (.Q(N7454), .DIN1(N7288), .DIN2(N2779), .DIN3(N2790));
and3s1 U1936 (.Q(N7455), .DIN1(N7276), .DIN2(N1327), .DIN3(N2790));
and3s1 U1937 (.Q(N7456), .DIN1(N7270), .DIN2(N1327), .DIN3(N2790));
and3s1 U1938 (.Q(N7457), .DIN1(N7310), .DIN2(N3075), .DIN3(N3086));
and3s1 U1939 (.Q(N7458), .DIN1(N7304), .DIN2(N1731), .DIN3(N3086));
and3s1 U1940 (.Q(N7459), .DIN1(N7294), .DIN2(N2801), .DIN3(N2812));
and3s1 U1941 (.Q(N7460), .DIN1(N7282), .DIN2(N1351), .DIN3(N2812));
and3s1 U1942 (.Q(N7461), .DIN1(N7288), .DIN2(N2801), .DIN3(N2812));
and3s1 U1943 (.Q(N7462), .DIN1(N7276), .DIN2(N1351), .DIN3(N2812));
and3s1 U1944 (.Q(N7463), .DIN1(N7270), .DIN2(N1351), .DIN3(N2812));
and3s1 U1945 (.Q(N7464), .DIN1(N7250), .DIN2(N603), .DIN3(N599));
hi1s1 U1946 (.Q(N7465), .DIN(N7310));
hi1s1 U1947 (.Q(N7466), .DIN(N7294));
hi1s1 U1948 (.Q(N7467), .DIN(N7288));
hi1s1 U1949 (.Q(N7468), .DIN(N7301));
or4s1 U1950 (.Q(N7469), .DIN1(N7016), .DIN2(N7364), .DIN3(N3660), .DIN4(N2626));
hi1s1 U1951 (.Q(N7470), .DIN(N7304));
hi1s1 U1952 (.Q(N7471), .DIN(N7282));
hi1s1 U1953 (.Q(N7472), .DIN(N7276));
hi1s1 U1954 (.Q(N7473), .DIN(N7270));
nb1s1 U1955 (.Q(N7474), .DIN(N7394));
nb1s1 U1956 (.Q(N7476), .DIN(N7397));
and2s1 U1957 (.Q(N7479), .DIN1(N7301), .DIN2(N3068));
and3s1 U1958 (.Q(N7481), .DIN1(N7245), .DIN2(N1793), .DIN3(N3158));
and3s1 U1959 (.Q(N7482), .DIN1(N7242), .DIN2(N1793), .DIN3(N3158));
and3s1 U1960 (.Q(N7483), .DIN1(N7239), .DIN2(N1793), .DIN3(N3158));
and3s1 U1961 (.Q(N7484), .DIN1(N7236), .DIN2(N1793), .DIN3(N3158));
and3s1 U1962 (.Q(N7485), .DIN1(N7263), .DIN2(N1807), .DIN3(N3180));
and3s1 U1963 (.Q(N7486), .DIN1(N7260), .DIN2(N1807), .DIN3(N3180));
and3s1 U1964 (.Q(N7487), .DIN1(N7257), .DIN2(N1807), .DIN3(N3180));
and3s1 U1965 (.Q(N7488), .DIN1(N7250), .DIN2(N1807), .DIN3(N3180));
nnd2s1 U1966 (.Q(N7489), .DIN1(N6979), .DIN2(N7250));
nnd2s1 U1967 (.Q(N7492), .DIN1(N6516), .DIN2(N7405));
nnd2s1 U1968 (.Q(N7493), .DIN1(N6526), .DIN2(N7407));
nnd2s1 U1969 (.Q(N7498), .DIN1(N6592), .DIN2(N7415));
nnd2s1 U1970 (.Q(N7499), .DIN1(N6599), .DIN2(N7417));
nnd2s1 U1971 (.Q(N7500), .DIN1(N6609), .DIN2(N7419));
and9s1 U1972 (.Q(N7503), .DIN1(N7105), .DIN2(N7166), .DIN3(N7167), .DIN4(N7168), .DIN5(N7169), .DIN6(N7424), .DIN7(N7425), .DIN8(N7426), .DIN9(N7427));
and9s1 U1973 (.Q(N7504), .DIN1(N6640), .DIN2(N7110), .DIN3(N7170), .DIN4(N7171), .DIN5(N7172), .DIN6(N7428), .DIN7(N7429), .DIN8(N7430), .DIN9(N7431));
or4s1 U1974 (.Q(N7505), .DIN1(N7433), .DIN2(N7434), .DIN3(N3616), .DIN4(N2585));
and2s1 U1975 (.Q(N7506), .DIN1(N7435), .DIN2(N2675));
or4s1 U1976 (.Q(N7507), .DIN1(N7339), .DIN2(N7436), .DIN3(N3622), .DIN4(N2592));
or4s1 U1977 (.Q(N7508), .DIN1(N7437), .DIN2(N7438), .DIN3(N3623), .DIN4(N2593));
or4s1 U1978 (.Q(N7509), .DIN1(N7439), .DIN2(N7440), .DIN3(N3624), .DIN4(N2594));
or4s1 U1979 (.Q(N7510), .DIN1(N7441), .DIN2(N7442), .DIN3(N3627), .DIN4(N2595));
and2s1 U1980 (.Q(N7511), .DIN1(N7443), .DIN2(N2750));
or4s1 U1981 (.Q(N7512), .DIN1(N7341), .DIN2(N7444), .DIN3(N3633), .DIN4(N2601));
or4s1 U1982 (.Q(N7513), .DIN1(N7445), .DIN2(N7446), .DIN3(N3634), .DIN4(N2602));
or4s1 U1983 (.Q(N7514), .DIN1(N7447), .DIN2(N7448), .DIN3(N3635), .DIN4(N2603));
or4s1 U1984 (.Q(N7515), .DIN1(N7450), .DIN2(N7451), .DIN3(N3646), .DIN4(N2610));
or4s1 U1985 (.Q(N7516), .DIN1(N7452), .DIN2(N7453), .DIN3(N3647), .DIN4(N2611));
or4s1 U1986 (.Q(N7517), .DIN1(N7454), .DIN2(N7455), .DIN3(N3648), .DIN4(N2612));
or4s1 U1987 (.Q(N7518), .DIN1(N7349), .DIN2(N7456), .DIN3(N3649), .DIN4(N2613));
or4s1 U1988 (.Q(N7519), .DIN1(N7457), .DIN2(N7458), .DIN3(N3654), .DIN4(N2618));
or4s1 U1989 (.Q(N7520), .DIN1(N7459), .DIN2(N7460), .DIN3(N3655), .DIN4(N2619));
or4s1 U1990 (.Q(N7521), .DIN1(N7461), .DIN2(N7462), .DIN3(N3656), .DIN4(N2620));
or4s1 U1991 (.Q(N7522), .DIN1(N7357), .DIN2(N7463), .DIN3(N3657), .DIN4(N2621));
or4s1 U1992 (.Q(N7525), .DIN1(N4741), .DIN2(N7114), .DIN3(N2624), .DIN4(N7464));
and3s1 U1993 (.Q(N7526), .DIN1(N7468), .DIN2(N3119), .DIN3(N3130));
hi1s1 U1994 (.Q(N7527), .DIN(N7394));
hi1s1 U1995 (.Q(N7528), .DIN(N7397));
hi1s1 U1996 (.Q(N7529), .DIN(N7402));
and2s1 U1997 (.Q(N7530), .DIN1(N7402), .DIN2(N3068));
or3s1 U1998 (.Q(N7531), .DIN1(N4981), .DIN2(N7481), .DIN3(N3801));
or3s1 U1999 (.Q(N7537), .DIN1(N4982), .DIN2(N7482), .DIN3(N3802));
or3s1 U2000 (.Q(N7543), .DIN1(N4983), .DIN2(N7483), .DIN3(N3803));
or3s1 U2001 (.Q(N7549), .DIN1(N5165), .DIN2(N7484), .DIN3(N3804));
or3s1 U2002 (.Q(N7555), .DIN1(N4985), .DIN2(N7485), .DIN3(N3806));
or3s1 U2003 (.Q(N7561), .DIN1(N4986), .DIN2(N7486), .DIN3(N3807));
or3s1 U2004 (.Q(N7567), .DIN1(N4547), .DIN2(N7487), .DIN3(N3808));
or3s1 U2005 (.Q(N7573), .DIN1(N4987), .DIN2(N7488), .DIN3(N3809));
nnd2s1 U2006 (.Q(N7579), .DIN1(N7492), .DIN2(N7406));
nnd2s1 U2007 (.Q(N7582), .DIN1(N7493), .DIN2(N7408));
hi1s1 U2008 (.Q(N7585), .DIN(N7409));
nnd2s1 U2009 (.Q(N7586), .DIN1(N7409), .DIN2(N6894));
hi1s1 U2010 (.Q(N7587), .DIN(N7412));
nnd2s1 U2011 (.Q(N7588), .DIN1(N7412), .DIN2(N6900));
nnd2s1 U2012 (.Q(N7589), .DIN1(N7498), .DIN2(N7416));
nnd2s1 U2013 (.Q(N7592), .DIN1(N7499), .DIN2(N7418));
nnd2s1 U2014 (.Q(N7595), .DIN1(N7500), .DIN2(N7420));
hi1s1 U2015 (.Q(N7598), .DIN(N7421));
nnd2s1 U2016 (.Q(N7599), .DIN1(N7421), .DIN2(N6919));
and2s1 U2017 (.Q(N7600), .DIN1(N7505), .DIN2(N2647));
and2s1 U2018 (.Q(N7601), .DIN1(N7507), .DIN2(N2675));
and2s1 U2019 (.Q(N7602), .DIN1(N7508), .DIN2(N2675));
and2s1 U2020 (.Q(N7603), .DIN1(N7509), .DIN2(N2675));
and2s1 U2021 (.Q(N7604), .DIN1(N7510), .DIN2(N2722));
and2s1 U2022 (.Q(N7605), .DIN1(N7512), .DIN2(N2750));
and2s1 U2023 (.Q(N7606), .DIN1(N7513), .DIN2(N2750));
and2s1 U2024 (.Q(N7607), .DIN1(N7514), .DIN2(N2750));
and2s1 U2025 (.Q(N7624), .DIN1(N6979), .DIN2(N7489));
and2s1 U2026 (.Q(N7625), .DIN1(N7489), .DIN2(N7250));
and2s1 U2027 (.Q(N7626), .DIN1(N1149), .DIN2(N7525));
and5s1 U2028 (.Q(N7631), .DIN1(N562), .DIN2(N7527), .DIN3(N7528), .DIN4(N6805), .DIN5(N6930));
and3s1 U2029 (.Q(N7636), .DIN1(N7529), .DIN2(N3097), .DIN3(N3108));
nnd2s1 U2030 (.Q(N7657), .DIN1(N6539), .DIN2(N7585));
nnd2s1 U2031 (.Q(N7658), .DIN1(N6556), .DIN2(N7587));
nnd2s1 U2032 (.Q(N7665), .DIN1(N6622), .DIN2(N7598));
and3s1 U2033 (.Q(N7666), .DIN1(N7555), .DIN2(N2653), .DIN3(N2664));
and3s1 U2034 (.Q(N7667), .DIN1(N7531), .DIN2(N1161), .DIN3(N2664));
and3s1 U2035 (.Q(N7668), .DIN1(N7561), .DIN2(N2653), .DIN3(N2664));
and3s1 U2036 (.Q(N7669), .DIN1(N7537), .DIN2(N1161), .DIN3(N2664));
and3s1 U2037 (.Q(N7670), .DIN1(N7567), .DIN2(N2653), .DIN3(N2664));
and3s1 U2038 (.Q(N7671), .DIN1(N7543), .DIN2(N1161), .DIN3(N2664));
and3s1 U2039 (.Q(N7672), .DIN1(N7573), .DIN2(N2653), .DIN3(N2664));
and3s1 U2040 (.Q(N7673), .DIN1(N7549), .DIN2(N1161), .DIN3(N2664));
and3s1 U2041 (.Q(N7674), .DIN1(N7555), .DIN2(N2728), .DIN3(N2739));
and3s1 U2042 (.Q(N7675), .DIN1(N7531), .DIN2(N1223), .DIN3(N2739));
and3s1 U2043 (.Q(N7676), .DIN1(N7561), .DIN2(N2728), .DIN3(N2739));
and3s1 U2044 (.Q(N7677), .DIN1(N7537), .DIN2(N1223), .DIN3(N2739));
and3s1 U2045 (.Q(N7678), .DIN1(N7567), .DIN2(N2728), .DIN3(N2739));
and3s1 U2046 (.Q(N7679), .DIN1(N7543), .DIN2(N1223), .DIN3(N2739));
and3s1 U2047 (.Q(N7680), .DIN1(N7573), .DIN2(N2728), .DIN3(N2739));
and3s1 U2048 (.Q(N7681), .DIN1(N7549), .DIN2(N1223), .DIN3(N2739));
and3s1 U2049 (.Q(N7682), .DIN1(N7573), .DIN2(N3075), .DIN3(N3086));
and3s1 U2050 (.Q(N7683), .DIN1(N7549), .DIN2(N1731), .DIN3(N3086));
and3s1 U2051 (.Q(N7684), .DIN1(N7573), .DIN2(N3041), .DIN3(N3052));
and3s1 U2052 (.Q(N7685), .DIN1(N7549), .DIN2(N1697), .DIN3(N3052));
and3s1 U2053 (.Q(N7686), .DIN1(N7567), .DIN2(N3041), .DIN3(N3052));
and3s1 U2054 (.Q(N7687), .DIN1(N7543), .DIN2(N1697), .DIN3(N3052));
and3s1 U2055 (.Q(N7688), .DIN1(N7561), .DIN2(N3041), .DIN3(N3052));
and3s1 U2056 (.Q(N7689), .DIN1(N7537), .DIN2(N1697), .DIN3(N3052));
and3s1 U2057 (.Q(N7690), .DIN1(N7555), .DIN2(N3041), .DIN3(N3052));
and3s1 U2058 (.Q(N7691), .DIN1(N7531), .DIN2(N1697), .DIN3(N3052));
and3s1 U2059 (.Q(N7692), .DIN1(N7567), .DIN2(N3075), .DIN3(N3086));
and3s1 U2060 (.Q(N7693), .DIN1(N7543), .DIN2(N1731), .DIN3(N3086));
and3s1 U2061 (.Q(N7694), .DIN1(N7561), .DIN2(N3075), .DIN3(N3086));
and3s1 U2062 (.Q(N7695), .DIN1(N7537), .DIN2(N1731), .DIN3(N3086));
and3s1 U2063 (.Q(N7696), .DIN1(N7555), .DIN2(N3075), .DIN3(N3086));
and3s1 U2064 (.Q(N7697), .DIN1(N7531), .DIN2(N1731), .DIN3(N3086));
or2s1 U2065 (.Q(N7698), .DIN1(N7624), .DIN2(N7625));
hi1s1 U2066 (.Q(N7699), .DIN(N7573));
hi1s1 U2067 (.Q(N7700), .DIN(N7567));
hi1s1 U2068 (.Q(N7701), .DIN(N7561));
hi1s1 U2069 (.Q(N7702), .DIN(N7555));
and3s1 U2070 (.Q(N7703), .DIN1(N1156), .DIN2(N7631), .DIN3(N245));
hi1s1 U2071 (.Q(N7704), .DIN(N7549));
hi1s1 U2072 (.Q(N7705), .DIN(N7543));
hi1s1 U2073 (.Q(N7706), .DIN(N7537));
hi1s1 U2074 (.Q(N7707), .DIN(N7531));
hi1s1 U2075 (.Q(N7708), .DIN(N7579));
nnd2s1 U2076 (.Q( tempN7709 ), .DIN1(N7579), .DIN2(N6739));
hi1s1 U2077 (.Q(N7710), .DIN(N7582));
nnd2s1 U2078 (.Q(N7711), .DIN1(N7582), .DIN2(N6744));
nnd2s1 U2079 (.Q(N7712), .DIN1(N7657), .DIN2(N7586));
nnd2s1 U2080 (.Q(N7715), .DIN1(N7658), .DIN2(N7588));
hi1s1 U2081 (.Q(N7718), .DIN(N7589));
nnd2s1 U2082 (.Q(N7719), .DIN1(N7589), .DIN2(N6772));
hi1s1 U2083 (.Q(N7720), .DIN(N7592));
nnd2s1 U2084 (.Q(N7721), .DIN1(N7592), .DIN2(N6776));
hi1s1 U2085 (.Q(N7722), .DIN(N7595));
nnd2s1 U2086 (.Q(N7723), .DIN1(N7595), .DIN2(N5733));
nnd2s1 U2087 (.Q(N7724), .DIN1(N7665), .DIN2(N7599));
or4s1 U2088 (.Q(N7727), .DIN1(N7666), .DIN2(N7667), .DIN3(N3617), .DIN4(N2586));
or4s1 U2089 (.Q(N7728), .DIN1(N7668), .DIN2(N7669), .DIN3(N3618), .DIN4(N2587));
or4s1 U2090 (.Q(N7729), .DIN1(N7670), .DIN2(N7671), .DIN3(N3619), .DIN4(N2588));
or4s1 U2091 (.Q(N7730), .DIN1(N7672), .DIN2(N7673), .DIN3(N3620), .DIN4(N2589));
or4s1 U2092 (.Q(N7731), .DIN1(N7674), .DIN2(N7675), .DIN3(N3628), .DIN4(N2596));
or4s1 U2093 (.Q(N7732), .DIN1(N7676), .DIN2(N7677), .DIN3(N3629), .DIN4(N2597));
or4s1 U2094 (.Q(N7733), .DIN1(N7678), .DIN2(N7679), .DIN3(N3630), .DIN4(N2598));
or4s1 U2095 (.Q(N7734), .DIN1(N7680), .DIN2(N7681), .DIN3(N3631), .DIN4(N2599));
or4s1 U2096 (.Q(N7735), .DIN1(N7682), .DIN2(N7683), .DIN3(N3638), .DIN4(N2604));
or4s1 U2097 (.Q(N7736), .DIN1(N7684), .DIN2(N7685), .DIN3(N3642), .DIN4(N2606));
or4s1 U2098 (.Q(N7737), .DIN1(N7686), .DIN2(N7687), .DIN3(N3643), .DIN4(N2607));
or4s1 U2099 (.Q(N7738), .DIN1(N7688), .DIN2(N7689), .DIN3(N3644), .DIN4(N2608));
or4s1 U2100 (.Q(N7739), .DIN1(N7690), .DIN2(N7691), .DIN3(N3645), .DIN4(N2609));
or4s1 U2101 (.Q(N7740), .DIN1(N7692), .DIN2(N7693), .DIN3(N3651), .DIN4(N2615));
or4s1 U2102 (.Q(N7741), .DIN1(N7694), .DIN2(N7695), .DIN3(N3652), .DIN4(N2616));
or4s1 U2103 (.Q(N7742), .DIN1(N7696), .DIN2(N7697), .DIN3(N3653), .DIN4(N2617));
nnd2s1 U2104 (.Q(N7743), .DIN1(N6271), .DIN2(N7708));
nnd2s1 U2105 (.Q(N7744), .DIN1(N6283), .DIN2(N7710));
nnd2s1 U2106 (.Q(N7749), .DIN1(N6341), .DIN2(N7718));
nnd2s1 U2107 (.Q(N7750), .DIN1(N6347), .DIN2(N7720));
nnd2s1 U2108 (.Q(N7751), .DIN1(N5214), .DIN2(N7722));
and2s1 U2109 (.Q(N7754), .DIN1(N7727), .DIN2(N2647));
and2s1 U2110 (.Q(N7755), .DIN1(N7728), .DIN2(N2647));
and2s1 U2111 (.Q(N7756), .DIN1(N7729), .DIN2(N2647));
and2s1 U2112 (.Q(N7757), .DIN1(N7730), .DIN2(N2647));
and2s1 U2113 (.Q(N7758), .DIN1(N7731), .DIN2(N2722));
and2s1 U2114 (.Q(N7759), .DIN1(N7732), .DIN2(N2722));
and2s1 U2115 (.Q(N7760), .DIN1(N7733), .DIN2(N2722));
and2s1 U2116 (.Q(N7761), .DIN1(N7734), .DIN2(N2722));
nnd2s1 U2117 (.Q(N7762), .DIN1(N7743), .DIN2(N7709));
nnd2s1 U2118 (.Q(N7765), .DIN1(N7744), .DIN2(N7711));
hi1s1 U2119 (.Q(N7768), .DIN(N7712));
nnd2s1 U2120 (.Q(N7769), .DIN1(N7712), .DIN2(N6751));
hi1s1 U2121 (.Q(N7770), .DIN(N7715));
nnd2s1 U2122 (.Q(N7771), .DIN1(N7715), .DIN2(N6760));
nnd2s1 U2123 (.Q(N7772), .DIN1(N7749), .DIN2(N7719));
nnd2s1 U2124 (.Q(N7775), .DIN1(N7750), .DIN2(N7721));
nnd2s1 U2125 (.Q(N7778), .DIN1(N7751), .DIN2(N7723));
hi1s1 U2126 (.Q(N7781), .DIN(N7724));
nnd2s1 U2127 (.Q(N7782), .DIN1(N7724), .DIN2(N5735));
nnd2s1 U2128 (.Q(N7787), .DIN1(N6295), .DIN2(N7768));
nnd2s1 U2129 (.Q(N7788), .DIN1(N6313), .DIN2(N7770));
nnd2s1 U2130 (.Q(N7795), .DIN1(N5220), .DIN2(N7781));
hi1s1 U2131 (.Q(N7796), .DIN(N7762));
nnd2s1 U2132 (.Q(N7797), .DIN1(N7762), .DIN2(N6740));
hi1s1 U2133 (.Q(N7798), .DIN(N7765));
nnd2s1 U2134 (.Q(N7799), .DIN1(N7765), .DIN2(N6745));
nnd2s1 U2135 (.Q(N7800), .DIN1(N7787), .DIN2(N7769));
nnd2s1 U2136 (.Q(N7803), .DIN1(N7788), .DIN2(N7771));
hi1s1 U2137 (.Q(N7806), .DIN(N7772));
nnd2s1 U2138 (.Q(N7807), .DIN1(N7772), .DIN2(N6773));
hi1s1 U2139 (.Q(N7808), .DIN(N7775));
nnd2s1 U2140 (.Q(N7809), .DIN1(N7775), .DIN2(N6777));
hi1s1 U2141 (.Q(N7810), .DIN(N7778));
nnd2s1 U2142 (.Q(N7811), .DIN1(N7778), .DIN2(N6782));
nnd2s1 U2143 (.Q(N7812), .DIN1(N7795), .DIN2(N7782));
nnd2s1 U2144 (.Q(N7815), .DIN1(N6274), .DIN2(N7796));
nnd2s1 U2145 (.Q(N7816), .DIN1(N6286), .DIN2(N7798));
nnd2s1 U2146 (.Q(N7821), .DIN1(N6344), .DIN2(N7806));
nnd2s1 U2147 (.Q(N7822), .DIN1(N6350), .DIN2(N7808));
nnd2s1 U2148 (.Q(N7823), .DIN1(N6353), .DIN2(N7810));
nnd2s1 U2149 (.Q(N7826), .DIN1(N7815), .DIN2(N7797));
nnd2s1 U2150 (.Q(N7829), .DIN1(N7816), .DIN2(N7799));
hi1s1 U2151 (.Q(N7832), .DIN(N7800));
nnd2s1 U2152 (.Q(N7833), .DIN1(N7800), .DIN2(N6752));
hi1s1 U2153 (.Q(N7834), .DIN(N7803));
nnd2s1 U2154 (.Q(N7835), .DIN1(N7803), .DIN2(N6761));
nnd2s1 U2155 (.Q(N7836), .DIN1(N7821), .DIN2(N7807));
nnd2s1 U2156 (.Q(N7839), .DIN1(N7822), .DIN2(N7809));
nnd2s1 U2157 (.Q(N7842), .DIN1(N7823), .DIN2(N7811));
hi1s1 U2158 (.Q(N7845), .DIN(N7812));
nnd2s1 U2159 (.Q(N7846), .DIN1(N7812), .DIN2(N6790));
nnd2s1 U2160 (.Q(N7851), .DIN1(N6298), .DIN2(N7832));
nnd2s1 U2161 (.Q(N7852), .DIN1(N6316), .DIN2(N7834));
nnd2s1 U2162 (.Q(N7859), .DIN1(N6364), .DIN2(N7845));
hi1s1 U2163 (.Q(N7860), .DIN(N7826));
nnd2s1 U2164 (.Q(N7861), .DIN1(N7826), .DIN2(N6741));
hi1s1 U2165 (.Q(N7862), .DIN(N7829));
nnd2s1 U2166 (.Q(N7863), .DIN1(N7829), .DIN2(N6746));
nnd2s1 U2167 (.Q(N7864), .DIN1(N7851), .DIN2(N7833));
nnd2s1 U2168 (.Q(N7867), .DIN1(N7852), .DIN2(N7835));
hi1s1 U2169 (.Q(N7870), .DIN(N7836));
nnd2s1 U2170 (.Q(N7871), .DIN1(N7836), .DIN2(N5730));
hi1s1 U2171 (.Q(N7872), .DIN(N7839));
nnd2s1 U2172 (.Q(N7873), .DIN1(N7839), .DIN2(N5732));
hi1s1 U2173 (.Q(N7874), .DIN(N7842));
nnd2s1 U2174 (.Q(N7875), .DIN1(N7842), .DIN2(N6783));
nnd2s1 U2175 (.Q(N7876), .DIN1(N7859), .DIN2(N7846));
nnd2s1 U2176 (.Q(N7879), .DIN1(N6277), .DIN2(N7860));
nnd2s1 U2177 (.Q(N7880), .DIN1(N6289), .DIN2(N7862));
nnd2s1 U2178 (.Q(N7885), .DIN1(N5199), .DIN2(N7870));
nnd2s1 U2179 (.Q(N7886), .DIN1(N5208), .DIN2(N7872));
nnd2s1 U2180 (.Q(N7887), .DIN1(N6356), .DIN2(N7874));
nnd2s1 U2181 (.Q(N7890), .DIN1(N7879), .DIN2(N7861));
nnd2s1 U2182 (.Q(N7893), .DIN1(N7880), .DIN2(N7863));
hi1s1 U2183 (.Q(N7896), .DIN(N7864));
nnd2s1 U2184 (.Q(N7897), .DIN1(N7864), .DIN2(N6753));
hi1s1 U2185 (.Q(N7898), .DIN(N7867));
nnd2s1 U2186 (.Q(N7899), .DIN1(N7867), .DIN2(N6762));
nnd2s1 U2187 (.Q(N7900), .DIN1(N7885), .DIN2(N7871));
nnd2s1 U2188 (.Q(N7903), .DIN1(N7886), .DIN2(N7873));
nnd2s1 U2189 (.Q(N7906), .DIN1(N7887), .DIN2(N7875));
hi1s1 U2190 (.Q(N7909), .DIN(N7876));
nnd2s1 U2191 (.Q(N7910), .DIN1(N7876), .DIN2(N6791));
nnd2s1 U2192 (.Q(N7917), .DIN1(N6301), .DIN2(N7896));
nnd2s1 U2193 (.Q(N7918), .DIN1(N6319), .DIN2(N7898));
nnd2s1 U2194 (.Q(N7923), .DIN1(N6367), .DIN2(N7909));
hi1s1 U2195 (.Q(N7924), .DIN(N7890));
nnd2s1 U2196 (.Q(N7925), .DIN1(N7890), .DIN2(N6680));
hi1s1 U2197 (.Q(N7926), .DIN(N7893));
nnd2s1 U2198 (.Q(N7927), .DIN1(N7893), .DIN2(N6681));
hi1s1 U2199 (.Q(N7928), .DIN(N7900));
nnd2s1 U2200 (.Q(N7929), .DIN1(N7900), .DIN2(N5690));
hi1s1 U2201 (.Q(N7930), .DIN(N7903));
nnd2s1 U2202 (.Q(N7931), .DIN1(N7903), .DIN2(N5691));
nnd2s1 U2203 (.Q(N7932), .DIN1(N7917), .DIN2(N7897));
nnd2s1 U2204 (.Q(N7935), .DIN1(N7918), .DIN2(N7899));
hi1s1 U2205 (.Q(N7938), .DIN(N7906));
nnd2s1 U2206 (.Q(N7939), .DIN1(N7906), .DIN2(N6784));
nnd2s1 U2207 (.Q(N7940), .DIN1(N7923), .DIN2(N7910));
nnd2s1 U2208 (.Q(N7943), .DIN1(N6280), .DIN2(N7924));
nnd2s1 U2209 (.Q(N7944), .DIN1(N6292), .DIN2(N7926));
nnd2s1 U2210 (.Q(N7945), .DIN1(N5202), .DIN2(N7928));
nnd2s1 U2211 (.Q(N7946), .DIN1(N5211), .DIN2(N7930));
nnd2s1 U2212 (.Q(N7951), .DIN1(N6359), .DIN2(N7938));
nnd2s1 U2213 (.Q(N7954), .DIN1(N7943), .DIN2(N7925));
nnd2s1 U2214 (.Q(N7957), .DIN1(N7944), .DIN2(N7927));
nnd2s1 U2215 (.Q(N7960), .DIN1(N7945), .DIN2(N7929));
nnd2s1 U2216 (.Q(N7963), .DIN1(N7946), .DIN2(N7931));
hi1s1 U2217 (.Q(N7966), .DIN(N7932));
nnd2s1 U2218 (.Q(N7967), .DIN1(N7932), .DIN2(N6754));
hi1s1 U2219 (.Q(N7968), .DIN(N7935));
nnd2s1 U2220 (.Q(N7969), .DIN1(N7935), .DIN2(N6755));
nnd2s1 U2221 (.Q(N7970), .DIN1(N7951), .DIN2(N7939));
hi1s1 U2222 (.Q(N7973), .DIN(N7940));
nnd2s1 U2223 (.Q(N7974), .DIN1(N7940), .DIN2(N6785));
nnd2s1 U2224 (.Q(N7984), .DIN1(N6304), .DIN2(N7966));
nnd2s1 U2225 (.Q(N7985), .DIN1(N6322), .DIN2(N7968));
nnd2s1 U2226 (.Q(N7987), .DIN1(N6370), .DIN2(N7973));
and3s1 U2227 (.Q(N7988), .DIN1(N7957), .DIN2(N6831), .DIN3(N1157));
and3s1 U2228 (.Q(N7989), .DIN1(N7954), .DIN2(N6415), .DIN3(N1157));
and3s1 U2229 (.Q(N7990), .DIN1(N7957), .DIN2(N7041), .DIN3(N566));
and3s1 U2230 (.Q(N7991), .DIN1(N7954), .DIN2(N7177), .DIN3(N566));
hi1s1 U2231 (.Q(N7992), .DIN(N7970));
nnd2s1 U2232 (.Q(N7993), .DIN1(N7970), .DIN2(N6448));
and3s1 U2233 (.Q(N7994), .DIN1(N7963), .DIN2(N6857), .DIN3(N1219));
and3s1 U2234 (.Q(N7995), .DIN1(N7960), .DIN2(N6441), .DIN3(N1219));
and3s1 U2235 (.Q(N7996), .DIN1(N7963), .DIN2(N7065), .DIN3(N583));
and3s1 U2236 (.Q(N7997), .DIN1(N7960), .DIN2(N7182), .DIN3(N583));
nnd2s1 U2237 (.Q(N7998), .DIN1(N7984), .DIN2(N7967));
nnd2s1 U2238 (.Q(N8001), .DIN1(N7985), .DIN2(N7969));
nnd2s1 U2239 (.Q(N8004), .DIN1(N7987), .DIN2(N7974));
nnd2s1 U2240 (.Q(N8009), .DIN1(N6051), .DIN2(N7992));
or4s1 U2241 (.Q(N8013), .DIN1(N7988), .DIN2(N7989), .DIN3(N7990), .DIN4(N7991));
or4s1 U2242 (.Q(N8017), .DIN1(N7994), .DIN2(N7995), .DIN3(N7996), .DIN4(N7997));
hi1s1 U2243 (.Q(N8020), .DIN(N7998));
nnd2s1 U2244 (.Q(N8021), .DIN1(N7998), .DIN2(N6682));
hi1s1 U2245 (.Q(N8022), .DIN(N8001));
nnd2s1 U2246 (.Q(N8023), .DIN1(N8001), .DIN2(N6683));
nnd2s1 U2247 (.Q(N8025), .DIN1(N8009), .DIN2(N7993));
hi1s1 U2248 (.Q(N8026), .DIN(N8004));
nnd2s1 U2249 (.Q(N8027), .DIN1(N8004), .DIN2(N6449));
nnd2s1 U2250 (.Q(N8031), .DIN1(N6307), .DIN2(N8020));
nnd2s1 U2251 (.Q(N8032), .DIN1(N6310), .DIN2(N8022));
hi1s1 U2252 (.Q(N8033), .DIN(N8013));
nnd2s1 U2253 (.Q(N8034), .DIN1(N6054), .DIN2(N8026));
and2s1 U2254 (.Q(N8035), .DIN1(N583), .DIN2(N8025));
hi1s1 U2255 (.Q(N8036), .DIN(N8017));
nnd2s1 U2256 (.Q(N8037), .DIN1(N8031), .DIN2(N8021));
nnd2s1 U2257 (.Q(N8038), .DIN1(N8032), .DIN2(N8023));
nnd2s1 U2258 (.Q(N8039), .DIN1(N8034), .DIN2(N8027));
hi1s1 U2259 (.Q(N8040), .DIN(N8038));
and2s1 U2260 (.Q(N8041), .DIN1(N566), .DIN2(N8037));
hi1s1 U2261 (.Q(N8042), .DIN(N8039));
and2s1 U2262 (.Q(N8043), .DIN1(N8040), .DIN2(N1157));
and2s1 U2263 (.Q(N8044), .DIN1(N8042), .DIN2(N1219));
or2s1 U2264 (.Q(N8045), .DIN1(N8043), .DIN2(N8041));
or2s1 U2265 (.Q(N8048), .DIN1(N8044), .DIN2(N8035));
nnd2s1 U2266 (.Q(N8055), .DIN1(N8045), .DIN2(N8033));
hi1s1 U2267 (.Q(N8056), .DIN(N8045));
nnd2s1 U2268 (.Q(N8057), .DIN1(N8048), .DIN2(N8036));
hi1s1 U2269 (.Q(N8058), .DIN(N8048));
nnd2s1 U2270 (.Q(N8059), .DIN1(N8013), .DIN2(N8056));
nnd2s1 U2271 (.Q(N8060), .DIN1(N8017), .DIN2(N8058));
nnd2s1 U2272 (.Q(N8061), .DIN1(N8055), .DIN2(N8059));
nnd2s1 U2273 (.Q(N8064), .DIN1(N8057), .DIN2(N8060));
and3s1 U2274 (.Q(N8071), .DIN1(N8064), .DIN2(N1777), .DIN3(N3130));
and3s1 U2275 (.Q(N8072), .DIN1(N8061), .DIN2(N1761), .DIN3(N3108));
hi1s1 U2276 (.Q(N8073), .DIN(N8061));
hi1s1 U2277 (.Q(N8074), .DIN(N8064));
or4s1 U2278 (.Q(N8075), .DIN1(N7526), .DIN2(N8071), .DIN3(N3659), .DIN4(N2625));
or4s1 U2279 (.Q(N8076), .DIN1(N7636), .DIN2(N8072), .DIN3(N3661), .DIN4(N2627));
and2s1 U2280 (.Q(N8077), .DIN1(N8073), .DIN2(N1727));
and2s1 U2281 (.Q(N8078), .DIN1(N8074), .DIN2(N1727));
or2s1 U2282 (.Q(N8079), .DIN1(N7530), .DIN2(N8077));
or2s1 U2283 (.Q(N8082), .DIN1(N7479), .DIN2(N8078));
and2s1 U2284 (.Q(N8089), .DIN1(N8079), .DIN2(N3063));
and2s1 U2285 (.Q(N8090), .DIN1(N8082), .DIN2(N3063));
and2s1 U2286 (.Q(N8091), .DIN1(N8079), .DIN2(N3063));
and2s1 U2287 (.Q(N8092), .DIN1(N8082), .DIN2(N3063));
or2s1 U2288 (.Q(N8093), .DIN1(N8089), .DIN2(N3071));
or2s1 U2289 (.Q(N8096), .DIN1(N8090), .DIN2(N3072));
or2s1 U2290 (.Q(N8099), .DIN1(N8091), .DIN2(N3073));
or2s1 U2291 (.Q(N8102), .DIN1(N8092), .DIN2(N3074));
and3s1 U2292 (.Q(N8113), .DIN1(N8102), .DIN2(N2779), .DIN3(N2790));
and3s1 U2293 (.Q(N8114), .DIN1(N8099), .DIN2(N1327), .DIN3(N2790));
and3s1 U2294 (.Q(N8115), .DIN1(N8102), .DIN2(N2801), .DIN3(N2812));
and3s1 U2295 (.Q(N8116), .DIN1(N8099), .DIN2(N1351), .DIN3(N2812));
and3s1 U2296 (.Q(N8117), .DIN1(N8096), .DIN2(N2681), .DIN3(N2692));
and3s1 U2297 (.Q(N8118), .DIN1(N8093), .DIN2(N1185), .DIN3(N2692));
and3s1 U2298 (.Q(N8119), .DIN1(N8096), .DIN2(N2756), .DIN3(N2767));
and3s1 U2299 (.Q(N8120), .DIN1(N8093), .DIN2(N1247), .DIN3(N2767));
or4s1 U2300 (.Q(N8121), .DIN1(N8117), .DIN2(N8118), .DIN3(N3662), .DIN4(N2703));
or4s1 U2301 (.Q(N8122), .DIN1(N8119), .DIN2(N8120), .DIN3(N3663), .DIN4(N2778));
or4s1 U2302 (.Q(N8123), .DIN1(N8113), .DIN2(N8114), .DIN3(N3650), .DIN4(N2614));
or4s1 U2303 (.Q(N8124), .DIN1(N8115), .DIN2(N8116), .DIN3(N3658), .DIN4(N2622));
and2s1 U2304 (.Q(N8125), .DIN1(N8121), .DIN2(N2675));
and2s1 U2305 (.Q(N8126), .DIN1(N8122), .DIN2(N2750));
hi1s1 U2306 (.Q(N8127), .DIN(N8125));
hi1s1 U2307 (.Q(N8128), .DIN(N8126));
  and3s1 troj52_0U1 ( .DIN1(troj52_0n1), .DIN2(troj52_0n2), .DIN3(troj52_0n3), .Q(Trigger_en52_0) );
  and3s1 troj52_0U2 ( .DIN1(N7441), .DIN2(N6180), .DIN3(N7697), .Q(troj52_0n3) );
  nor2s1 troj52_0U3 ( .DIN1(N6935), .DIN2(troj52_0n4), .Q(troj52_0n2) );
  i1s1 troj52_0U4 ( .DIN(N6091), .Q(troj52_0n4) );
  and2s1 troj52_0U5 ( .DIN1(N6172), .DIN2(N6133), .Q(troj52_0n1) );
    xor2s1 trojan52_0  (.DIN1(tempN7709), .DIN2(Trigger_en52_0), .Q(N7709) );

endmodule
