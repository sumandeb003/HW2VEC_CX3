
module s13207 ( CK, g1, g10, g1000, g1006, g1008, g1015, g1016, g1017, g1080, 
        g11, g1193, g1194, g1195, g1196, g1197, g1198, g1201, g1202, g1203, 
        g1205, g1206, g1234, g1246, g1553, g1554, g1724, g1783, g1798, g1804, 
        g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g206, 
        g21, g22, g23, g24, g25, g26, g2662, g27, g28, g2844, g2888, g29, g291, 
        g30, g3077, g3096, g31, g3130, g3159, g3191, g32, g37, g372, g3829, 
        g3854, g3856, g3857, g3859, g3860, g41, g42, g4267, g43, g4316, g4370, 
        g4371, g4372, g4373, g44, g45, g453, g4655, g4657, g4660, g4661, g4663, 
        g4664, g49, g5143, g5164, g534, g5571, g5669, g5678, g5682, g5684, 
        g5687, g5729, g594, g6207, g6212, g6223, g6236, g6269, g6288, g6289, 
        g6290, g6291, g6292, g6293, g6294, g6295, g6296, g6297, g6298, g6299, 
        g6300, g6301, g6302, g6303, g6304, g6305, g6306, g6307, g6308, g633, 
        g634, g635, g6376, g6425, g645, g647, g648, g6648, g6653, g6675, g6849, 
        g6850, g6895, g690, g6909, g694, g698, g702, g7048, g7063, g7103, g722, 
        g723, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, 
        g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, 
        g7505, g7506, g7507, g7508, g751, g7514, g752, g753, g754, g755, g756, 
        g757, g7729, g7730, g7731, g7732, g7763, g781, g785, g786, g795, g8216, 
        g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9, g9128, 
        g9132, g9204, g9280, g929, g9297, g9299, g9305, g9308, g9310, g9312, 
        g9314, g9378, g941, g955, g962, test_se, test_si, test_so );
  input CK, g1, g10, g1000, g1008, g1016, g1080, g11, g1194, g1196, g1198,
         g1202, g1203, g1206, g1234, g1553, g1554, g21, g22, g23, g24, g25,
         g26, g27, g28, g29, g30, g31, g32, g37, g41, g42, g43, g44, g45, g49,
         g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722,
         g723, g751, g752, g753, g754, g755, g756, g757, g781, g786, g795, g9,
         g929, g941, g955, g962, test_se, test_si;
  output g1006, g1015, g1017, g1193, g1195, g1197, g1201, g1205, g1246, g1724,
         g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894,
         g1911, g1944, g206, g2662, g2844, g2888, g291, g3077, g3096, g3130,
         g3159, g3191, g372, g3829, g3854, g3856, g3857, g3859, g3860, g4267,
         g4316, g4370, g4371, g4372, g4373, g453, g4655, g4657, g4660, g4661,
         g4663, g4664, g5143, g5164, g534, g5571, g5669, g5678, g5682, g5684,
         g5687, g5729, g594, g6207, g6212, g6223, g6236, g6269, g6288, g6289,
         g6290, g6291, g6292, g6293, g6294, g6295, g6296, g6297, g6298, g6299,
         g6300, g6301, g6302, g6303, g6304, g6305, g6306, g6307, g6308, g6376,
         g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063,
         g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291,
         g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504,
         g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g7763,
         g785, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958,
         g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312,
         g9314, g9378, test_so;
  wire   g3077, g3860, g5143, g5729, g594, g6269, g6288, g6289, g6290, g6291,
         g6292, g6293, g6294, g6296, g6297, g6298, g6299, g6300, g6301, g6302,
         g6303, g6304, g6305, g6306, g6307, g6308, g6376, g6909, g7504, g7505,
         g7506, g7507, g7508, g7729, g7730, g7731, g7732, g8216, g8217, g8218,
         g8219, g8663, g9132, g9204, g7739, g162, g673, g677, n2119, g146,
         g734, g714, n2039, g706, g855, g665, g859, g150, g661, g158, g2654,
         g669, g685, g174, g681, n1525, g730, g710, g718, n1477, n1480, n1482,
         n1484, n1486, n1488, n1490, n1492, n1494, n1496, n1428, n1502, n1504,
         n1506, n1508, n1511, n1513, n1429, n1412, n1414, n1413, g9389, n1388,
         g9375, g9376, g9374, g9373, g9372, g9360, g9362, g5153, g5154, g5155,
         g5156, \DFF_270/net495 , g179, g5149, \DFF_404/net629 , g180, g5157,
         g5150, g5147, g5151, n1391, g5148, n1409, g5152, g9145, g9134, n1470,
         n1440, g9133, g2653, g9117, g9116, g9115, g9114, g9113, g9112, g9111,
         g9110, g9109, g9108, g9107, g9106, g9105, g9104, g9103, g9102, g9101,
         g9100, g9099, g9098, g9097, g9096, g9095, g9094, g9093, g9092, g9091,
         g9090, g9089, g9088, g9087, g9086, g9085, g9036, g9035, g9034, n1433,
         g9033, g9032, g9031, g9030, g9029, g9028, g9027, g9026, g8960, g8959,
         n1459, g8957, g999, \DFF_160/net385 , g8875, g8874, g8873, g8871,
         g8870, n1446, g8869, n1401, g8867, g8865, g8864, g8678, n1451, g8676,
         n1403, g8675, g8674, n1402, g8673, g8672, g8671, g954, g8670, g953,
         g8669, g952, g8668, g951, g8667, g950, n1386, g8666, g949, g8665,
         g948, n1387, g8664, g944, n1471, g7104, g8227, g8226, g8225, g8224,
         n1460, g973, g7775, n1419, g7774, g7773, g7772, g7771, n1455, g7770,
         g7769, g7768, n1430, g7767, g7766, n1453, g7765, g976, g7762, g7761,
         g7759, g7758, g7757, n1463, g7756, n1431, n1397, n1444, g7733, g7530,
         n1424, g7529, g7528, g7527, n1422, g3851, g7525, n1462, g7524, g7523,
         g7522, n1441, n1461, g7521, g7520, g7519, n1396, n1407, g7518, g7517,
         g7516, n1393, g7515, n1464, g7513, g7512, n1472, g7511, g7510, g7309,
         g93, g7308, g7307, n1473, g98, g7306, g103, g7305, g108, g7304, g3847,
         g3848, g7303, g7302, g3850, g7301, g3852, g3844, g7300, n1400, g7299,
         g7119, n1410, g7118, g113, g7117, g117, g7116, g121, g7115, g125,
         g7114, g129, g7113, g133, g7112, n1449, g7111, g1253, g7110, g7109,
         g7108, g7107, g7106, n1475, g984, g7102, n1469, g12, g7101, n1405,
         n1468, n1417, n1465, g7100, g7099, n1432, g3855, n1423, n1395, n1383,
         n1380, n1421, n1394, n1382, n1379, g6891, g6890, g6889, g6888, g6887,
         g6886, g6885, g6884, g6883, g6882, g6881, g6880, g6879, g6878, g6877,
         g6876, g6875, g6874, g6873, g6872, g6871, g6870, g6869, g6868, g6867,
         g6866, g6865, n1408, g6864, n1411, n1390, g6863, g6862, g6861, n1474,
         g137, g6859, g6858, g6857, g6856, g6855, n1454, g6854, g6853, g6852,
         n1445, \DFF_144/net369 , \DFF_622/net847 , \DFF_381/net606 ,
         \DFF_371/net596 , g1033, g6392, g3845, g3846, g6391, n1420, g6386,
         g6385, \DFF_373/net598 , g6384, g6383, g6382, g1266, g6381, g6380,
         g6379, g6378, g6377, g6372, \DFF_605/net830 , g6371, g6370, g587,
         g6369, g583, g6368, g579, g6367, g566, g6366, g556, g6365, g543,
         g6364, g539, g6363, g535, g595, \DFF_550/net775 , g6362, g517, g6361,
         g516, g6360, g479, g6359, g478, g6358, g477, g6357, g476, g6356, g475,
         g6355, g474, g6354, g458, g6353, g457, g6352, g456, g6351, g455,
         g6350, g454, g533, \DFF_286/net511 , g6349, g436, g6348, g435, g6347,
         g398, g6346, g397, g6345, g396, g6344, g395, g6343, g394, g6342, g393,
         g6341, g377, g6340, g376, g6339, g375, g6338, g374, g6337, g373, g452,
         \DFF_171/net396 , g6336, g355, g6335, g354, g6334, g317, g6333, g316,
         g6332, g315, g6331, g314, g6330, g313, g6329, g312, g6328, g296,
         g6327, g295, g6326, g294, g6325, g293, g6324, g292, g371,
         \DFF_365/net590 , g6323, g274, g6322, g273, g6321, g236, g6320, g235,
         g6319, g234, g6318, g233, g6317, g232, g6316, g231, g6315, g215,
         g6314, g214, g6313, g213, g6312, g212, g6311, g211, g290,
         \DFF_342/net567 , g5746, g5745, g5180, g5744, g5177, g5743, g141,
         g5742, g145, g5740, g5739, g5738, g5737, g5736, g5173, g5735, g5733,
         g5161, g210, g5732, g5160, g205, g5731, g5159, g195, g5730, g5158,
         g186, g5187, g5186, n1415, g5185, n1452, g5184, g5183, g5181, g5182,
         n1458, g5179, n1399, g5178, n1398, g5175, g5174, g5172,
         \DFF_630/net855 , n1456, \DFF_66/net291 , \DFF_517/net742 ,
         \DFF_313/net538 , g5170, g5169, g5168, \DFF_391/net616 , g5167, g5166,
         g5165, g5163, n1457, g4669, g4668, g4665, g4658, \DFF_422/net647 ,
         \DFF_63/net288 , \DFF_412/net637 , \DFF_635/net860 , \DFF_260/net485 ,
         \DFF_24/net249 , \DFF_140/net365 , \DFF_518/net743 , \DFF_527/net752 ,
         \DFF_180/net405 , g4656, g1269, g1268, \DFF_175/net400 ,
         \DFF_98/net323 , g1398, \DFF_218/net443 , g1391, \DFF_402/net627 ,
         g1401, \DFF_252/net477 , g1395, \DFF_377/net602 , \DFF_84/net309 ,
         \DFF_200/net425 , \DFF_314/net539 , \DFF_564/net789 ,
         \DFF_521/net746 , \DFF_101/net326 , \DFF_619/net844 ,
         \DFF_155/net380 , \DFF_597/net822 , \DFF_20/net245 , g6843, g201,
         g4650, g1204, g94, g1311, g1310, g1159, g1393, g1192, g4642, n1384,
         g3863, g2661, g1155, g1154, g1147, g6841, g2673, g4649, g4646, g1157,
         g1390, g1191, g1403, g1402, g1200, g1199, g200, g1396, g2663, g1399,
         g1312, g1153, g1185, g4651, g4639, g4641, g99, g4648, n1385, g1244,
         g4643, g4644, g1270, g1271, g1005, g1004, g4667, g5146, g4640, g2644,
         g1309, g4647, g2659, g4645, g5145, g1404, g890, g199, n1418, g1156,
         n1416, g1014, g1146, g92, g646, g104, g1308, g109, g2672, n1381,
         g1012, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1389, n1392, n1404, n1406,
         n1425, n1426, n1427, n1434, n1435, n1436, n1437, n1438, n1439, n1442,
         n1443, n1447, n1448, n1450, n1466, n1467, n1476, n1478, n1479, n1481,
         n1483, n1485, n1487, n1489, n1491, n1493, n1495, n1497, n1498, n1499,
         n1500, n1501, n1503, n1505, n1507, n1509, n1510, n1512, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638;

wire Trigger_en1_0,  troj1_0n1,  troj1_0n2,  troj1_0n3,  troj1_0n4,  troj1_0n5,  troj1_0n6,  troj1_0n7,  tempg9027,  Trigger_en1_1,  troj1_1n1,  troj1_1n2,  troj1_1n3,  troj1_1n4,  troj1_1n5,  tempg9112;

  assign g7295 = 1'b1;
  assign g7294 = 1'b1;
  assign g7293 = 1'b1;
  assign g7292 = 1'b1;
  assign g7291 = 1'b1;
  assign g7290 = 1'b1;
  assign g7289 = 1'b1;
  assign g7288 = 1'b1;
  assign g7287 = 1'b1;
  assign g7286 = 1'b1;
  assign g7285 = 1'b1;
  assign g7284 = 1'b1;
  assign g7283 = 1'b1;
  assign g8661 = 1'b0;
  assign g1017 = g3077;
  assign g3859 = g3860;
  assign g3829 = g3860;
  assign g5143 = g1554;
  assign g5729 = g49;
  assign g534 = g594;
  assign g453 = g594;
  assign g372 = g594;
  assign g291 = g594;
  assign g206 = g594;
  assign g6269 = g1000;
  assign g6288 = g9;
  assign g6289 = g1;
  assign g6290 = g11;
  assign g6291 = g10;
  assign g6292 = g22;
  assign g6293 = g23;
  assign g6294 = g24;
  assign g6296 = g26;
  assign g6297 = g27;
  assign g6298 = g28;
  assign g6299 = g21;
  assign g6300 = g29;
  assign g6301 = g30;
  assign g6302 = g31;
  assign g6303 = g32;
  assign g6304 = g37;
  assign g6305 = g41;
  assign g6306 = g42;
  assign g6307 = g44;
  assign g6308 = g45;
  assign g6295 = g6376;
  assign g6376 = g25;
  assign g6909 = g1008;
  assign g5669 = g7504;
  assign g5678 = g7505;
  assign g5682 = g7506;
  assign g5684 = g7507;
  assign g5687 = g7508;
  assign g6207 = g7729;
  assign g6212 = g7730;
  assign g6236 = g7731;
  assign g6223 = g7732;
  assign g6648 = g8216;
  assign g6653 = g8217;
  assign g6425 = g8218;
  assign g6675 = g8219;
  assign g7063 = g8663;
  assign g8234 = g9132;
  assign g9128 = g9204;

  nor2s3 U3 ( .DIN1(n893), .DIN2(n894), .Q(n2298) );
  xor2s3 U4 ( .DIN1(n896), .DIN2(n2248), .Q(n2300) );
  nnd2s3 U5 ( .DIN1(n2054), .DIN2(n1465), .Q(n2119) );
  nnd2s3 U6 ( .DIN1(n752), .DIN2(n897), .Q(n2039) );
  nnd3s3 U7 ( .DIN1(n881), .DIN2(n791), .DIN3(n898), .Q(n897) );
  nnd2s3 U8 ( .DIN1(n853), .DIN2(n899), .Q(n1525) );
  nnd4s2 U9 ( .DIN1(n898), .DIN2(g9389), .DIN3(n879), .DIN4(n881), .Q(n899) );
  or2s3 U10 ( .DIN1(g9389), .DIN2(n1388), .Q(g9378) );
  nnd2s3 U11 ( .DIN1(n900), .DIN2(n901), .Q(g9389) );
  nnd2s3 U12 ( .DIN1(n902), .DIN2(n879), .Q(n901) );
  xor2s3 U13 ( .DIN1(n757), .DIN2(n688), .Q(n902) );
  nnd2s3 U14 ( .DIN1(n903), .DIN2(g6307), .Q(n900) );
  xor2s3 U15 ( .DIN1(n904), .DIN2(n905), .Q(n903) );
  xor2s3 U16 ( .DIN1(n906), .DIN2(n907), .Q(n905) );
  xor2s3 U17 ( .DIN1(g9360), .DIN2(g9373), .Q(n907) );
  xor2s3 U18 ( .DIN1(n2296), .DIN2(g9362), .Q(n906) );
  xor2s3 U19 ( .DIN1(n908), .DIN2(n909), .Q(n904) );
  xor2s3 U20 ( .DIN1(g9374), .DIN2(g9375), .Q(n909) );
  xnr2s3 U21 ( .DIN1(g9372), .DIN2(g9376), .Q(n908) );
  or2s3 U22 ( .DIN1(g9376), .DIN2(n1388), .Q(g9314) );
  or5s3 U23 ( .DIN1(n910), .DIN2(n911), .DIN3(n912), .DIN4(n913), .DIN5(n914), 
        .Q(g9376) );
  or5s3 U24 ( .DIN1(n915), .DIN2(n916), .DIN3(n917), .DIN4(n918), .DIN5(n919), 
        .Q(n914) );
  nor2s3 U25 ( .DIN1(n2120), .DIN2(n920), .Q(n918) );
  nor2s3 U26 ( .DIN1(n2017), .DIN2(n921), .Q(n917) );
  nor2s3 U27 ( .DIN1(n2025), .DIN2(n922), .Q(n916) );
  nor2s3 U28 ( .DIN1(n2079), .DIN2(n923), .Q(n915) );
  nnd3s3 U29 ( .DIN1(n924), .DIN2(n925), .DIN3(n926), .Q(n913) );
  or2s3 U30 ( .DIN1(n927), .DIN2(n2106), .Q(n926) );
  nnd2s3 U31 ( .DIN1(n626), .DIN2(n928), .Q(n925) );
  or5s3 U32 ( .DIN1(n929), .DIN2(n930), .DIN3(n931), .DIN4(n932), .DIN5(n933), 
        .Q(n928) );
  nor2s3 U33 ( .DIN1(n2155), .DIN2(n934), .Q(n933) );
  nor2s3 U34 ( .DIN1(n2146), .DIN2(n935), .Q(n932) );
  nor2s3 U35 ( .DIN1(n2252), .DIN2(n936), .Q(n931) );
  nor2s3 U36 ( .DIN1(n1511), .DIN2(n937), .Q(n930) );
  nor2s3 U37 ( .DIN1(n938), .DIN2(n939), .Q(n929) );
  nor5s3 U38 ( .DIN1(n940), .DIN2(n941), .DIN3(n942), .DIN4(n943), .DIN5(n944), 
        .Q(n938) );
  nor2s3 U39 ( .DIN1(n2009), .DIN2(n945), .Q(n944) );
  nor2s3 U40 ( .DIN1(n946), .DIN2(n884), .Q(n942) );
  nor2s3 U42 ( .DIN1(n2186), .DIN2(n948), .Q(n940) );
  nnd2s3 U43 ( .DIN1(n629), .DIN2(n795), .Q(n924) );
  nor2s3 U44 ( .DIN1(n2033), .DIN2(n949), .Q(n912) );
  nor2s3 U45 ( .DIN1(n1987), .DIN2(n950), .Q(n911) );
  nor2s3 U46 ( .DIN1(n2163), .DIN2(n951), .Q(n910) );
  or2s3 U47 ( .DIN1(g9375), .DIN2(n1388), .Q(g9312) );
  nnd2s3 U48 ( .DIN1(n952), .DIN2(n953), .Q(g9375) );
  nor6s3 U49 ( .DIN1(n954), .DIN2(n955), .DIN3(n956), .DIN4(n957), .DIN5(n958), 
        .DIN6(n959), .Q(n953) );
  nor2s3 U50 ( .DIN1(n1989), .DIN2(n950), .Q(n959) );
  nor2s3 U51 ( .DIN1(n2166), .DIN2(n951), .Q(n958) );
  nor2s3 U52 ( .DIN1(n1988), .DIN2(n960), .Q(n957) );
  nor2s3 U53 ( .DIN1(n2041), .DIN2(n961), .Q(n956) );
  nor2s3 U54 ( .DIN1(n962), .DIN2(n963), .Q(n955) );
  nor5s3 U55 ( .DIN1(n964), .DIN2(n965), .DIN3(n966), .DIN4(n967), .DIN5(n968), 
        .Q(n962) );
  nor2s3 U56 ( .DIN1(n1429), .DIN2(n937), .Q(n968) );
  nor2s3 U57 ( .DIN1(n969), .DIN2(n939), .Q(n967) );
  nor5s3 U58 ( .DIN1(n970), .DIN2(n971), .DIN3(n972), .DIN4(n943), .DIN5(n973), 
        .Q(n969) );
  nor2s3 U59 ( .DIN1(n2008), .DIN2(n945), .Q(n973) );
  and2s3 U60 ( .DIN1(n642), .DIN2(g633), .Q(n972) );
  nor2s3 U62 ( .DIN1(n2178), .DIN2(n948), .Q(n970) );
  nor2s3 U63 ( .DIN1(n2251), .DIN2(n936), .Q(n966) );
  nor2s3 U64 ( .DIN1(n2152), .DIN2(n934), .Q(n965) );
  nor2s3 U65 ( .DIN1(n2139), .DIN2(n935), .Q(n964) );
  nor2s3 U66 ( .DIN1(n2107), .DIN2(n927), .Q(n954) );
  nor6s3 U67 ( .DIN1(n974), .DIN2(n975), .DIN3(n976), .DIN4(n919), .DIN5(n977), 
        .DIN6(n978), .Q(n952) );
  nor2s3 U68 ( .DIN1(n2121), .DIN2(n920), .Q(n978) );
  nor2s3 U69 ( .DIN1(n2016), .DIN2(n921), .Q(n977) );
  nor2s3 U70 ( .DIN1(n1990), .DIN2(n923), .Q(n976) );
  nor2s3 U71 ( .DIN1(n2032), .DIN2(n949), .Q(n975) );
  nor2s3 U72 ( .DIN1(n2024), .DIN2(n922), .Q(n974) );
  or2s3 U73 ( .DIN1(g9374), .DIN2(n1388), .Q(g9310) );
  nnd2s3 U74 ( .DIN1(n979), .DIN2(n980), .Q(g9374) );
  nor6s3 U75 ( .DIN1(n981), .DIN2(n982), .DIN3(n983), .DIN4(n984), .DIN5(n985), 
        .DIN6(n986), .Q(n980) );
  nor2s3 U76 ( .DIN1(n1992), .DIN2(n950), .Q(n986) );
  nor2s3 U77 ( .DIN1(n2160), .DIN2(n951), .Q(n985) );
  nor2s3 U78 ( .DIN1(n1991), .DIN2(n960), .Q(n984) );
  nor2s3 U79 ( .DIN1(n2040), .DIN2(n961), .Q(n983) );
  nor2s3 U80 ( .DIN1(n987), .DIN2(n963), .Q(n982) );
  nor5s3 U81 ( .DIN1(n988), .DIN2(n989), .DIN3(n990), .DIN4(n991), .DIN5(n992), 
        .Q(n987) );
  nor2s3 U82 ( .DIN1(n1496), .DIN2(n937), .Q(n992) );
  nor2s3 U83 ( .DIN1(n993), .DIN2(n939), .Q(n991) );
  nor5s3 U84 ( .DIN1(n994), .DIN2(n995), .DIN3(n996), .DIN4(n943), .DIN5(n997), 
        .Q(n993) );
  nor2s3 U85 ( .DIN1(n2007), .DIN2(n945), .Q(n997) );
  and2s3 U86 ( .DIN1(n642), .DIN2(g634), .Q(n996) );
  nor2s3 U88 ( .DIN1(n2179), .DIN2(n948), .Q(n994) );
  nor2s3 U89 ( .DIN1(n2250), .DIN2(n936), .Q(n990) );
  nor2s3 U90 ( .DIN1(n934), .DIN2(n694), .Q(n989) );
  nor2s3 U91 ( .DIN1(n2140), .DIN2(n935), .Q(n988) );
  nor2s3 U92 ( .DIN1(n2108), .DIN2(n927), .Q(n981) );
  nor6s3 U93 ( .DIN1(n998), .DIN2(n999), .DIN3(n1000), .DIN4(n919), .DIN5(
        n1001), .DIN6(n1002), .Q(n979) );
  nor2s3 U94 ( .DIN1(n2122), .DIN2(n920), .Q(n1002) );
  nor2s3 U95 ( .DIN1(n2015), .DIN2(n921), .Q(n1001) );
  nor2s3 U96 ( .DIN1(n2065), .DIN2(n923), .Q(n1000) );
  nor2s3 U97 ( .DIN1(n2031), .DIN2(n949), .Q(n999) );
  nor2s3 U98 ( .DIN1(n2023), .DIN2(n922), .Q(n998) );
  or2s3 U99 ( .DIN1(g9373), .DIN2(n1388), .Q(g9308) );
  or5s3 U100 ( .DIN1(n1003), .DIN2(n1004), .DIN3(n1005), .DIN4(n1006), .DIN5(
        n1007), .Q(g9373) );
  or5s3 U101 ( .DIN1(n1008), .DIN2(n919), .DIN3(n1009), .DIN4(n1010), .DIN5(
        n1011), .Q(n1007) );
  or5s3 U102 ( .DIN1(n1012), .DIN2(n1013), .DIN3(n1014), .DIN4(n1015), .DIN5(
        n1016), .Q(n1011) );
  nor2s3 U103 ( .DIN1(n2123), .DIN2(n920), .Q(n1016) );
  nor2s3 U104 ( .DIN1(n2115), .DIN2(n1017), .Q(n1015) );
  nor2s3 U105 ( .DIN1(n2129), .DIN2(n1018), .Q(n1014) );
  nor2s3 U106 ( .DIN1(n2014), .DIN2(n921), .Q(n1013) );
  nor2s3 U107 ( .DIN1(n2022), .DIN2(n922), .Q(n1012) );
  nor2s3 U108 ( .DIN1(n2247), .DIN2(n1019), .Q(n1010) );
  nor2s3 U109 ( .DIN1(n2234), .DIN2(n1020), .Q(n1009) );
  nor2s3 U110 ( .DIN1(n2221), .DIN2(n1021), .Q(n1008) );
  nnd4s2 U111 ( .DIN1(n1022), .DIN2(n1023), .DIN3(n1024), .DIN4(n1025), .Q(
        n1006) );
  nnd2s3 U112 ( .DIN1(n627), .DIN2(g5156), .Q(n1025) );
  nnd2s3 U113 ( .DIN1(n638), .DIN2(g179), .Q(n1024) );
  nnd2s3 U114 ( .DIN1(n639), .DIN2(n781), .Q(n1023) );
  nnd2s3 U115 ( .DIN1(n636), .DIN2(n840), .Q(n1022) );
  nnd3s3 U116 ( .DIN1(n1026), .DIN2(n1027), .DIN3(n1028), .Q(n1005) );
  or2s3 U117 ( .DIN1(n927), .DIN2(n2109), .Q(n1028) );
  nnd2s3 U118 ( .DIN1(n626), .DIN2(n1029), .Q(n1027) );
  or5s3 U119 ( .DIN1(n1030), .DIN2(n1031), .DIN3(n1032), .DIN4(n1033), .DIN5(
        n1034), .Q(n1029) );
  nor2s3 U120 ( .DIN1(n2153), .DIN2(n934), .Q(n1034) );
  nor2s3 U121 ( .DIN1(n2141), .DIN2(n935), .Q(n1033) );
  nor2s3 U122 ( .DIN1(n2249), .DIN2(n936), .Q(n1032) );
  nor2s3 U123 ( .DIN1(n1412), .DIN2(n937), .Q(n1031) );
  nor2s3 U124 ( .DIN1(n1035), .DIN2(n939), .Q(n1030) );
  nor5s3 U125 ( .DIN1(n1036), .DIN2(n943), .DIN3(n1037), .DIN4(n1038), .DIN5(
        n1039), .Q(n1035) );
  nor2s3 U126 ( .DIN1(n2006), .DIN2(n945), .Q(n1039) );
  nor2s3 U127 ( .DIN1(n2182), .DIN2(n1040), .Q(n1038) );
  nor2s3 U128 ( .DIN1(n1041), .DIN2(n889), .Q(n1037) );
  nnd4s2 U129 ( .DIN1(n1042), .DIN2(n1043), .DIN3(n1044), .DIN4(n1045), .Q(
        n1036) );
  nnd2s3 U130 ( .DIN1(g635), .DIN2(n642), .Q(n1045) );
  nnd2s3 U131 ( .DIN1(n630), .DIN2(n829), .Q(n1044) );
  nnd2s3 U133 ( .DIN1(n1046), .DIN2(n670), .Q(n1042) );
  nnd2s3 U134 ( .DIN1(n629), .DIN2(n720), .Q(n1026) );
  nor2s3 U135 ( .DIN1(n2159), .DIN2(n951), .Q(n1004) );
  nor2s3 U136 ( .DIN1(n1047), .DIN2(\DFF_270/net495 ), .Q(n1003) );
  or2s3 U137 ( .DIN1(g9372), .DIN2(n1388), .Q(g9305) );
  or5s3 U138 ( .DIN1(n1048), .DIN2(n1049), .DIN3(n1050), .DIN4(n1051), .DIN5(
        n1052), .Q(g9372) );
  or5s3 U139 ( .DIN1(n1053), .DIN2(n919), .DIN3(n1054), .DIN4(n1055), .DIN5(
        n1056), .Q(n1052) );
  or5s3 U140 ( .DIN1(n1057), .DIN2(n1058), .DIN3(n1059), .DIN4(n1060), .DIN5(
        n1061), .Q(n1056) );
  nor2s3 U141 ( .DIN1(n2124), .DIN2(n920), .Q(n1061) );
  nor2s3 U142 ( .DIN1(n2114), .DIN2(n1017), .Q(n1060) );
  nor2s3 U143 ( .DIN1(n2128), .DIN2(n1018), .Q(n1059) );
  nor2s3 U144 ( .DIN1(n2013), .DIN2(n921), .Q(n1058) );
  nor2s3 U145 ( .DIN1(n2021), .DIN2(n922), .Q(n1057) );
  nor2s3 U146 ( .DIN1(n2246), .DIN2(n1019), .Q(n1055) );
  nor2s3 U147 ( .DIN1(n2233), .DIN2(n1020), .Q(n1054) );
  nor2s3 U148 ( .DIN1(n2220), .DIN2(n1021), .Q(n1053) );
  nnd4s2 U149 ( .DIN1(n1062), .DIN2(n1063), .DIN3(n1064), .DIN4(n1065), .Q(
        n1051) );
  nnd2s3 U150 ( .DIN1(n627), .DIN2(g5149), .Q(n1065) );
  nnd2s3 U151 ( .DIN1(n638), .DIN2(g180), .Q(n1064) );
  nnd2s3 U152 ( .DIN1(n639), .DIN2(n724), .Q(n1063) );
  or2s3 U153 ( .DIN1(n923), .DIN2(n2278), .Q(n1062) );
  nnd3s3 U154 ( .DIN1(n1066), .DIN2(n1067), .DIN3(n1068), .Q(n1050) );
  or2s3 U155 ( .DIN1(n927), .DIN2(n2110), .Q(n1068) );
  nnd2s3 U156 ( .DIN1(n626), .DIN2(n1069), .Q(n1067) );
  or5s3 U157 ( .DIN1(n1070), .DIN2(n1071), .DIN3(n1072), .DIN4(n1073), .DIN5(
        n1074), .Q(n1069) );
  nor2s3 U158 ( .DIN1(n2148), .DIN2(n934), .Q(n1074) );
  nor2s3 U159 ( .DIN1(n2142), .DIN2(n935), .Q(n1073) );
  nor2s3 U160 ( .DIN1(n2256), .DIN2(n936), .Q(n1072) );
  and2s3 U161 ( .DIN1(n640), .DIN2(n2304), .Q(n1071) );
  nor2s3 U162 ( .DIN1(n1075), .DIN2(n939), .Q(n1070) );
  nor5s3 U163 ( .DIN1(n1076), .DIN2(n943), .DIN3(n1077), .DIN4(n1078), .DIN5(
        n1079), .Q(n1075) );
  nor2s3 U164 ( .DIN1(n2005), .DIN2(n945), .Q(n1079) );
  nor2s3 U165 ( .DIN1(n2184), .DIN2(n1040), .Q(n1078) );
  nor2s3 U166 ( .DIN1(n1041), .DIN2(n888), .Q(n1077) );
  nnd4s2 U167 ( .DIN1(n1080), .DIN2(n1081), .DIN3(n1082), .DIN4(n1083), .Q(
        n1076) );
  nnd2s3 U168 ( .DIN1(g645), .DIN2(n642), .Q(n1083) );
  nnd2s3 U169 ( .DIN1(n630), .DIN2(n675), .Q(n1082) );
  nnd2s3 U171 ( .DIN1(n2306), .DIN2(n647), .Q(n1080) );
  nnd2s3 U172 ( .DIN1(n629), .DIN2(n741), .Q(n1066) );
  nor2s3 U173 ( .DIN1(n2162), .DIN2(n951), .Q(n1049) );
  nor2s3 U174 ( .DIN1(n1047), .DIN2(\DFF_404/net629 ), .Q(n1048) );
  or2s3 U175 ( .DIN1(n2296), .DIN2(n1388), .Q(g9299) );
  nnd2s3 U176 ( .DIN1(n1084), .DIN2(n1085), .Q(n2296) );
  nor6s3 U177 ( .DIN1(n1086), .DIN2(n1087), .DIN3(n1088), .DIN4(n1089), .DIN5(
        n1090), .DIN6(n1091), .Q(n1085) );
  nor2s3 U178 ( .DIN1(n2245), .DIN2(n1019), .Q(n1091) );
  nor2s3 U179 ( .DIN1(n1418), .DIN2(n923), .Q(n1090) );
  nor2s3 U180 ( .DIN1(n2219), .DIN2(n1021), .Q(n1089) );
  nor2s3 U181 ( .DIN1(n1092), .DIN2(n963), .Q(n1088) );
  nor6s3 U182 ( .DIN1(n1093), .DIN2(n1094), .DIN3(n1095), .DIN4(n1096), .DIN5(
        n1097), .DIN6(n1098), .Q(n1092) );
  nor2s3 U183 ( .DIN1(n2143), .DIN2(n935), .Q(n1098) );
  nor2s3 U184 ( .DIN1(n2255), .DIN2(n936), .Q(n1097) );
  nor2s3 U185 ( .DIN1(n2147), .DIN2(n934), .Q(n1096) );
  nor2s3 U186 ( .DIN1(n1099), .DIN2(n939), .Q(n1095) );
  nor5s3 U187 ( .DIN1(n1100), .DIN2(n943), .DIN3(n1101), .DIN4(n1102), .DIN5(
        n1103), .Q(n1099) );
  nor2s3 U188 ( .DIN1(n2004), .DIN2(n945), .Q(n1103) );
  nor2s3 U189 ( .DIN1(n2183), .DIN2(n1040), .Q(n1102) );
  nor2s3 U190 ( .DIN1(n1041), .DIN2(n887), .Q(n1101) );
  nnd4s2 U191 ( .DIN1(n1104), .DIN2(n1105), .DIN3(n1106), .DIN4(n1107), .Q(
        n1100) );
  nnd2s3 U192 ( .DIN1(n642), .DIN2(n810), .Q(n1107) );
  nnd2s3 U193 ( .DIN1(n630), .DIN2(n684), .Q(n1106) );
  nnd2s3 U195 ( .DIN1(n2305), .DIN2(n871), .Q(n1104) );
  nor2s3 U196 ( .DIN1(n2054), .DIN2(n1108), .Q(n1094) );
  nor2s3 U197 ( .DIN1(n1414), .DIN2(n937), .Q(n1093) );
  nor2s3 U198 ( .DIN1(n2168), .DIN2(n1109), .Q(n1087) );
  or5s3 U199 ( .DIN1(n1110), .DIN2(n1111), .DIN3(n1112), .DIN4(n1113), .DIN5(
        n1114), .Q(n1086) );
  nor2s3 U200 ( .DIN1(n2232), .DIN2(n1020), .Q(n1114) );
  nor2s3 U201 ( .DIN1(n2116), .DIN2(n1018), .Q(n1113) );
  nor2s3 U202 ( .DIN1(n1995), .DIN2(n950), .Q(n1112) );
  nor2s3 U203 ( .DIN1(n2157), .DIN2(n951), .Q(n1111) );
  nor2s3 U204 ( .DIN1(n1994), .DIN2(n1047), .Q(n1110) );
  nor6s3 U205 ( .DIN1(n1115), .DIN2(n1116), .DIN3(n1117), .DIN4(n1118), .DIN5(
        n1119), .DIN6(n1120), .Q(n1084) );
  nor2s3 U206 ( .DIN1(n2111), .DIN2(n927), .Q(n1120) );
  nor2s3 U207 ( .DIN1(n2045), .DIN2(n961), .Q(n1119) );
  nor2s3 U208 ( .DIN1(n2012), .DIN2(n921), .Q(n1118) );
  nor2s3 U209 ( .DIN1(n2028), .DIN2(n949), .Q(n1117) );
  nor2s3 U210 ( .DIN1(n1993), .DIN2(n960), .Q(n1116) );
  nnd4s2 U211 ( .DIN1(n792), .DIN2(n1121), .DIN3(n1122), .DIN4(n1123), .Q(
        n1115) );
  or2s3 U212 ( .DIN1(n922), .DIN2(n2020), .Q(n1123) );
  or2s3 U213 ( .DIN1(n1017), .DIN2(n2103), .Q(n1122) );
  or2s3 U214 ( .DIN1(n920), .DIN2(n2125), .Q(n1121) );
  or2s3 U215 ( .DIN1(g9360), .DIN2(n1388), .Q(g9297) );
  nnd2s3 U216 ( .DIN1(n1124), .DIN2(n1125), .Q(g9360) );
  nor6s3 U217 ( .DIN1(n1126), .DIN2(n1127), .DIN3(n1128), .DIN4(n1129), .DIN5(
        n1130), .DIN6(n1131), .Q(n1125) );
  nor2s3 U218 ( .DIN1(n1132), .DIN2(n963), .Q(n1131) );
  nor6s3 U219 ( .DIN1(n1133), .DIN2(n1134), .DIN3(n1135), .DIN4(n1136), .DIN5(
        n1137), .DIN6(n1138), .Q(n1132) );
  nor2s3 U220 ( .DIN1(n2144), .DIN2(n935), .Q(n1138) );
  nor2s3 U221 ( .DIN1(n2254), .DIN2(n936), .Q(n1137) );
  nor2s3 U222 ( .DIN1(n2149), .DIN2(n934), .Q(n1136) );
  nor2s3 U223 ( .DIN1(n1139), .DIN2(n939), .Q(n1135) );
  nor6s3 U224 ( .DIN1(n1140), .DIN2(n1141), .DIN3(n1142), .DIN4(n1143), .DIN5(
        n943), .DIN6(n1144), .Q(n1139) );
  nor2s3 U225 ( .DIN1(n1145), .DIN2(n853), .Q(n1144) );
  nor2s3 U226 ( .DIN1(n1041), .DIN2(n886), .Q(n1143) );
  nor2s3 U227 ( .DIN1(n2011), .DIN2(n945), .Q(n1142) );
  nor2s3 U228 ( .DIN1(n2185), .DIN2(n1040), .Q(n1141) );
  nnd4s2 U229 ( .DIN1(n1146), .DIN2(n1147), .DIN3(n1148), .DIN4(n1149), .Q(
        n1140) );
  nnd2s3 U230 ( .DIN1(g647), .DIN2(n642), .Q(n1149) );
  or2s3 U231 ( .DIN1(n948), .DIN2(n2176), .Q(n1148) );
  nnd2s3 U233 ( .DIN1(n1046), .DIN2(n788), .Q(n1146) );
  nor2s3 U234 ( .DIN1(n1469), .DIN2(n1108), .Q(n1134) );
  nor2s3 U235 ( .DIN1(n1428), .DIN2(n937), .Q(n1133) );
  nor2s3 U236 ( .DIN1(n2170), .DIN2(n1109), .Q(n1130) );
  nor2s3 U237 ( .DIN1(n2044), .DIN2(n961), .Q(n1129) );
  nor2s3 U238 ( .DIN1(n1997), .DIN2(n1047), .Q(n1128) );
  nor2s3 U239 ( .DIN1(n2113), .DIN2(n927), .Q(n1127) );
  or5s3 U240 ( .DIN1(n1150), .DIN2(n1151), .DIN3(n1152), .DIN4(n1153), .DIN5(
        n1154), .Q(n1126) );
  nor2s3 U241 ( .DIN1(n2101), .DIN2(n923), .Q(n1154) );
  nor2s3 U242 ( .DIN1(n2035), .DIN2(n949), .Q(n1153) );
  nor2s3 U243 ( .DIN1(n1999), .DIN2(n960), .Q(n1152) );
  nor2s3 U244 ( .DIN1(n1998), .DIN2(n950), .Q(n1151) );
  nor2s3 U245 ( .DIN1(n2156), .DIN2(n951), .Q(n1150) );
  nor6s3 U246 ( .DIN1(n1155), .DIN2(n1156), .DIN3(n1157), .DIN4(n1158), .DIN5(
        n1159), .DIN6(n1160), .Q(n1124) );
  nor2s3 U247 ( .DIN1(n2019), .DIN2(n921), .Q(n1160) );
  nor2s3 U248 ( .DIN1(n2027), .DIN2(n922), .Q(n1159) );
  nor2s3 U249 ( .DIN1(n2117), .DIN2(n1018), .Q(n1158) );
  nor2s3 U250 ( .DIN1(n2127), .DIN2(n920), .Q(n1157) );
  nor2s3 U251 ( .DIN1(n2104), .DIN2(n1017), .Q(n1156) );
  nnd4s2 U252 ( .DIN1(n792), .DIN2(n1161), .DIN3(n1162), .DIN4(n1163), .Q(
        n1155) );
  nnd2s3 U253 ( .DIN1(n631), .DIN2(n674), .Q(n1163) );
  nnd2s3 U254 ( .DIN1(n634), .DIN2(n828), .Q(n1162) );
  nnd2s3 U255 ( .DIN1(n2307), .DIN2(n842), .Q(n1161) );
  or2s3 U256 ( .DIN1(g9362), .DIN2(n1388), .Q(g9280) );
  nnd2s3 U257 ( .DIN1(n1164), .DIN2(n1165), .Q(g9362) );
  nor6s3 U258 ( .DIN1(n1166), .DIN2(n1167), .DIN3(n1168), .DIN4(n1169), .DIN5(
        n1170), .DIN6(n1171), .Q(n1165) );
  nor2s3 U259 ( .DIN1(n1172), .DIN2(n963), .Q(n1171) );
  or4s3 U260 ( .DIN1(n636), .DIN2(n637), .DIN3(n1173), .DIN4(n1174), .Q(n963)
         );
  or5s3 U261 ( .DIN1(n1175), .DIN2(n632), .DIN3(n638), .DIN4(n628), .DIN5(n635), .Q(n1174) );
  nnd3s3 U262 ( .DIN1(n1047), .DIN2(n950), .DIN3(n1176), .Q(n1173) );
  nor4s3 U263 ( .DIN1(n1177), .DIN2(n1178), .DIN3(n1179), .DIN4(n1180), .Q(
        n1172) );
  nor2s3 U264 ( .DIN1(n1181), .DIN2(n939), .Q(n1180) );
  nnd3s3 U265 ( .DIN1(n1182), .DIN2(n1183), .DIN3(n1184), .Q(n939) );
  nnd2s3 U266 ( .DIN1(n1185), .DIN2(n1391), .Q(n1184) );
  nor6s3 U267 ( .DIN1(n1186), .DIN2(n1187), .DIN3(n1188), .DIN4(n1189), .DIN5(
        n943), .DIN6(n1190), .Q(n1181) );
  nor2s3 U268 ( .DIN1(n1145), .DIN2(n752), .Q(n1190) );
  nor5s3 U269 ( .DIN1(n2305), .DIN2(n947), .DIN3(n643), .DIN4(n641), .DIN5(
        n1191), .Q(n943) );
  nnd4s2 U270 ( .DIN1(n1192), .DIN2(n1040), .DIN3(n946), .DIN4(n948), .Q(n1191) );
  nnd2s3 U271 ( .DIN1(n1193), .DIN2(n1194), .Q(n1192) );
  nnd3s3 U272 ( .DIN1(n1195), .DIN2(n803), .DIN3(n1193), .Q(n1145) );
  nor2s3 U273 ( .DIN1(n1041), .DIN2(n885), .Q(n1189) );
  nnd2s3 U274 ( .DIN1(n1196), .DIN2(n1194), .Q(n1041) );
  nor2s3 U275 ( .DIN1(n2010), .DIN2(n945), .Q(n1188) );
  nor2s3 U276 ( .DIN1(n2187), .DIN2(n1040), .Q(n1187) );
  nnd2s3 U277 ( .DIN1(n1196), .DIN2(n1197), .Q(n1040) );
  nnd4s2 U278 ( .DIN1(n1198), .DIN2(n1199), .DIN3(n1200), .DIN4(n1201), .Q(
        n1186) );
  nnd2s3 U279 ( .DIN1(g648), .DIN2(n642), .Q(n1201) );
  nnd2s3 U280 ( .DIN1(n1196), .DIN2(n1195), .Q(n946) );
  or2s3 U281 ( .DIN1(n948), .DIN2(n2177), .Q(n1200) );
  nnd2s3 U282 ( .DIN1(n1196), .DIN2(n1202), .Q(n948) );
  and2s3 U283 ( .DIN1(n1193), .DIN2(n1409), .Q(n1196) );
  nor5s3 U284 ( .DIN1(n2136), .DIN2(n2137), .DIN3(n2138), .DIN4(n1444), .DIN5(
        n786), .Q(n1193) );
  and4s2 U286 ( .DIN1(n1409), .DIN2(n786), .DIN3(n1197), .DIN4(n1203), .Q(n947) );
  nor4s3 U287 ( .DIN1(n1444), .DIN2(n2138), .DIN3(n2137), .DIN4(n2136), .Q(
        n1203) );
  nnd2s3 U288 ( .DIN1(n2306), .DIN2(n820), .Q(n1198) );
  nor2s3 U289 ( .DIN1(n2145), .DIN2(n935), .Q(n1179) );
  nnd2s3 U290 ( .DIN1(n713), .DIN2(n1195), .Q(n935) );
  nor2s3 U291 ( .DIN1(n2150), .DIN2(n934), .Q(n1178) );
  nnd2s3 U292 ( .DIN1(n1202), .DIN2(n712), .Q(n934) );
  nnd4s2 U293 ( .DIN1(n1204), .DIN2(n1205), .DIN3(n1206), .DIN4(n1207), .Q(
        n1177) );
  nnd3s3 U294 ( .DIN1(n1197), .DIN2(n836), .DIN3(n712), .Q(n1207) );
  or2s3 U295 ( .DIN1(n1108), .DIN2(n1471), .Q(n1206) );
  nnd2s3 U296 ( .DIN1(n713), .DIN2(n1202), .Q(n1108) );
  nnd2s3 U297 ( .DIN1(n1208), .DIN2(n786), .Q(n1182) );
  nnd2s3 U298 ( .DIN1(n640), .DIN2(n860), .Q(n1205) );
  nnd2s3 U299 ( .DIN1(n641), .DIN2(n1391), .Q(n937) );
  nnd2s3 U300 ( .DIN1(n1185), .DIN2(n1195), .Q(n945) );
  or2s3 U301 ( .DIN1(n936), .DIN2(n2253), .Q(n1204) );
  nnd2s3 U302 ( .DIN1(n1185), .DIN2(n1202), .Q(n936) );
  nor2s3 U303 ( .DIN1(n2165), .DIN2(n1109), .Q(n1170) );
  nnd2s3 U304 ( .DIN1(n1194), .DIN2(n712), .Q(n1109) );
  nor2s3 U305 ( .DIN1(n2043), .DIN2(n961), .Q(n1169) );
  nnd2s3 U306 ( .DIN1(n711), .DIN2(n1202), .Q(n961) );
  nor2s3 U307 ( .DIN1(n2000), .DIN2(n1047), .Q(n1168) );
  nnd2s3 U308 ( .DIN1(n1197), .DIN2(n1209), .Q(n1047) );
  nor2s3 U309 ( .DIN1(n2112), .DIN2(n927), .Q(n1167) );
  nnd2s3 U310 ( .DIN1(n1210), .DIN2(n1202), .Q(n927) );
  or5s3 U311 ( .DIN1(n1211), .DIN2(n1212), .DIN3(n1213), .DIN4(n1214), .DIN5(
        n1215), .Q(n1166) );
  nor2s3 U312 ( .DIN1(n2003), .DIN2(n923), .Q(n1215) );
  nnd2s3 U313 ( .DIN1(n1194), .DIN2(n1209), .Q(n923) );
  nor2s3 U314 ( .DIN1(n2034), .DIN2(n949), .Q(n1214) );
  nnd2s3 U315 ( .DIN1(n1175), .DIN2(n1195), .Q(n949) );
  nor2s3 U316 ( .DIN1(n2002), .DIN2(n960), .Q(n1213) );
  nnd2s3 U317 ( .DIN1(n1195), .DIN2(n1209), .Q(n960) );
  nor2s3 U318 ( .DIN1(n2001), .DIN2(n950), .Q(n1212) );
  nnd2s3 U319 ( .DIN1(n1202), .DIN2(n1209), .Q(n950) );
  and3s3 U320 ( .DIN1(n1391), .DIN2(n1216), .DIN3(n1409), .Q(n1209) );
  nor2s3 U321 ( .DIN1(n2158), .DIN2(n951), .Q(n1211) );
  nnd2s3 U322 ( .DIN1(n1195), .DIN2(n712), .Q(n951) );
  nnd2s3 U323 ( .DIN1(n1208), .DIN2(n1391), .Q(n1183) );
  and3s3 U324 ( .DIN1(n1217), .DIN2(n866), .DIN3(n1409), .Q(n1208) );
  nor6s3 U325 ( .DIN1(n1218), .DIN2(n1219), .DIN3(n1220), .DIN4(n1221), .DIN5(
        n1222), .DIN6(n1223), .Q(n1164) );
  nor2s3 U326 ( .DIN1(n2018), .DIN2(n921), .Q(n1223) );
  nnd2s3 U327 ( .DIN1(n711), .DIN2(n1195), .Q(n921) );
  nor2s3 U328 ( .DIN1(n2026), .DIN2(n922), .Q(n1222) );
  nnd2s3 U329 ( .DIN1(n1175), .DIN2(n1202), .Q(n922) );
  nor2s3 U330 ( .DIN1(n1397), .DIN2(n1431), .Q(n1202) );
  nor2s3 U331 ( .DIN1(n2118), .DIN2(n1018), .Q(n1221) );
  nnd2s3 U332 ( .DIN1(n1194), .DIN2(n1210), .Q(n1018) );
  nor2s3 U333 ( .DIN1(n2126), .DIN2(n920), .Q(n1220) );
  nnd2s3 U334 ( .DIN1(n1210), .DIN2(n1195), .Q(n920) );
  nor2s3 U335 ( .DIN1(n644), .DIN2(n1397), .Q(n1195) );
  nor2s3 U336 ( .DIN1(n2105), .DIN2(n1017), .Q(n1219) );
  nnd2s3 U337 ( .DIN1(n1210), .DIN2(n1197), .Q(n1017) );
  and3s3 U338 ( .DIN1(n786), .DIN2(n803), .DIN3(n1216), .Q(n1210) );
  nnd4s2 U339 ( .DIN1(n792), .DIN2(n1224), .DIN3(n1225), .DIN4(n1226), .Q(
        n1218) );
  nnd2s3 U340 ( .DIN1(n631), .DIN2(n807), .Q(n1226) );
  nnd2s3 U341 ( .DIN1(n634), .DIN2(n753), .Q(n1225) );
  nnd2s3 U342 ( .DIN1(n2307), .DIN2(n848), .Q(n1224) );
  nnd2s3 U343 ( .DIN1(n1227), .DIN2(n1228), .Q(g9204) );
  nnd2s3 U344 ( .DIN1(g6303), .DIN2(g6301), .Q(n1228) );
  nnd2s3 U345 ( .DIN1(g6302), .DIN2(n877), .Q(n1227) );
  nnd2s3 U346 ( .DIN1(n1229), .DIN2(n1230), .Q(g9145) );
  nnd2s3 U347 ( .DIN1(n1231), .DIN2(n743), .Q(n1230) );
  nnd2s3 U348 ( .DIN1(n678), .DIN2(n745), .Q(n1229) );
  nnd2s3 U349 ( .DIN1(n1232), .DIN2(n1233), .Q(g9134) );
  nnd2s3 U350 ( .DIN1(n1234), .DIN2(n743), .Q(n1233) );
  nnd2s3 U351 ( .DIN1(n654), .DIN2(n1235), .Q(n1234) );
  nnd2s3 U352 ( .DIN1(n1440), .DIN2(n1236), .Q(n1235) );
  nnd2s3 U353 ( .DIN1(n1470), .DIN2(n1231), .Q(n1232) );
  nor2s3 U355 ( .DIN1(n1239), .DIN2(n778), .Q(g9133) );
  nnd2s3 U356 ( .DIN1(n1240), .DIN2(n1241), .Q(g9117) );
  nnd2s3 U358 ( .DIN1(n1237), .DIN2(n730), .Q(n1240) );
  nnd2s3 U359 ( .DIN1(n1243), .DIN2(n1244), .Q(g9116) );
  nnd2s3 U360 ( .DIN1(n2305), .DIN2(n727), .Q(n1244) );
  or2s3 U361 ( .DIN1(n2306), .DIN2(n2004), .Q(n1243) );
  nnd2s3 U362 ( .DIN1(n1245), .DIN2(n1246), .Q(g9115) );
  nnd2s3 U363 ( .DIN1(n1046), .DIN2(n749), .Q(n1246) );
  or2s3 U364 ( .DIN1(n2305), .DIN2(n2005), .Q(n1245) );
  nnd2s3 U365 ( .DIN1(n1247), .DIN2(n1248), .Q(g9114) );
  nnd2s3 U366 ( .DIN1(n2306), .DIN2(n721), .Q(n1248) );
  or2s3 U367 ( .DIN1(n1046), .DIN2(n2006), .Q(n1247) );
  nnd2s3 U368 ( .DIN1(n1249), .DIN2(n1250), .Q(g9113) );
  nnd2s3 U369 ( .DIN1(n2305), .DIN2(n821), .Q(n1250) );
  or2s3 U370 ( .DIN1(n2306), .DIN2(n2007), .Q(n1249) );
  nnd2s3 U371 ( .DIN1(n1251), .DIN2(n1252), .Q( tempg9112 ) );
  nnd2s3 U372 ( .DIN1(n1046), .DIN2(n857), .Q(n1252) );
  or2s3 U373 ( .DIN1(n2305), .DIN2(n2008), .Q(n1251) );
  nnd2s3 U374 ( .DIN1(n1253), .DIN2(n1254), .Q(g9111) );
  nnd2s3 U375 ( .DIN1(n2306), .DIN2(n835), .Q(n1254) );
  or2s3 U376 ( .DIN1(n1046), .DIN2(n2009), .Q(n1253) );
  nnd2s3 U377 ( .DIN1(n1255), .DIN2(n1256), .Q(g9110) );
  nnd2s3 U378 ( .DIN1(n2305), .DIN2(n686), .Q(n1256) );
  or2s3 U379 ( .DIN1(n2306), .DIN2(n2010), .Q(n1255) );
  nnd2s3 U380 ( .DIN1(n1257), .DIN2(n1258), .Q(g9109) );
  nnd2s3 U381 ( .DIN1(n1046), .DIN2(n800), .Q(n1258) );
  or2s3 U382 ( .DIN1(n2306), .DIN2(n2011), .Q(n1257) );
  and3s3 U383 ( .DIN1(n1259), .DIN2(n786), .DIN3(n1185), .Q(n1046) );
  and3s3 U384 ( .DIN1(n803), .DIN2(n866), .DIN3(n1217), .Q(n1185) );
  nnd2s3 U385 ( .DIN1(n1260), .DIN2(n1261), .Q(g9108) );
  nnd2s3 U386 ( .DIN1(n2307), .DIN2(n676), .Q(n1261) );
  or2s3 U387 ( .DIN1(n2309), .DIN2(n2012), .Q(n1260) );
  nnd2s3 U388 ( .DIN1(n1262), .DIN2(n1263), .Q(g9107) );
  nnd2s3 U389 ( .DIN1(n2307), .DIN2(n672), .Q(n1263) );
  or2s3 U390 ( .DIN1(n2309), .DIN2(n2013), .Q(n1262) );
  nnd2s3 U391 ( .DIN1(n1264), .DIN2(n1265), .Q(g9106) );
  nnd2s3 U392 ( .DIN1(n2307), .DIN2(n718), .Q(n1265) );
  or2s3 U393 ( .DIN1(n2308), .DIN2(n2014), .Q(n1264) );
  nnd2s3 U394 ( .DIN1(n1266), .DIN2(n1267), .Q(g9105) );
  nnd2s3 U395 ( .DIN1(n2307), .DIN2(n798), .Q(n1267) );
  or2s3 U396 ( .DIN1(n2308), .DIN2(n2015), .Q(n1266) );
  nnd2s3 U397 ( .DIN1(n1268), .DIN2(n1269), .Q(g9104) );
  nnd2s3 U398 ( .DIN1(n2307), .DIN2(n815), .Q(n1269) );
  or2s3 U399 ( .DIN1(n2308), .DIN2(n2016), .Q(n1268) );
  nnd2s3 U400 ( .DIN1(n1270), .DIN2(n1271), .Q(g9103) );
  nnd2s3 U401 ( .DIN1(n2307), .DIN2(n740), .Q(n1271) );
  or2s3 U402 ( .DIN1(n2308), .DIN2(n2017), .Q(n1270) );
  nnd2s3 U403 ( .DIN1(n1272), .DIN2(n1273), .Q(g9102) );
  nnd2s3 U404 ( .DIN1(n2307), .DIN2(n715), .Q(n1273) );
  or2s3 U405 ( .DIN1(n2308), .DIN2(n2018), .Q(n1272) );
  nnd2s3 U406 ( .DIN1(n1274), .DIN2(n1275), .Q(g9101) );
  nnd2s3 U407 ( .DIN1(n2307), .DIN2(n847), .Q(n1275) );
  or2s3 U408 ( .DIN1(n2308), .DIN2(n2019), .Q(n1274) );
  nnd2s3 U409 ( .DIN1(n1276), .DIN2(n1277), .Q(g9100) );
  nnd2s3 U410 ( .DIN1(n631), .DIN2(n811), .Q(n1277) );
  or2s3 U411 ( .DIN1(n631), .DIN2(n2020), .Q(n1276) );
  nnd2s3 U412 ( .DIN1(n1278), .DIN2(n1279), .Q(g9099) );
  nnd2s3 U413 ( .DIN1(n631), .DIN2(n782), .Q(n1279) );
  or2s3 U414 ( .DIN1(n631), .DIN2(n2021), .Q(n1278) );
  nnd2s3 U415 ( .DIN1(n1280), .DIN2(n1281), .Q(g9098) );
  nnd2s3 U416 ( .DIN1(n631), .DIN2(n852), .Q(n1281) );
  or2s3 U417 ( .DIN1(n631), .DIN2(n2022), .Q(n1280) );
  nnd2s3 U418 ( .DIN1(n1282), .DIN2(n1283), .Q(g9097) );
  nnd2s3 U419 ( .DIN1(n631), .DIN2(n680), .Q(n1283) );
  or2s3 U420 ( .DIN1(n631), .DIN2(n2023), .Q(n1282) );
  nnd2s3 U421 ( .DIN1(n1284), .DIN2(n1285), .Q(g9096) );
  nnd2s3 U422 ( .DIN1(n631), .DIN2(n677), .Q(n1285) );
  or2s3 U423 ( .DIN1(n631), .DIN2(n2024), .Q(n1284) );
  nnd2s3 U424 ( .DIN1(n1286), .DIN2(n1287), .Q(g9095) );
  nnd2s3 U425 ( .DIN1(n631), .DIN2(n785), .Q(n1287) );
  or2s3 U426 ( .DIN1(n631), .DIN2(n2025), .Q(n1286) );
  nnd2s3 U427 ( .DIN1(n1288), .DIN2(n1289), .Q(g9094) );
  nnd2s3 U428 ( .DIN1(n631), .DIN2(n873), .Q(n1289) );
  or2s3 U429 ( .DIN1(n631), .DIN2(n2026), .Q(n1288) );
  nnd2s3 U430 ( .DIN1(n1290), .DIN2(n1291), .Q(g9093) );
  nnd2s3 U431 ( .DIN1(n631), .DIN2(n748), .Q(n1291) );
  or2s3 U432 ( .DIN1(n631), .DIN2(n2027), .Q(n1290) );
  nnd3s3 U433 ( .DIN1(n1175), .DIN2(n1197), .DIN3(n792), .Q(n1020) );
  nor2s3 U434 ( .DIN1(n780), .DIN2(n1431), .Q(n1197) );
  nnd2s3 U435 ( .DIN1(n1292), .DIN2(n1293), .Q(g9092) );
  nnd2s3 U436 ( .DIN1(n634), .DIN2(n783), .Q(n1293) );
  or2s3 U437 ( .DIN1(n634), .DIN2(n2028), .Q(n1292) );
  nnd2s3 U438 ( .DIN1(n1294), .DIN2(n1295), .Q(g9091) );
  nnd2s3 U439 ( .DIN1(n634), .DIN2(n738), .Q(n1295) );
  nnd2s3 U440 ( .DIN1(n1019), .DIN2(n724), .Q(n1294) );
  nnd2s3 U441 ( .DIN1(n1296), .DIN2(n1297), .Q(g9090) );
  nnd2s3 U442 ( .DIN1(n634), .DIN2(n833), .Q(n1297) );
  nnd2s3 U443 ( .DIN1(n1019), .DIN2(n781), .Q(n1296) );
  nnd2s3 U444 ( .DIN1(n1298), .DIN2(n1299), .Q(g9089) );
  nnd2s3 U445 ( .DIN1(n634), .DIN2(n868), .Q(n1299) );
  or2s3 U446 ( .DIN1(n634), .DIN2(n2031), .Q(n1298) );
  nnd2s3 U447 ( .DIN1(n1300), .DIN2(n1301), .Q(g9088) );
  nnd2s3 U448 ( .DIN1(n634), .DIN2(n844), .Q(n1301) );
  or2s3 U449 ( .DIN1(n634), .DIN2(n2032), .Q(n1300) );
  nnd2s3 U450 ( .DIN1(n1302), .DIN2(n1303), .Q(g9087) );
  nnd2s3 U451 ( .DIN1(n634), .DIN2(n754), .Q(n1303) );
  or2s3 U452 ( .DIN1(n634), .DIN2(n2033), .Q(n1302) );
  nnd2s3 U453 ( .DIN1(n1304), .DIN2(n1305), .Q(g9086) );
  nnd2s3 U454 ( .DIN1(n634), .DIN2(n862), .Q(n1305) );
  or2s3 U455 ( .DIN1(n634), .DIN2(n2034), .Q(n1304) );
  nnd2s3 U456 ( .DIN1(n1306), .DIN2(n1307), .Q(g9085) );
  nnd2s3 U457 ( .DIN1(n634), .DIN2(n710), .Q(n1307) );
  or2s3 U458 ( .DIN1(n634), .DIN2(n2035), .Q(n1306) );
  nnd2s3 U459 ( .DIN1(n1259), .DIN2(n1175), .Q(n1019) );
  and3s3 U460 ( .DIN1(n1216), .DIN2(n786), .DIN3(n1409), .Q(n1175) );
  nor2s3 U461 ( .DIN1(n1308), .DIN2(n1309), .Q(g9036) );
  xnr2s3 U462 ( .DIN1(n2061), .DIN2(n1310), .Q(n1309) );
  nnd2s3 U463 ( .DIN1(n1311), .DIN2(n1312), .Q(g9035) );
  nnd2s3 U465 ( .DIN1(n1237), .DIN2(n706), .Q(n1311) );
  nnd2s3 U466 ( .DIN1(n1313), .DIN2(n1314), .Q(n1237) );
  nnd2s3 U467 ( .DIN1(n1242), .DIN2(n1236), .Q(n1314) );
  nnd3s3 U468 ( .DIN1(n683), .DIN2(n706), .DIN3(n656), .Q(n1242) );
  and2s3 U469 ( .DIN1(n1315), .DIN2(n1316), .Q(g9034) );
  nnd3s3 U470 ( .DIN1(n1317), .DIN2(g9132), .DIN3(n664), .Q(n1315) );
  nnd3s3 U471 ( .DIN1(n2049), .DIN2(n823), .DIN3(n2048), .Q(n1317) );
  nnd2s3 U472 ( .DIN1(n1319), .DIN2(n1320), .Q(g9033) );
  nnd2s3 U473 ( .DIN1(n2307), .DIN2(n770), .Q(n1320) );
  nnd2s3 U474 ( .DIN1(n1021), .DIN2(n741), .Q(n1319) );
  nnd2s3 U475 ( .DIN1(n1321), .DIN2(n1322), .Q(g9032) );
  nnd2s3 U476 ( .DIN1(n2307), .DIN2(n681), .Q(n1322) );
  nnd2s3 U477 ( .DIN1(n1021), .DIN2(n720), .Q(n1321) );
  nnd2s3 U478 ( .DIN1(n1323), .DIN2(n1324), .Q(g9031) );
  nnd2s3 U479 ( .DIN1(n2307), .DIN2(n817), .Q(n1324) );
  or2s3 U480 ( .DIN1(n2308), .DIN2(n2040), .Q(n1323) );
  nnd2s3 U481 ( .DIN1(n1325), .DIN2(n1326), .Q(g9030) );
  nnd2s3 U482 ( .DIN1(n2308), .DIN2(n812), .Q(n1326) );
  or2s3 U483 ( .DIN1(n2308), .DIN2(n2041), .Q(n1325) );
  nnd2s3 U484 ( .DIN1(n1327), .DIN2(n1328), .Q(g9029) );
  nnd2s3 U485 ( .DIN1(n2308), .DIN2(n806), .Q(n1328) );
  nnd2s3 U486 ( .DIN1(n1021), .DIN2(n795), .Q(n1327) );
  nnd2s3 U487 ( .DIN1(n1329), .DIN2(n1330), .Q(g9028) );
  nnd2s3 U488 ( .DIN1(n2308), .DIN2(n789), .Q(n1330) );
  or2s3 U489 ( .DIN1(n2308), .DIN2(n2043), .Q(n1329) );
  nnd2s3 U490 ( .DIN1(n1331), .DIN2(n1332), .Q( tempg9027 ) );
  nnd2s3 U491 ( .DIN1(n2308), .DIN2(n697), .Q(n1332) );
  or2s3 U492 ( .DIN1(n2309), .DIN2(n2044), .Q(n1331) );
  nnd2s3 U493 ( .DIN1(n1333), .DIN2(n1334), .Q(g9026) );
  nnd2s3 U494 ( .DIN1(n2308), .DIN2(n779), .Q(n1334) );
  or2s3 U495 ( .DIN1(n2309), .DIN2(n2045), .Q(n1333) );
  nnd2s3 U496 ( .DIN1(n711), .DIN2(n1259), .Q(n1021) );
  and2s3 U497 ( .DIN1(n792), .DIN2(n1194), .Q(n1259) );
  nor2s3 U498 ( .DIN1(n644), .DIN2(n780), .Q(n1194) );
  nnd3s3 U499 ( .DIN1(n1216), .DIN2(n803), .DIN3(n1391), .Q(n1176) );
  and2s3 U500 ( .DIN1(n1444), .DIN2(n1217), .Q(n1216) );
  and3s3 U501 ( .DIN1(n2137), .DIN2(n2138), .DIN3(n2136), .Q(n1217) );
  and3s3 U502 ( .DIN1(n1335), .DIN2(n1310), .DIN3(n649), .Q(g8960) );
  or2s3 U503 ( .DIN1(n1336), .DIN2(n2058), .Q(n1310) );
  nnd2s3 U504 ( .DIN1(n2058), .DIN2(n1336), .Q(n1335) );
  nnd2s3 U505 ( .DIN1(n1337), .DIN2(n1338), .Q(g8959) );
  nnd2s3 U507 ( .DIN1(n1340), .DIN2(n683), .Q(n1337) );
  nnd2s3 U508 ( .DIN1(g6289), .DIN2(n1341), .Q(g8958) );
  nnd3s3 U509 ( .DIN1(n1342), .DIN2(n831), .DIN3(n1343), .Q(n1341) );
  nnd2s3 U510 ( .DIN1(n876), .DIN2(g9132), .Q(n1342) );
  nor2s3 U511 ( .DIN1(n652), .DIN2(n1344), .Q(g8957) );
  nor2s3 U512 ( .DIN1(n797), .DIN2(n1318), .Q(n1344) );
  or3s3 U513 ( .DIN1(n666), .DIN2(n1345), .DIN3(n1346), .Q(n1318) );
  nor4s3 U514 ( .DIN1(g6269), .DIN2(g6289), .DIN3(n2050), .DIN4(n695), .Q(
        n1346) );
  nor6s3 U515 ( .DIN1(g6850), .DIN2(g6909), .DIN3(g1016), .DIN4(
        \DFF_160/net385 ), .DIN5(n875), .DIN6(n876), .Q(n1345) );
  and2s3 U516 ( .DIN1(n649), .DIN2(n1348), .Q(g8875) );
  nnd2s3 U517 ( .DIN1(n1349), .DIN2(n1350), .Q(n1348) );
  nnd3s3 U518 ( .DIN1(n1351), .DIN2(n751), .DIN3(n2064), .Q(n1350) );
  nnd2s3 U519 ( .DIN1(n1336), .DIN2(n822), .Q(n1349) );
  nnd3s3 U520 ( .DIN1(n822), .DIN2(n751), .DIN3(n1351), .Q(n1336) );
  nor2s3 U521 ( .DIN1(n722), .DIN2(n1352), .Q(g8874) );
  xnr2s3 U522 ( .DIN1(n2072), .DIN2(n1353), .Q(n1352) );
  nnd2s3 U523 ( .DIN1(n1354), .DIN2(n1355), .Q(g8873) );
  nnd2s3 U525 ( .DIN1(n1340), .DIN2(n784), .Q(n1354) );
  nnd2s3 U526 ( .DIN1(n1313), .DIN2(n1356), .Q(n1340) );
  nnd2s3 U527 ( .DIN1(n1339), .DIN2(n1236), .Q(n1356) );
  nnd2s3 U528 ( .DIN1(n657), .DIN2(n784), .Q(n1339) );
  nnd2s3 U529 ( .DIN1(g6289), .DIN2(n1358), .Q(g8872) );
  nnd2s3 U530 ( .DIN1(n1343), .DIN2(n831), .Q(n1358) );
  nnd2s3 U531 ( .DIN1(n1359), .DIN2(n1360), .Q(g8871) );
  nnd3s3 U532 ( .DIN1(n1361), .DIN2(n841), .DIN3(n1362), .Q(n1360) );
  and3s3 U533 ( .DIN1(n1446), .DIN2(n1363), .DIN3(n1362), .Q(g8870) );
  nnd2s3 U534 ( .DIN1(n1361), .DIN2(n1364), .Q(n1363) );
  or2s3 U535 ( .DIN1(n1433), .DIN2(n2049), .Q(n1364) );
  nnd2s3 U536 ( .DIN1(n1359), .DIN2(n1365), .Q(g8869) );
  nnd2s3 U537 ( .DIN1(n1362), .DIN2(n1433), .Q(n1365) );
  and3s3 U538 ( .DIN1(n1366), .DIN2(g43), .DIN3(n1367), .Q(n1362) );
  or2s3 U539 ( .DIN1(n1361), .DIN2(n841), .Q(n1367) );
  nnd2s3 U540 ( .DIN1(n1433), .DIN2(n2049), .Q(n1361) );
  nnd3s3 U541 ( .DIN1(g43), .DIN2(n851), .DIN3(n1366), .Q(n1359) );
  nnd2s3 U542 ( .DIN1(n1401), .DIN2(g9132), .Q(n1366) );
  nor5s3 U543 ( .DIN1(n1368), .DIN2(n1369), .DIN3(n876), .DIN4(n2052), .DIN5(
        n875), .Q(g8867) );
  nor4s3 U544 ( .DIN1(n1368), .DIN2(g6269), .DIN3(g6289), .DIN4(n2050), .Q(
        g8865) );
  and2s3 U545 ( .DIN1(g43), .DIN2(g7298), .Q(g8864) );
  nor2s3 U546 ( .DIN1(n1308), .DIN2(n1370), .Q(g8678) );
  xor2s3 U547 ( .DIN1(n2063), .DIN2(n1351), .Q(n1370) );
  nor2s3 U548 ( .DIN1(n1371), .DIN2(n1451), .Q(n1351) );
  nor2s3 U549 ( .DIN1(n1403), .DIN2(n1372), .Q(g8676) );
  xnr2s3 U550 ( .DIN1(n2167), .DIN2(n1373), .Q(n1372) );
  and3s3 U551 ( .DIN1(n1373), .DIN2(n830), .DIN3(n1374), .Q(g8675) );
  nnd2s3 U552 ( .DIN1(n2169), .DIN2(n1375), .Q(n1374) );
  or2s3 U553 ( .DIN1(n1375), .DIN2(n2169), .Q(n1373) );
  nnd3s3 U554 ( .DIN1(n1376), .DIN2(n1377), .DIN3(n1402), .Q(g8674) );
  nnd4s2 U555 ( .DIN1(n690), .DIN2(n1378), .DIN3(n685), .DIN4(n729), .Q(n1377)
         );
  nnd2s3 U556 ( .DIN1(n1353), .DIN2(n809), .Q(n1376) );
  or2s3 U557 ( .DIN1(n1378), .DIN2(n2134), .Q(n1353) );
  nnd2s3 U558 ( .DIN1(n1389), .DIN2(n1392), .Q(g8673) );
  nnd2s3 U560 ( .DIN1(n1404), .DIN2(n846), .Q(n1389) );
  nnd2s3 U561 ( .DIN1(n1313), .DIN2(n1406), .Q(n1404) );
  nnd2s3 U562 ( .DIN1(n1357), .DIN2(n1236), .Q(n1406) );
  nnd3s3 U563 ( .DIN1(n838), .DIN2(n846), .DIN3(n658), .Q(n1357) );
  and2s3 U564 ( .DIN1(g43), .DIN2(g7103), .Q(g8672) );
  nnd2s3 U565 ( .DIN1(n1425), .DIN2(n1426), .Q(g8671) );
  nnd2s3 U566 ( .DIN1(n1427), .DIN2(g954), .Q(n1426) );
  nnd2s3 U567 ( .DIN1(n736), .DIN2(n860), .Q(n1425) );
  nnd2s3 U568 ( .DIN1(n1434), .DIN2(n1435), .Q(g8670) );
  nnd2s3 U569 ( .DIN1(n1427), .DIN2(g953), .Q(n1435) );
  nnd2s3 U570 ( .DIN1(n736), .DIN2(n843), .Q(n1434) );
  nnd2s3 U571 ( .DIN1(n1436), .DIN2(n1437), .Q(g8669) );
  nnd2s3 U572 ( .DIN1(n1427), .DIN2(g952), .Q(n1437) );
  nnd2s3 U573 ( .DIN1(n736), .DIN2(n772), .Q(n1436) );
  nnd2s3 U574 ( .DIN1(n1438), .DIN2(n1439), .Q(g8668) );
  nnd2s3 U575 ( .DIN1(n1427), .DIN2(g951), .Q(n1439) );
  nnd2s3 U576 ( .DIN1(n736), .DIN2(n2304), .Q(n1438) );
  nnd2s3 U577 ( .DIN1(n1442), .DIN2(n1443), .Q(g8667) );
  nnd2s3 U578 ( .DIN1(n1427), .DIN2(g950), .Q(n1443) );
  nnd2s3 U579 ( .DIN1(n736), .DIN2(n854), .Q(n1442) );
  nnd2s3 U580 ( .DIN1(n1447), .DIN2(n1448), .Q(g8666) );
  nnd2s3 U581 ( .DIN1(n1427), .DIN2(g949), .Q(n1448) );
  nnd2s3 U582 ( .DIN1(n736), .DIN2(n793), .Q(n1447) );
  nnd2s3 U583 ( .DIN1(n1450), .DIN2(n1466), .Q(g8665) );
  nnd2s3 U584 ( .DIN1(n1427), .DIN2(g948), .Q(n1466) );
  nnd2s3 U585 ( .DIN1(n736), .DIN2(n687), .Q(n1450) );
  nnd2s3 U586 ( .DIN1(n736), .DIN2(n1511), .Q(g8664) );
  nor2s3 U587 ( .DIN1(n1308), .DIN2(n1467), .Q(g8227) );
  xnr2s3 U588 ( .DIN1(n1451), .DIN2(n1371), .Q(n1467) );
  nnd2s3 U589 ( .DIN1(n1476), .DIN2(n1478), .Q(g8226) );
  nnd2s3 U590 ( .DIN1(n1479), .DIN2(n796), .Q(n1478) );
  xor2s3 U591 ( .DIN1(g7732), .DIN2(n1483), .Q(n1479) );
  nnd2s3 U592 ( .DIN1(n1481), .DIN2(n2057), .Q(n1476) );
  nnd2s3 U593 ( .DIN1(n1402), .DIN2(n1485), .Q(g8225) );
  xor2s3 U594 ( .DIN1(n729), .DIN2(n1487), .Q(n1485) );
  nnd2s3 U595 ( .DIN1(n690), .DIN2(n685), .Q(n1487) );
  nnd2s3 U596 ( .DIN1(n1491), .DIN2(n1493), .Q(g8224) );
  nnd2s3 U598 ( .DIN1(n1497), .DIN2(n838), .Q(n1491) );
  nor2s3 U599 ( .DIN1(n1498), .DIN2(n1308), .Q(g7775) );
  and2s3 U600 ( .DIN1(n1499), .DIN2(n1500), .Q(n1498) );
  nnd3s3 U601 ( .DIN1(n1501), .DIN2(n824), .DIN3(n1503), .Q(n1500) );
  nnd2s3 U602 ( .DIN1(n1371), .DIN2(n705), .Q(n1499) );
  or2s3 U603 ( .DIN1(n1501), .DIN2(n698), .Q(n1371) );
  or4s3 U604 ( .DIN1(n1505), .DIN2(n2062), .DIN3(n2059), .DIN4(n2055), .Q(
        n1501) );
  nor2s3 U605 ( .DIN1(n1308), .DIN2(n1507), .Q(g7774) );
  xor2s3 U606 ( .DIN1(n824), .DIN2(n650), .Q(n1507) );
  and3s3 U607 ( .DIN1(n1509), .DIN2(n650), .DIN3(n649), .Q(g7773) );
  nor2s3 U608 ( .DIN1(n1510), .DIN2(n2062), .Q(n1503) );
  nnd2s3 U609 ( .DIN1(n2062), .DIN2(n1510), .Q(n1509) );
  nor2s3 U610 ( .DIN1(n1512), .DIN2(n1308), .Q(g7772) );
  and2s3 U611 ( .DIN1(n1514), .DIN2(n1515), .Q(n1512) );
  nnd3s3 U612 ( .DIN1(n1505), .DIN2(n648), .DIN3(n1516), .Q(n1515) );
  nnd2s3 U613 ( .DIN1(n1510), .DIN2(n867), .Q(n1514) );
  nor2s3 U614 ( .DIN1(n1308), .DIN2(n1517), .Q(g7771) );
  xor2s3 U615 ( .DIN1(n2067), .DIN2(n1516), .Q(n1517) );
  nor2s3 U616 ( .DIN1(n1518), .DIN2(n1455), .Q(n1516) );
  nor2s3 U617 ( .DIN1(n1308), .DIN2(n1519), .Q(g7770) );
  xnr2s3 U618 ( .DIN1(n1455), .DIN2(n1518), .Q(n1519) );
  and3s3 U619 ( .DIN1(n1520), .DIN2(n1518), .DIN3(n649), .Q(g7769) );
  nnd2s3 U620 ( .DIN1(n1483), .DIN2(n1521), .Q(n1308) );
  nnd2s3 U621 ( .DIN1(n1481), .DIN2(n1522), .Q(n1521) );
  xor2s3 U622 ( .DIN1(n2056), .DIN2(n2057), .Q(n1522) );
  or5s3 U623 ( .DIN1(n1523), .DIN2(n1510), .DIN3(n1481), .DIN4(n1524), .DIN5(
        n1526), .Q(n1483) );
  or4s3 U624 ( .DIN1(n1451), .DIN2(n2064), .DIN3(n2063), .DIN4(n2058), .Q(
        n1526) );
  nor2s3 U625 ( .DIN1(n2060), .DIN2(n1527), .Q(n1524) );
  nor2s3 U626 ( .DIN1(n2062), .DIN2(n2061), .Q(n1527) );
  nor2s3 U627 ( .DIN1(n797), .DIN2(n2065), .Q(n1481) );
  or2s3 U628 ( .DIN1(n1505), .DIN2(n698), .Q(n1510) );
  or4s3 U629 ( .DIN1(n1455), .DIN2(n2068), .DIN3(n2067), .DIN4(n2066), .Q(
        n1505) );
  nor2s3 U630 ( .DIN1(n840), .DIN2(n705), .Q(n1523) );
  or2s3 U631 ( .DIN1(n698), .DIN2(n2066), .Q(n1518) );
  nnd2s3 U632 ( .DIN1(n2066), .DIN2(n698), .Q(n1520) );
  and3s3 U633 ( .DIN1(n1375), .DIN2(n830), .DIN3(n1528), .Q(g7768) );
  nnd2s3 U634 ( .DIN1(n1430), .DIN2(n1529), .Q(n1528) );
  nnd2s3 U635 ( .DIN1(n1530), .DIN2(n669), .Q(n1529) );
  or3s3 U636 ( .DIN1(n1430), .DIN2(n2164), .DIN3(n689), .Q(n1375) );
  or5s3 U637 ( .DIN1(n2069), .DIN2(g7423), .DIN3(n2299), .DIN4(g7425), .DIN5(
        g7424), .Q(g7767) );
  nor2s3 U638 ( .DIN1(n1378), .DIN2(n2072), .Q(n2299) );
  nnd4s2 U639 ( .DIN1(n685), .DIN2(n759), .DIN3(n1531), .DIN4(n1532), .Q(n1378) );
  and3s3 U640 ( .DIN1(n809), .DIN2(n729), .DIN3(n733), .Q(n1532) );
  nnd2s3 U641 ( .DIN1(n1402), .DIN2(n1533), .Q(g7766) );
  xor2s3 U642 ( .DIN1(n685), .DIN2(n1489), .Q(n1533) );
  nnd2s3 U643 ( .DIN1(n1534), .DIN2(n1535), .Q(g7765) );
  nnd2s3 U645 ( .DIN1(n1497), .DIN2(n814), .Q(n1534) );
  nnd2s3 U646 ( .DIN1(n1313), .DIN2(n1536), .Q(n1497) );
  nnd2s3 U647 ( .DIN1(n1495), .DIN2(n1236), .Q(n1536) );
  nnd2s3 U648 ( .DIN1(n659), .DIN2(n814), .Q(n1495) );
  xnr2s3 U649 ( .DIN1(g786), .DIN2(n1538), .Q(g7763) );
  nnd2s3 U650 ( .DIN1(n1539), .DIN2(n750), .Q(n1538) );
  xor2s3 U651 ( .DIN1(n750), .DIN2(n1539), .Q(g7762) );
  xor2s3 U652 ( .DIN1(n2084), .DIN2(n1416), .Q(g7761) );
  nor2s3 U653 ( .DIN1(n1540), .DIN2(n1541), .Q(g7759) );
  nor2s3 U654 ( .DIN1(n1542), .DIN2(n856), .Q(n1540) );
  nor2s3 U655 ( .DIN1(n2089), .DIN2(n1543), .Q(n1542) );
  nor2s3 U656 ( .DIN1(n1541), .DIN2(n1544), .Q(g7758) );
  xnr2s3 U657 ( .DIN1(n2089), .DIN2(n1543), .Q(n1544) );
  nnd2s3 U658 ( .DIN1(n1545), .DIN2(n1546), .Q(g7757) );
  nnd3s3 U659 ( .DIN1(n731), .DIN2(n813), .DIN3(n1463), .Q(n1546) );
  nnd2s3 U660 ( .DIN1(g7756), .DIN2(n864), .Q(n1545) );
  nor2s3 U661 ( .DIN1(n813), .DIN2(n1541), .Q(g7756) );
  nor2s3 U662 ( .DIN1(n1986), .DIN2(n2278), .Q(g7739) );
  and2s3 U663 ( .DIN1(n1547), .DIN2(n1548), .Q(g7733) );
  nnd3s3 U664 ( .DIN1(n1549), .DIN2(n757), .DIN3(n688), .Q(n1548) );
  nnd2s3 U665 ( .DIN1(n1550), .DIN2(n1551), .Q(n1547) );
  nnd2s3 U666 ( .DIN1(n1549), .DIN2(n757), .Q(n1551) );
  xor2s3 U667 ( .DIN1(n1552), .DIN2(n1553), .Q(n1550) );
  xor2s3 U668 ( .DIN1(n1554), .DIN2(n1555), .Q(n1553) );
  xor2s3 U669 ( .DIN1(n1496), .DIN2(n1429), .Q(n1555) );
  xor2s3 U670 ( .DIN1(n2304), .DIN2(n1511), .Q(n1554) );
  xor2s3 U671 ( .DIN1(n1556), .DIN2(n1557), .Q(n1552) );
  xor2s3 U672 ( .DIN1(n1428), .DIN2(n1414), .Q(n1557) );
  xor2s3 U673 ( .DIN1(n854), .DIN2(n1413), .Q(n1556) );
  nnd2s3 U674 ( .DIN1(\DFF_98/net323 ), .DIN2(\DFF_175/net400 ), .Q(g7731) );
  nor2s3 U675 ( .DIN1(n1403), .DIN2(n1558), .Q(g7530) );
  xor2s3 U676 ( .DIN1(n669), .DIN2(n689), .Q(n1558) );
  and3s3 U677 ( .DIN1(n689), .DIN2(n830), .DIN3(n1559), .Q(g7529) );
  nnd2s3 U678 ( .DIN1(n1424), .DIN2(n1560), .Q(n1559) );
  nor2s3 U679 ( .DIN1(n1560), .DIN2(n1424), .Q(n1530) );
  and3s3 U680 ( .DIN1(n1560), .DIN2(n830), .DIN3(n1561), .Q(g7528) );
  nnd2s3 U681 ( .DIN1(n704), .DIN2(n1562), .Q(n1561) );
  or2s3 U682 ( .DIN1(n704), .DIN2(n1562), .Q(n1560) );
  nnd3s3 U683 ( .DIN1(n1563), .DIN2(n893), .DIN3(n1422), .Q(g7527) );
  or4s3 U684 ( .DIN1(n2264), .DIN2(n2263), .DIN3(n2262), .DIN4(n2261), .Q(n893) );
  xor2s3 U685 ( .DIN1(n2263), .DIN2(n1564), .Q(n1563) );
  nnd2s3 U686 ( .DIN1(n1565), .DIN2(n1566), .Q(g7525) );
  nnd2s3 U688 ( .DIN1(n1567), .DIN2(n714), .Q(n1565) );
  nnd2s3 U689 ( .DIN1(n1568), .DIN2(n1569), .Q(g7524) );
  nnd2s3 U691 ( .DIN1(n1567), .DIN2(n850), .Q(n1568) );
  nnd2s3 U692 ( .DIN1(n1313), .DIN2(n1571), .Q(n1567) );
  nnd2s3 U693 ( .DIN1(n1570), .DIN2(n1236), .Q(n1571) );
  nnd2s3 U694 ( .DIN1(n1572), .DIN2(n1573), .Q(g7523) );
  nnd2s3 U696 ( .DIN1(n1575), .DIN2(n662), .Q(n1572) );
  nnd2s3 U697 ( .DIN1(n1313), .DIN2(n1576), .Q(n1575) );
  nnd2s3 U698 ( .DIN1(n1574), .DIN2(n1236), .Q(n1576) );
  nnd2s3 U699 ( .DIN1(n1577), .DIN2(n1578), .Q(g7522) );
  nnd2s3 U701 ( .DIN1(n1579), .DIN2(n692), .Q(n1577) );
  nnd2s3 U702 ( .DIN1(n1313), .DIN2(n1580), .Q(n1579) );
  nnd2s3 U703 ( .DIN1(n1441), .DIN2(n1236), .Q(n1580) );
  nnd3s3 U704 ( .DIN1(n1581), .DIN2(n1582), .DIN3(n1402), .Q(g7521) );
  nnd3s3 U705 ( .DIN1(n1583), .DIN2(n759), .DIN3(n2075), .Q(n1582) );
  nnd2s3 U706 ( .DIN1(n1489), .DIN2(n733), .Q(n1581) );
  nnd3s3 U707 ( .DIN1(n759), .DIN2(n733), .DIN3(n1583), .Q(n1489) );
  nnd2s3 U708 ( .DIN1(n1584), .DIN2(n1585), .Q(g7520) );
  nnd2s3 U710 ( .DIN1(n678), .DIN2(n874), .Q(n1584) );
  nnd2s3 U711 ( .DIN1(n1586), .DIN2(n1587), .Q(g7519) );
  and3s3 U713 ( .DIN1(n1236), .DIN2(n679), .DIN3(n1419), .Q(n1238) );
  nnd2s3 U714 ( .DIN1(n1588), .DIN2(n858), .Q(n1586) );
  nnd2s3 U715 ( .DIN1(n1313), .DIN2(n1589), .Q(n1588) );
  nnd2s3 U716 ( .DIN1(n1537), .DIN2(n1236), .Q(n1589) );
  nnd3s3 U717 ( .DIN1(n714), .DIN2(n858), .DIN3(n660), .Q(n1537) );
  nnd2s3 U718 ( .DIN1(n661), .DIN2(n850), .Q(n1570) );
  nnd3s3 U719 ( .DIN1(n692), .DIN2(n662), .DIN3(n874), .Q(n1574) );
  nnd2s3 U720 ( .DIN1(n1236), .DIN2(n1590), .Q(n1313) );
  nnd2s3 U721 ( .DIN1(n1419), .DIN2(n679), .Q(n1590) );
  nnd2s3 U722 ( .DIN1(n745), .DIN2(n679), .Q(n1236) );
  and3s3 U723 ( .DIN1(n725), .DIN2(n797), .DIN3(n2079), .Q(g7518) );
  nnd3s3 U724 ( .DIN1(g43), .DIN2(g1033), .DIN3(n1446), .Q(g9132) );
  nor2s3 U725 ( .DIN1(g43), .DIN2(n1591), .Q(g7517) );
  xor2s3 U726 ( .DIN1(n653), .DIN2(n1592), .Q(n1591) );
  and3s3 U727 ( .DIN1(n1592), .DIN2(g6850), .DIN3(n1593), .Q(g7516) );
  nnd2s3 U728 ( .DIN1(n1464), .DIN2(n1393), .Q(n1593) );
  or2s3 U729 ( .DIN1(n1464), .DIN2(n1393), .Q(n1592) );
  and3s3 U730 ( .DIN1(n1347), .DIN2(g6850), .DIN3(n1393), .Q(g7515) );
  nnd3s3 U731 ( .DIN1(n1393), .DIN2(n653), .DIN3(n1464), .Q(n1347) );
  nor2s3 U732 ( .DIN1(n1401), .DIN2(g7104), .Q(g7514) );
  nnd2s3 U733 ( .DIN1(n1594), .DIN2(n1595), .Q(g7513) );
  nnd2s3 U734 ( .DIN1(n787), .DIN2(n1596), .Q(n1595) );
  nnd2s3 U735 ( .DIN1(n826), .DIN2(n1597), .Q(n1596) );
  nnd2s3 U736 ( .DIN1(g786), .DIN2(n750), .Q(n1597) );
  nnd2s3 U737 ( .DIN1(n1598), .DIN2(n826), .Q(n1594) );
  nnd2s3 U738 ( .DIN1(n1599), .DIN2(n1600), .Q(g7512) );
  nnd3s3 U739 ( .DIN1(n1539), .DIN2(n750), .DIN3(g786), .Q(n1600) );
  nor2s3 U740 ( .DIN1(n1598), .DIN2(n2083), .Q(n1539) );
  nnd2s3 U741 ( .DIN1(n1601), .DIN2(n1598), .Q(n1599) );
  or3s3 U742 ( .DIN1(n1472), .DIN2(n2084), .DIN3(n1416), .Q(n1598) );
  nnd2s3 U743 ( .DIN1(n1472), .DIN2(n1602), .Q(n1601) );
  or2s3 U744 ( .DIN1(n1416), .DIN2(n2084), .Q(n1602) );
  nnd2s3 U745 ( .DIN1(n731), .DIN2(n1603), .Q(g7511) );
  nnd2s3 U746 ( .DIN1(n1604), .DIN2(n1543), .Q(n1603) );
  nnd2s3 U747 ( .DIN1(n732), .DIN2(n1605), .Q(n1604) );
  nnd2s3 U748 ( .DIN1(n731), .DIN2(n1606), .Q(g7510) );
  xor2s3 U749 ( .DIN1(n2092), .DIN2(n1607), .Q(n1606) );
  nor2s3 U750 ( .DIN1(n1463), .DIN2(n2093), .Q(n1607) );
  nnd2s3 U751 ( .DIN1(g781), .DIN2(n896), .Q(n1541) );
  or3s3 U752 ( .DIN1(n2090), .DIN2(n2089), .DIN3(n1543), .Q(n896) );
  or2s3 U753 ( .DIN1(n732), .DIN2(n1605), .Q(n1543) );
  or3s3 U754 ( .DIN1(n2093), .DIN2(n2092), .DIN3(n1463), .Q(n1605) );
  nnd3s3 U755 ( .DIN1(n898), .DIN2(n880), .DIN3(n2081), .Q(n919) );
  nnd2s3 U756 ( .DIN1(g6307), .DIN2(n881), .Q(n1549) );
  nor2s3 U757 ( .DIN1(g6306), .DIN2(g6305), .Q(n898) );
  nnd2s3 U758 ( .DIN1(n881), .DIN2(n1608), .Q(g7474) );
  nnd2s3 U759 ( .DIN1(n1388), .DIN2(n737), .Q(n1608) );
  nnd2s3 U760 ( .DIN1(n1609), .DIN2(n1610), .Q(g7309) );
  xor2s3 U762 ( .DIN1(n693), .DIN2(n1612), .Q(n1611) );
  nnd2s3 U763 ( .DIN1(n719), .DIN2(g93), .Q(n1609) );
  nor2s3 U764 ( .DIN1(n1613), .DIN2(n719), .Q(g7308) );
  nor2s3 U765 ( .DIN1(n1614), .DIN2(g7504), .Q(n1613) );
  nor2s3 U766 ( .DIN1(n693), .DIN2(n1612), .Q(n1614) );
  nnd2s3 U767 ( .DIN1(n1615), .DIN2(n1616), .Q(g7307) );
  nnd3s3 U769 ( .DIN1(n802), .DIN2(n808), .DIN3(n1618), .Q(n1612) );
  nnd2s3 U770 ( .DIN1(n1473), .DIN2(n1619), .Q(n1617) );
  nnd2s3 U771 ( .DIN1(n1618), .DIN2(n808), .Q(n1619) );
  nnd2s3 U772 ( .DIN1(n719), .DIN2(g98), .Q(n1615) );
  nnd2s3 U773 ( .DIN1(n1620), .DIN2(n1621), .Q(g7306) );
  xor2s3 U775 ( .DIN1(n808), .DIN2(n1618), .Q(n1622) );
  nor2s3 U776 ( .DIN1(n1623), .DIN2(n2087), .Q(n1618) );
  nnd2s3 U777 ( .DIN1(n719), .DIN2(g103), .Q(n1620) );
  nnd2s3 U778 ( .DIN1(n1624), .DIN2(n1625), .Q(g7305) );
  xor2s3 U780 ( .DIN1(n1623), .DIN2(n2087), .Q(n1626) );
  nnd2s3 U781 ( .DIN1(n719), .DIN2(g108), .Q(n1624) );
  nor2s3 U782 ( .DIN1(n869), .DIN2(n1627), .Q(g7304) );
  xnr2s3 U783 ( .DIN1(n2262), .DIN2(n1628), .Q(n1627) );
  and3s3 U784 ( .DIN1(n1629), .DIN2(n1628), .DIN3(n1422), .Q(g7303) );
  or2s3 U785 ( .DIN1(n1630), .DIN2(n2261), .Q(n1628) );
  nnd2s3 U786 ( .DIN1(n2261), .DIN2(n1630), .Q(n1629) );
  and2s3 U787 ( .DIN1(n1422), .DIN2(n1631), .Q(g7302) );
  nnd2s3 U788 ( .DIN1(n1632), .DIN2(n1633), .Q(n1631) );
  nnd3s3 U789 ( .DIN1(n1564), .DIN2(n861), .DIN3(n2264), .Q(n1633) );
  nnd2s3 U790 ( .DIN1(n1630), .DIN2(n777), .Q(n1632) );
  nnd3s3 U791 ( .DIN1(n777), .DIN2(n861), .DIN3(n1564), .Q(n1630) );
  nor2s3 U792 ( .DIN1(n894), .DIN2(n2171), .Q(n1564) );
  or4s3 U793 ( .DIN1(n1449), .DIN2(n2267), .DIN3(n2266), .DIN4(n2265), .Q(n894) );
  nor2s3 U794 ( .DIN1(n869), .DIN2(n1634), .Q(g7301) );
  xor2s3 U795 ( .DIN1(n2267), .DIN2(n1635), .Q(n1634) );
  nor2s3 U796 ( .DIN1(n2265), .DIN2(n1636), .Q(n1635) );
  nnd2s3 U798 ( .DIN1(n1638), .DIN2(n756), .Q(n1637) );
  xor2s3 U799 ( .DIN1(n1639), .DIN2(n1480), .Q(n1638) );
  nnd2s3 U800 ( .DIN1(n1402), .DIN2(n1640), .Q(g7299) );
  xor2s3 U801 ( .DIN1(n2088), .DIN2(n1583), .Q(n1640) );
  nor2s3 U802 ( .DIN1(n875), .DIN2(n667), .Q(g7298) );
  and3s3 U803 ( .DIN1(n1562), .DIN2(n830), .DIN3(n1641), .Q(g7119) );
  nnd2s3 U804 ( .DIN1(n1410), .DIN2(n1642), .Q(n1641) );
  or2s3 U805 ( .DIN1(n1643), .DIN2(n1408), .Q(n1642) );
  or3s3 U806 ( .DIN1(n1408), .DIN2(n1410), .DIN3(n1643), .Q(n1562) );
  nnd2s3 U807 ( .DIN1(n1644), .DIN2(n1645), .Q(g7118) );
  nnd3s3 U809 ( .DIN1(n2095), .DIN2(n1647), .DIN3(n2094), .Q(n1623) );
  nnd2s3 U810 ( .DIN1(n744), .DIN2(n1648), .Q(n1646) );
  nnd2s3 U811 ( .DIN1(n2095), .DIN2(n1647), .Q(n1648) );
  nnd2s3 U812 ( .DIN1(n719), .DIN2(g113), .Q(n1644) );
  nnd2s3 U813 ( .DIN1(n1649), .DIN2(n1650), .Q(g7117) );
  xor2s3 U815 ( .DIN1(n2095), .DIN2(n1647), .Q(n1651) );
  nor2s3 U816 ( .DIN1(n1652), .DIN2(n2096), .Q(n1647) );
  nnd2s3 U817 ( .DIN1(n719), .DIN2(g117), .Q(n1649) );
  nnd2s3 U818 ( .DIN1(n1653), .DIN2(n1654), .Q(g7116) );
  xor2s3 U820 ( .DIN1(n1652), .DIN2(n2096), .Q(n1655) );
  nnd2s3 U821 ( .DIN1(n719), .DIN2(g121), .Q(n1653) );
  nnd2s3 U822 ( .DIN1(n1656), .DIN2(n1657), .Q(g7115) );
  nnd3s3 U824 ( .DIN1(n1659), .DIN2(n768), .DIN3(n2097), .Q(n1652) );
  nnd2s3 U825 ( .DIN1(n682), .DIN2(n1660), .Q(n1658) );
  nnd2s3 U826 ( .DIN1(n1659), .DIN2(n768), .Q(n1660) );
  nnd2s3 U827 ( .DIN1(n719), .DIN2(g125), .Q(n1656) );
  nnd2s3 U828 ( .DIN1(n1661), .DIN2(n1662), .Q(g7114) );
  xor2s3 U830 ( .DIN1(n768), .DIN2(n1659), .Q(n1663) );
  nor2s3 U831 ( .DIN1(n1664), .DIN2(n2099), .Q(n1659) );
  nnd2s3 U832 ( .DIN1(n719), .DIN2(g129), .Q(n1661) );
  nnd2s3 U833 ( .DIN1(n1665), .DIN2(n1666), .Q(g7113) );
  xor2s3 U835 ( .DIN1(n1664), .DIN2(n2099), .Q(n1667) );
  nnd2s3 U836 ( .DIN1(n719), .DIN2(g133), .Q(n1665) );
  nor2s3 U837 ( .DIN1(n869), .DIN2(n1668), .Q(g7112) );
  xnr2s3 U838 ( .DIN1(n2265), .DIN2(n1636), .Q(n1668) );
  nnd2s3 U839 ( .DIN1(n1669), .DIN2(n773), .Q(n1636) );
  nnd2s3 U840 ( .DIN1(g1253), .DIN2(n895), .Q(g7111) );
  nnd2s3 U841 ( .DIN1(n1670), .DIN2(n830), .Q(n895) );
  nnd2s3 U842 ( .DIN1(n1671), .DIN2(n1672), .Q(n1670) );
  nnd2s3 U843 ( .DIN1(n2172), .DIN2(n2173), .Q(n1672) );
  nnd3s3 U845 ( .DIN1(n755), .DIN2(n728), .DIN3(n1674), .Q(n1639) );
  nnd2s3 U846 ( .DIN1(n1675), .DIN2(n1488), .Q(n1673) );
  nnd2s3 U847 ( .DIN1(n1674), .DIN2(n728), .Q(n1675) );
  xor2s3 U849 ( .DIN1(n728), .DIN2(n702), .Q(n1676) );
  nnd2s3 U851 ( .DIN1(n1678), .DIN2(n702), .Q(n1677) );
  nor2s3 U852 ( .DIN1(n1679), .DIN2(n1490), .Q(n1674) );
  nnd2s3 U853 ( .DIN1(n1679), .DIN2(n1490), .Q(n1678) );
  nnd3s3 U854 ( .DIN1(n1680), .DIN2(n1681), .DIN3(n1402), .Q(g7107) );
  or3s3 U855 ( .DIN1(n1531), .DIN2(n2132), .DIN3(n1682), .Q(n1681) );
  or2s3 U856 ( .DIN1(n1583), .DIN2(n2100), .Q(n1680) );
  nor2s3 U857 ( .DIN1(n707), .DIN2(n2134), .Q(n1583) );
  nor4s3 U858 ( .DIN1(n1454), .DIN2(n2133), .DIN3(n2132), .DIN4(n2100), .Q(
        n1531) );
  xor2s3 U859 ( .DIN1(n776), .DIN2(n1683), .Q(g7106) );
  nnd2s3 U860 ( .DIN1(n1684), .DIN2(n1685), .Q(n1683) );
  or3s3 U861 ( .DIN1(n1456), .DIN2(n2175), .DIN3(n1407), .Q(n1685) );
  nnd2s3 U862 ( .DIN1(n2101), .DIN2(g43), .Q(n1369) );
  nor2s3 U863 ( .DIN1(n667), .DIN2(g6289), .Q(g7103) );
  nnd2s3 U864 ( .DIN1(n1686), .DIN2(n1687), .Q(g7102) );
  nnd2s3 U865 ( .DIN1(n1469), .DIN2(g6290), .Q(n1687) );
  nnd2s3 U866 ( .DIN1(n801), .DIN2(g12), .Q(n1686) );
  nnd3s3 U867 ( .DIN1(n1688), .DIN2(n1689), .DIN3(n1690), .Q(g7101) );
  or4s3 U868 ( .DIN1(n742), .DIN2(n1417), .DIN3(n1432), .DIN4(n1457), .Q(n1689) );
  nnd2s3 U869 ( .DIN1(n1468), .DIN2(n1691), .Q(n1688) );
  nnd2s3 U870 ( .DIN1(n1692), .DIN2(n1693), .Q(n1691) );
  nnd4s2 U871 ( .DIN1(n2102), .DIN2(n765), .DIN3(n1465), .DIN4(n742), .Q(n1693) );
  nnd2s3 U872 ( .DIN1(n1694), .DIN2(n1695), .Q(n1692) );
  nnd2s3 U873 ( .DIN1(n1417), .DIN2(n1696), .Q(n1695) );
  nnd2s3 U874 ( .DIN1(n1697), .DIN2(n1698), .Q(n1696) );
  nnd2s3 U875 ( .DIN1(n1465), .DIN2(n1699), .Q(n1697) );
  nnd3s3 U876 ( .DIN1(n1700), .DIN2(n1701), .DIN3(n1690), .Q(g7100) );
  nnd2s3 U877 ( .DIN1(g5164), .DIN2(n1698), .Q(n1690) );
  nnd3s3 U878 ( .DIN1(n849), .DIN2(n671), .DIN3(n1694), .Q(n1701) );
  nnd2s3 U879 ( .DIN1(n765), .DIN2(n1702), .Q(n1700) );
  nnd2s3 U880 ( .DIN1(n1703), .DIN2(n1704), .Q(n1702) );
  nnd2s3 U881 ( .DIN1(n2102), .DIN2(n742), .Q(n1704) );
  nnd2s3 U882 ( .DIN1(n2281), .DIN2(n1405), .Q(n1703) );
  nnd3s3 U883 ( .DIN1(n1705), .DIN2(n1706), .DIN3(n1707), .Q(g7099) );
  nnd2s3 U884 ( .DIN1(n1698), .DIN2(n766), .Q(n1707) );
  nnd2s3 U885 ( .DIN1(n1405), .DIN2(n1708), .Q(n1705) );
  nnd3s3 U886 ( .DIN1(n1709), .DIN2(n1710), .DIN3(n1432), .Q(n1708) );
  nnd4s2 U887 ( .DIN1(n1417), .DIN2(n1699), .DIN3(n1698), .DIN4(n671), .Q(
        n1710) );
  or5s3 U888 ( .DIN1(n863), .DIN2(n758), .DIN3(n747), .DIN4(n870), .DIN5(n1711), .Q(n1699) );
  nnd4s2 U889 ( .DIN1(n1383), .DIN2(n1382), .DIN3(n1380), .DIN4(n1379), .Q(
        n1711) );
  nnd2s3 U890 ( .DIN1(n1712), .DIN2(n763), .Q(n1709) );
  nnd2s3 U891 ( .DIN1(n717), .DIN2(n1417), .Q(n1712) );
  nnd2s3 U892 ( .DIN1(n1471), .DIN2(g944), .Q(g7048) );
  xor2s3 U893 ( .DIN1(n2103), .DIN2(n1506), .Q(g6891) );
  xor2s3 U894 ( .DIN1(n2104), .DIN2(n1490), .Q(g6890) );
  xor2s3 U895 ( .DIN1(n2105), .DIN2(n1477), .Q(g6889) );
  xor2s3 U896 ( .DIN1(n2106), .DIN2(n1482), .Q(g6888) );
  xor2s3 U897 ( .DIN1(n2107), .DIN2(n1508), .Q(g6887) );
  xor2s3 U898 ( .DIN1(n2108), .DIN2(n1492), .Q(g6886) );
  xor2s3 U899 ( .DIN1(n2109), .DIN2(n1502), .Q(g6885) );
  xor2s3 U900 ( .DIN1(n2110), .DIN2(n1486), .Q(g6884) );
  xor2s3 U901 ( .DIN1(n2111), .DIN2(n1484), .Q(g6883) );
  xor2s3 U902 ( .DIN1(n2112), .DIN2(n1513), .Q(g6882) );
  xor2s3 U903 ( .DIN1(n2113), .DIN2(n1494), .Q(g6881) );
  xor2s3 U904 ( .DIN1(n2114), .DIN2(n1488), .Q(g6880) );
  xor2s3 U905 ( .DIN1(n2115), .DIN2(n1480), .Q(g6879) );
  xor2s3 U906 ( .DIN1(n2116), .DIN2(n1506), .Q(g6878) );
  xor2s3 U907 ( .DIN1(n2117), .DIN2(n1490), .Q(g6877) );
  xor2s3 U908 ( .DIN1(n2118), .DIN2(n1477), .Q(g6876) );
  xor2s3 U909 ( .DIN1(n2120), .DIN2(n1482), .Q(g6875) );
  xor2s3 U910 ( .DIN1(n2121), .DIN2(n1508), .Q(g6874) );
  xor2s3 U911 ( .DIN1(n2122), .DIN2(n1492), .Q(g6873) );
  xor2s3 U912 ( .DIN1(n2123), .DIN2(n1502), .Q(g6872) );
  xor2s3 U913 ( .DIN1(n2124), .DIN2(n1486), .Q(g6871) );
  xor2s3 U914 ( .DIN1(n2125), .DIN2(n1484), .Q(g6870) );
  xor2s3 U915 ( .DIN1(n2126), .DIN2(n1513), .Q(g6869) );
  xor2s3 U916 ( .DIN1(n2127), .DIN2(n1494), .Q(g6868) );
  xor2s3 U917 ( .DIN1(n2128), .DIN2(n1488), .Q(g6867) );
  xor2s3 U918 ( .DIN1(n2129), .DIN2(n1480), .Q(g6866) );
  nor2s3 U919 ( .DIN1(n1403), .DIN2(n1713), .Q(g6865) );
  xnr2s3 U920 ( .DIN1(n1408), .DIN2(n1643), .Q(n1713) );
  and3s3 U921 ( .DIN1(n1643), .DIN2(n830), .DIN3(n1714), .Q(g6864) );
  nnd2s3 U922 ( .DIN1(n1420), .DIN2(n1715), .Q(n1714) );
  nnd2s3 U923 ( .DIN1(n825), .DIN2(n691), .Q(n1715) );
  or3s3 U924 ( .DIN1(n1411), .DIN2(n1420), .DIN3(n1390), .Q(n1643) );
  nnd2s3 U925 ( .DIN1(n1716), .DIN2(n1717), .Q(g6863) );
  nnd3s3 U926 ( .DIN1(n830), .DIN2(n691), .DIN3(n1390), .Q(n1717) );
  nnd2s3 U927 ( .DIN1(g6862), .DIN2(n825), .Q(n1716) );
  nor2s3 U928 ( .DIN1(n691), .DIN2(n1403), .Q(g6862) );
  nnd2s3 U929 ( .DIN1(n1718), .DIN2(n1719), .Q(g6861) );
  or3s3 U931 ( .DIN1(n2260), .DIN2(n2259), .DIN3(n1474), .Q(n1664) );
  nnd2s3 U932 ( .DIN1(n1474), .DIN2(n1721), .Q(n1720) );
  or2s3 U933 ( .DIN1(n2260), .DIN2(n2259), .Q(n1721) );
  nnd2s3 U934 ( .DIN1(n719), .DIN2(g137), .Q(n1718) );
  nnd2s3 U936 ( .DIN1(n1723), .DIN2(n1679), .Q(n1722) );
  or5s3 U937 ( .DIN1(n1513), .DIN2(n1494), .DIN3(n1477), .DIN4(n1724), .DIN5(
        n1725), .Q(n1679) );
  nnd2s3 U938 ( .DIN1(n1726), .DIN2(n1477), .Q(n1723) );
  nnd4s2 U939 ( .DIN1(n760), .DIN2(n701), .DIN3(n709), .DIN4(n739), .Q(n1726)
         );
  xor2s3 U941 ( .DIN1(n746), .DIN2(n1728), .Q(n1727) );
  or2s3 U942 ( .DIN1(n1729), .DIN2(n1508), .Q(n1728) );
  xor2s3 U944 ( .DIN1(n769), .DIN2(n1729), .Q(n1730) );
  nnd2s3 U945 ( .DIN1(n1684), .DIN2(n1731), .Q(g6856) );
  or3s3 U946 ( .DIN1(n2175), .DIN2(n2135), .DIN3(n1407), .Q(n1731) );
  nnd2s3 U947 ( .DIN1(n776), .DIN2(n872), .Q(n1684) );
  nor2s3 U948 ( .DIN1(n722), .DIN2(n1732), .Q(g6855) );
  xnr2s3 U949 ( .DIN1(n2132), .DIN2(n1682), .Q(n1732) );
  nnd2s3 U950 ( .DIN1(n1733), .DIN2(n845), .Q(n1682) );
  nor2s3 U951 ( .DIN1(n722), .DIN2(n1734), .Q(g6854) );
  xor2s3 U952 ( .DIN1(n1454), .DIN2(n1733), .Q(n1734) );
  nor2s3 U953 ( .DIN1(n2133), .DIN2(n2134), .Q(n1733) );
  nor2s3 U954 ( .DIN1(n1735), .DIN2(n722), .Q(g6853) );
  xnr2s3 U955 ( .DIN1(n2133), .DIN2(n2134), .Q(n1735) );
  nnd2s3 U956 ( .DIN1(n1736), .DIN2(n1737), .Q(g6852) );
  nnd2s3 U957 ( .DIN1(n1445), .DIN2(g1080), .Q(n1737) );
  nnd2s3 U958 ( .DIN1(n2135), .DIN2(n723), .Q(n1736) );
  and4s2 U959 ( .DIN1(n1694), .DIN2(n1417), .DIN3(n2248), .DIN4(n1738), .Q(
        g6849) );
  or5s3 U960 ( .DIN1(n1739), .DIN2(n1740), .DIN3(n1741), .DIN4(n1742), .DIN5(
        n1743), .Q(n1738) );
  nnd4s2 U961 ( .DIN1(n1744), .DIN2(n1745), .DIN3(n1746), .DIN4(n1747), .Q(
        n1743) );
  xnr2s3 U962 ( .DIN1(n1380), .DIN2(n2256), .Q(n1747) );
  xnr2s3 U963 ( .DIN1(n1383), .DIN2(n2255), .Q(n1746) );
  xor2s3 U964 ( .DIN1(n870), .DIN2(n2254), .Q(n1745) );
  xor2s3 U965 ( .DIN1(n758), .DIN2(n2253), .Q(n1744) );
  xor2s3 U966 ( .DIN1(n2251), .DIN2(n1382), .Q(n1742) );
  xor2s3 U967 ( .DIN1(n2252), .DIN2(n1379), .Q(n1741) );
  xor2s3 U968 ( .DIN1(n2249), .DIN2(n1421), .Q(n1740) );
  xor2s3 U969 ( .DIN1(n2250), .DIN2(n1394), .Q(n1739) );
  nor2s3 U970 ( .DIN1(n766), .DIN2(n742), .Q(n1694) );
  or5s3 U971 ( .DIN1(n1748), .DIN2(n1749), .DIN3(n1750), .DIN4(n1751), .DIN5(
        n1752), .Q(g6392) );
  nnd4s2 U972 ( .DIN1(n1753), .DIN2(n1754), .DIN3(n1755), .DIN4(n1756), .Q(
        n1752) );
  xnr2s3 U973 ( .DIN1(n2262), .DIN2(n2146), .Q(n1756) );
  xnr2s3 U974 ( .DIN1(n2145), .DIN2(n2266), .Q(n1755) );
  xor2s3 U975 ( .DIN1(n2144), .DIN2(n773), .Q(n1754) );
  xnr2s3 U976 ( .DIN1(n2143), .DIN2(n2265), .Q(n1753) );
  xor2s3 U977 ( .DIN1(n2141), .DIN2(n2263), .Q(n1751) );
  xor2s3 U978 ( .DIN1(n2142), .DIN2(n2267), .Q(n1750) );
  xor2s3 U979 ( .DIN1(n2139), .DIN2(n2261), .Q(n1749) );
  xor2s3 U980 ( .DIN1(n2140), .DIN2(n2264), .Q(n1748) );
  or5s3 U981 ( .DIN1(n691), .DIN2(n1757), .DIN3(n1758), .DIN4(n1759), .DIN5(
        n1760), .Q(g6391) );
  or5s3 U982 ( .DIN1(n1761), .DIN2(n1762), .DIN3(n1763), .DIN4(n1764), .DIN5(
        n1765), .Q(n1760) );
  xor2s3 U983 ( .DIN1(n2154), .DIN2(n2167), .Q(n1765) );
  xor2s3 U984 ( .DIN1(n2155), .DIN2(n2169), .Q(n1764) );
  xor2s3 U985 ( .DIN1(n2149), .DIN2(n1408), .Q(n1763) );
  xor2s3 U986 ( .DIN1(n2147), .DIN2(n1410), .Q(n1762) );
  xor2s3 U987 ( .DIN1(n2152), .DIN2(n1430), .Q(n1761) );
  nnd3s3 U988 ( .DIN1(n1766), .DIN2(n1767), .DIN3(n1390), .Q(n1759) );
  xor2s3 U989 ( .DIN1(n2151), .DIN2(n2164), .Q(n1767) );
  xor2s3 U990 ( .DIN1(n2148), .DIN2(n2161), .Q(n1766) );
  xor2s3 U991 ( .DIN1(n2150), .DIN2(n1420), .Q(n1758) );
  xor2s3 U992 ( .DIN1(n2153), .DIN2(n1424), .Q(n1757) );
  or5s3 U993 ( .DIN1(n1768), .DIN2(n1769), .DIN3(n1770), .DIN4(n1771), .DIN5(
        n1772), .Q(g6386) );
  or5s3 U994 ( .DIN1(n1773), .DIN2(n1774), .DIN3(n1775), .DIN4(n1776), .DIN5(
        n1777), .Q(n1772) );
  xor2s3 U995 ( .DIN1(n2163), .DIN2(n2164), .Q(n1777) );
  xor2s3 U996 ( .DIN1(n2165), .DIN2(n1430), .Q(n1776) );
  xor2s3 U997 ( .DIN1(n2167), .DIN2(n2168), .Q(n1775) );
  xor2s3 U998 ( .DIN1(n2169), .DIN2(n2170), .Q(n1774) );
  xor2s3 U999 ( .DIN1(n2166), .DIN2(n1424), .Q(n1773) );
  nnd3s3 U1000 ( .DIN1(n1778), .DIN2(n1779), .DIN3(n1780), .Q(n1771) );
  xnr2s3 U1001 ( .DIN1(n2162), .DIN2(n1408), .Q(n1780) );
  xor2s3 U1002 ( .DIN1(n2160), .DIN2(n2161), .Q(n1779) );
  xnr2s3 U1003 ( .DIN1(n2159), .DIN2(n1410), .Q(n1778) );
  xor2s3 U1004 ( .DIN1(n2157), .DIN2(n1420), .Q(n1770) );
  xor2s3 U1005 ( .DIN1(n2158), .DIN2(n1411), .Q(n1769) );
  xor2s3 U1006 ( .DIN1(n2156), .DIN2(n1390), .Q(n1768) );
  nnd2s3 U1007 ( .DIN1(\DFF_373/net598 ), .DIN2(n668), .Q(g6385) );
  nor2s3 U1008 ( .DIN1(n797), .DIN2(n2278), .Q(n2297) );
  nor2s3 U1009 ( .DIN1(n869), .DIN2(n1781), .Q(g6384) );
  xor2s3 U1010 ( .DIN1(n1449), .DIN2(n1669), .Q(n1781) );
  nor2s3 U1011 ( .DIN1(n2171), .DIN2(n2266), .Q(n1669) );
  nor2s3 U1012 ( .DIN1(n1782), .DIN2(n869), .Q(g6383) );
  xnr2s3 U1013 ( .DIN1(n2171), .DIN2(n2266), .Q(n1782) );
  nnd2s3 U1014 ( .DIN1(n1671), .DIN2(g1266), .Q(g6382) );
  nnd2s3 U1015 ( .DIN1(n1671), .DIN2(n816), .Q(g6381) );
  nnd2s3 U1016 ( .DIN1(n1671), .DIN2(n818), .Q(g6380) );
  and4s2 U1017 ( .DIN1(n1488), .DIN2(n839), .DIN3(n701), .DIN4(n1783), .Q(
        n1671) );
  and3s3 U1018 ( .DIN1(n834), .DIN2(n728), .DIN3(n726), .Q(n1783) );
  nnd3s3 U1019 ( .DIN1(n703), .DIN2(n769), .DIN3(n746), .Q(n1724) );
  nnd2s3 U1021 ( .DIN1(n1785), .DIN2(n1729), .Q(n1784) );
  nnd3s3 U1022 ( .DIN1(n703), .DIN2(n805), .DIN3(n1786), .Q(n1729) );
  nnd2s3 U1023 ( .DIN1(n1787), .DIN2(n1492), .Q(n1785) );
  nnd2s3 U1024 ( .DIN1(n1786), .DIN2(n805), .Q(n1787) );
  xor2s3 U1026 ( .DIN1(n805), .DIN2(n708), .Q(n1788) );
  nnd2s3 U1028 ( .DIN1(n1790), .DIN2(n708), .Q(n1789) );
  nor2s3 U1029 ( .DIN1(n1791), .DIN2(n1486), .Q(n1786) );
  nnd2s3 U1030 ( .DIN1(n1791), .DIN2(n1486), .Q(n1790) );
  nnd2s3 U1031 ( .DIN1(n1427), .DIN2(n1792), .Q(g6372) );
  nnd2s3 U1032 ( .DIN1(g4655), .DIN2(\DFF_605/net830 ), .Q(n1792) );
  or5s3 U1033 ( .DIN1(n1793), .DIN2(n1794), .DIN3(n1795), .DIN4(n1796), .DIN5(
        n1797), .Q(g6371) );
  nnd4s2 U1034 ( .DIN1(n1798), .DIN2(n1799), .DIN3(n1800), .DIN4(n1801), .Q(
        n1797) );
  and3s3 U1035 ( .DIN1(n1802), .DIN2(n1803), .DIN3(n1804), .Q(n1801) );
  or2s3 U1036 ( .DIN1(n887), .DIN2(n2183), .Q(n1804) );
  or2s3 U1037 ( .DIN1(n885), .DIN2(n2187), .Q(n1803) );
  or2s3 U1038 ( .DIN1(n886), .DIN2(n2185), .Q(n1802) );
  nnd2s3 U1039 ( .DIN1(n810), .DIN2(n684), .Q(n1800) );
  or2s3 U1040 ( .DIN1(n888), .DIN2(n2184), .Q(n1799) );
  or2s3 U1041 ( .DIN1(n889), .DIN2(n2182), .Q(n1798) );
  nnd4s2 U1042 ( .DIN1(n1805), .DIN2(n1806), .DIN3(n1807), .DIN4(n1808), .Q(
        n1796) );
  nnd2s3 U1043 ( .DIN1(g633), .DIN2(n804), .Q(n1808) );
  nnd2s3 U1044 ( .DIN1(g634), .DIN2(n790), .Q(n1807) );
  nnd2s3 U1045 ( .DIN1(g635), .DIN2(n829), .Q(n1806) );
  nnd2s3 U1046 ( .DIN1(g645), .DIN2(n675), .Q(n1805) );
  nor2s3 U1047 ( .DIN1(n2186), .DIN2(n884), .Q(n1795) );
  nor2s3 U1048 ( .DIN1(n2177), .DIN2(n883), .Q(n1794) );
  nor2s3 U1049 ( .DIN1(n2176), .DIN2(n882), .Q(n1793) );
  nnd2s3 U1050 ( .DIN1(n1809), .DIN2(n1810), .Q(g6370) );
  nnd2s3 U1051 ( .DIN1(n696), .DIN2(g587), .Q(n1810) );
  nnd2s3 U1052 ( .DIN1(n1811), .DIN2(n770), .Q(n1809) );
  nnd2s3 U1053 ( .DIN1(n1812), .DIN2(n1813), .Q(g6369) );
  nnd2s3 U1054 ( .DIN1(n696), .DIN2(g583), .Q(n1813) );
  nnd2s3 U1055 ( .DIN1(n1811), .DIN2(n681), .Q(n1812) );
  nnd2s3 U1056 ( .DIN1(n1814), .DIN2(n1815), .Q(g6368) );
  nnd2s3 U1057 ( .DIN1(n696), .DIN2(g579), .Q(n1815) );
  nnd2s3 U1058 ( .DIN1(n1811), .DIN2(n817), .Q(n1814) );
  nnd2s3 U1059 ( .DIN1(n1816), .DIN2(n1817), .Q(g6367) );
  nnd2s3 U1060 ( .DIN1(n696), .DIN2(g566), .Q(n1817) );
  nnd2s3 U1061 ( .DIN1(n1811), .DIN2(n812), .Q(n1816) );
  nnd2s3 U1062 ( .DIN1(n1818), .DIN2(n1819), .Q(g6366) );
  nnd2s3 U1063 ( .DIN1(n696), .DIN2(g556), .Q(n1819) );
  nnd2s3 U1064 ( .DIN1(n1811), .DIN2(n806), .Q(n1818) );
  nnd2s3 U1065 ( .DIN1(n1820), .DIN2(n1821), .Q(g6365) );
  nnd2s3 U1066 ( .DIN1(n696), .DIN2(g543), .Q(n1821) );
  nnd2s3 U1067 ( .DIN1(n1811), .DIN2(n789), .Q(n1820) );
  nnd2s3 U1068 ( .DIN1(n1822), .DIN2(n1823), .Q(g6364) );
  nnd2s3 U1069 ( .DIN1(n696), .DIN2(g539), .Q(n1823) );
  nnd2s3 U1070 ( .DIN1(n1811), .DIN2(n697), .Q(n1822) );
  nnd2s3 U1071 ( .DIN1(n1824), .DIN2(n1825), .Q(g6363) );
  nnd2s3 U1072 ( .DIN1(n696), .DIN2(g535), .Q(n1825) );
  nnd2s3 U1073 ( .DIN1(n1811), .DIN2(n779), .Q(n1824) );
  nnd2s3 U1074 ( .DIN1(g595), .DIN2(\DFF_550/net775 ), .Q(n1811) );
  nnd2s3 U1075 ( .DIN1(n1826), .DIN2(n1827), .Q(g6362) );
  nnd2s3 U1076 ( .DIN1(n794), .DIN2(g517), .Q(n1827) );
  nnd2s3 U1077 ( .DIN1(n1828), .DIN2(n686), .Q(n1826) );
  nnd2s3 U1078 ( .DIN1(n1829), .DIN2(n1830), .Q(g6361) );
  nnd2s3 U1079 ( .DIN1(n794), .DIN2(g516), .Q(n1830) );
  nnd2s3 U1080 ( .DIN1(n1828), .DIN2(n800), .Q(n1829) );
  nnd2s3 U1081 ( .DIN1(n1831), .DIN2(n1832), .Q(g6360) );
  nnd2s3 U1082 ( .DIN1(n794), .DIN2(g479), .Q(n1832) );
  nnd2s3 U1083 ( .DIN1(n1828), .DIN2(n727), .Q(n1831) );
  nnd2s3 U1084 ( .DIN1(n1833), .DIN2(n1834), .Q(g6359) );
  nnd2s3 U1085 ( .DIN1(n794), .DIN2(g478), .Q(n1834) );
  nnd2s3 U1086 ( .DIN1(n1828), .DIN2(n749), .Q(n1833) );
  nnd2s3 U1087 ( .DIN1(n1835), .DIN2(n1836), .Q(g6358) );
  nnd2s3 U1088 ( .DIN1(n794), .DIN2(g477), .Q(n1836) );
  nnd2s3 U1089 ( .DIN1(n1828), .DIN2(n721), .Q(n1835) );
  nnd2s3 U1090 ( .DIN1(n1837), .DIN2(n1838), .Q(g6357) );
  nnd2s3 U1091 ( .DIN1(n794), .DIN2(g476), .Q(n1838) );
  nnd2s3 U1092 ( .DIN1(n1828), .DIN2(n821), .Q(n1837) );
  nnd2s3 U1093 ( .DIN1(n1839), .DIN2(n1840), .Q(g6356) );
  nnd2s3 U1094 ( .DIN1(n794), .DIN2(g475), .Q(n1840) );
  nnd2s3 U1095 ( .DIN1(n1828), .DIN2(n857), .Q(n1839) );
  nnd2s3 U1096 ( .DIN1(n1841), .DIN2(n1842), .Q(g6355) );
  nnd2s3 U1097 ( .DIN1(n794), .DIN2(g474), .Q(n1842) );
  nnd2s3 U1098 ( .DIN1(n1828), .DIN2(n835), .Q(n1841) );
  nnd2s3 U1099 ( .DIN1(n1843), .DIN2(n1844), .Q(g6354) );
  nnd2s3 U1100 ( .DIN1(n794), .DIN2(g458), .Q(n1844) );
  nnd2s3 U1101 ( .DIN1(n1828), .DIN2(n820), .Q(n1843) );
  nnd2s3 U1102 ( .DIN1(n1845), .DIN2(n1846), .Q(g6353) );
  nnd2s3 U1103 ( .DIN1(n794), .DIN2(g457), .Q(n1846) );
  nnd2s3 U1104 ( .DIN1(n1828), .DIN2(n788), .Q(n1845) );
  nnd2s3 U1105 ( .DIN1(n1847), .DIN2(n1848), .Q(g6352) );
  nnd2s3 U1106 ( .DIN1(n794), .DIN2(g456), .Q(n1848) );
  nnd2s3 U1107 ( .DIN1(n1828), .DIN2(n871), .Q(n1847) );
  nnd2s3 U1108 ( .DIN1(n1849), .DIN2(n1850), .Q(g6351) );
  nnd2s3 U1109 ( .DIN1(n794), .DIN2(g455), .Q(n1850) );
  nnd2s3 U1110 ( .DIN1(n1828), .DIN2(n647), .Q(n1849) );
  nnd2s3 U1111 ( .DIN1(n1851), .DIN2(n1852), .Q(g6350) );
  nnd2s3 U1112 ( .DIN1(n794), .DIN2(g454), .Q(n1852) );
  nnd2s3 U1113 ( .DIN1(n1828), .DIN2(n670), .Q(n1851) );
  nnd2s3 U1114 ( .DIN1(g533), .DIN2(\DFF_286/net511 ), .Q(n1828) );
  nnd2s3 U1115 ( .DIN1(n1853), .DIN2(n1854), .Q(g6349) );
  nnd2s3 U1116 ( .DIN1(n832), .DIN2(g436), .Q(n1854) );
  nnd2s3 U1117 ( .DIN1(n1855), .DIN2(n715), .Q(n1853) );
  nnd2s3 U1118 ( .DIN1(n1856), .DIN2(n1857), .Q(g6348) );
  nnd2s3 U1119 ( .DIN1(n832), .DIN2(g435), .Q(n1857) );
  nnd2s3 U1120 ( .DIN1(n1855), .DIN2(n847), .Q(n1856) );
  nnd2s3 U1121 ( .DIN1(n1858), .DIN2(n1859), .Q(g6347) );
  nnd2s3 U1122 ( .DIN1(n832), .DIN2(g398), .Q(n1859) );
  nnd2s3 U1123 ( .DIN1(n1855), .DIN2(n676), .Q(n1858) );
  nnd2s3 U1124 ( .DIN1(n1860), .DIN2(n1861), .Q(g6346) );
  nnd2s3 U1125 ( .DIN1(n832), .DIN2(g397), .Q(n1861) );
  nnd2s3 U1126 ( .DIN1(n1855), .DIN2(n672), .Q(n1860) );
  nnd2s3 U1127 ( .DIN1(n1862), .DIN2(n1863), .Q(g6345) );
  nnd2s3 U1128 ( .DIN1(n832), .DIN2(g396), .Q(n1863) );
  nnd2s3 U1129 ( .DIN1(n1855), .DIN2(n718), .Q(n1862) );
  nnd2s3 U1130 ( .DIN1(n1864), .DIN2(n1865), .Q(g6344) );
  nnd2s3 U1131 ( .DIN1(n832), .DIN2(g395), .Q(n1865) );
  nnd2s3 U1132 ( .DIN1(n1855), .DIN2(n798), .Q(n1864) );
  nnd2s3 U1133 ( .DIN1(n1866), .DIN2(n1867), .Q(g6343) );
  nnd2s3 U1134 ( .DIN1(n832), .DIN2(g394), .Q(n1867) );
  nnd2s3 U1135 ( .DIN1(n1855), .DIN2(n815), .Q(n1866) );
  nnd2s3 U1136 ( .DIN1(n1868), .DIN2(n1869), .Q(g6342) );
  nnd2s3 U1137 ( .DIN1(n832), .DIN2(g393), .Q(n1869) );
  nnd2s3 U1138 ( .DIN1(n1855), .DIN2(n740), .Q(n1868) );
  nnd2s3 U1139 ( .DIN1(n1870), .DIN2(n1871), .Q(g6341) );
  nnd2s3 U1140 ( .DIN1(n832), .DIN2(g377), .Q(n1871) );
  nnd2s3 U1141 ( .DIN1(n1855), .DIN2(n848), .Q(n1870) );
  nnd2s3 U1142 ( .DIN1(n1872), .DIN2(n1873), .Q(g6340) );
  nnd2s3 U1143 ( .DIN1(n832), .DIN2(g376), .Q(n1873) );
  nnd2s3 U1144 ( .DIN1(n1855), .DIN2(n842), .Q(n1872) );
  nnd2s3 U1145 ( .DIN1(n1874), .DIN2(n1875), .Q(g6339) );
  nnd2s3 U1146 ( .DIN1(n832), .DIN2(g375), .Q(n1875) );
  or2s3 U1147 ( .DIN1(n832), .DIN2(n2219), .Q(n1874) );
  nnd2s3 U1148 ( .DIN1(n1876), .DIN2(n1877), .Q(g6338) );
  nnd2s3 U1149 ( .DIN1(n832), .DIN2(g374), .Q(n1877) );
  or2s3 U1150 ( .DIN1(n832), .DIN2(n2220), .Q(n1876) );
  nnd2s3 U1151 ( .DIN1(n1878), .DIN2(n1879), .Q(g6337) );
  nnd2s3 U1152 ( .DIN1(n832), .DIN2(g373), .Q(n1879) );
  or2s3 U1153 ( .DIN1(n832), .DIN2(n2221), .Q(n1878) );
  nnd2s3 U1154 ( .DIN1(g452), .DIN2(\DFF_171/net396 ), .Q(n1855) );
  nnd2s3 U1155 ( .DIN1(n1880), .DIN2(n1881), .Q(g6336) );
  nnd2s3 U1156 ( .DIN1(n762), .DIN2(g355), .Q(n1881) );
  nnd2s3 U1157 ( .DIN1(n1882), .DIN2(n873), .Q(n1880) );
  nnd2s3 U1158 ( .DIN1(n1883), .DIN2(n1884), .Q(g6335) );
  nnd2s3 U1159 ( .DIN1(n762), .DIN2(g354), .Q(n1884) );
  nnd2s3 U1160 ( .DIN1(n1882), .DIN2(n748), .Q(n1883) );
  nnd2s3 U1161 ( .DIN1(n1885), .DIN2(n1886), .Q(g6334) );
  nnd2s3 U1162 ( .DIN1(n762), .DIN2(g317), .Q(n1886) );
  nnd2s3 U1163 ( .DIN1(n1882), .DIN2(n811), .Q(n1885) );
  nnd2s3 U1164 ( .DIN1(n1887), .DIN2(n1888), .Q(g6333) );
  nnd2s3 U1165 ( .DIN1(n762), .DIN2(g316), .Q(n1888) );
  nnd2s3 U1166 ( .DIN1(n1882), .DIN2(n782), .Q(n1887) );
  nnd2s3 U1167 ( .DIN1(n1889), .DIN2(n1890), .Q(g6332) );
  nnd2s3 U1168 ( .DIN1(n762), .DIN2(g315), .Q(n1890) );
  nnd2s3 U1169 ( .DIN1(n1882), .DIN2(n852), .Q(n1889) );
  nnd2s3 U1170 ( .DIN1(n1891), .DIN2(n1892), .Q(g6331) );
  nnd2s3 U1171 ( .DIN1(n762), .DIN2(g314), .Q(n1892) );
  nnd2s3 U1172 ( .DIN1(n1882), .DIN2(n680), .Q(n1891) );
  nnd2s3 U1173 ( .DIN1(n1893), .DIN2(n1894), .Q(g6330) );
  nnd2s3 U1174 ( .DIN1(n762), .DIN2(g313), .Q(n1894) );
  nnd2s3 U1175 ( .DIN1(n1882), .DIN2(n677), .Q(n1893) );
  nnd2s3 U1176 ( .DIN1(n1895), .DIN2(n1896), .Q(g6329) );
  nnd2s3 U1177 ( .DIN1(n762), .DIN2(g312), .Q(n1896) );
  nnd2s3 U1178 ( .DIN1(n1882), .DIN2(n785), .Q(n1895) );
  nnd2s3 U1179 ( .DIN1(n1897), .DIN2(n1898), .Q(g6328) );
  nnd2s3 U1180 ( .DIN1(n762), .DIN2(g296), .Q(n1898) );
  nnd2s3 U1181 ( .DIN1(n1882), .DIN2(n807), .Q(n1897) );
  nnd2s3 U1182 ( .DIN1(n1899), .DIN2(n1900), .Q(g6327) );
  nnd2s3 U1183 ( .DIN1(n762), .DIN2(g295), .Q(n1900) );
  nnd2s3 U1184 ( .DIN1(n1882), .DIN2(n674), .Q(n1899) );
  nnd2s3 U1185 ( .DIN1(n1901), .DIN2(n1902), .Q(g6326) );
  nnd2s3 U1186 ( .DIN1(n762), .DIN2(g294), .Q(n1902) );
  or2s3 U1187 ( .DIN1(n762), .DIN2(n2232), .Q(n1901) );
  nnd2s3 U1188 ( .DIN1(n1903), .DIN2(n1904), .Q(g6325) );
  nnd2s3 U1189 ( .DIN1(n762), .DIN2(g293), .Q(n1904) );
  or2s3 U1190 ( .DIN1(n762), .DIN2(n2233), .Q(n1903) );
  nnd2s3 U1191 ( .DIN1(n1905), .DIN2(n1906), .Q(g6324) );
  nnd2s3 U1192 ( .DIN1(n762), .DIN2(g292), .Q(n1906) );
  or2s3 U1193 ( .DIN1(n762), .DIN2(n2234), .Q(n1905) );
  nnd2s3 U1194 ( .DIN1(g371), .DIN2(\DFF_365/net590 ), .Q(n1882) );
  nnd2s3 U1195 ( .DIN1(n1907), .DIN2(n1908), .Q(g6323) );
  nnd2s3 U1196 ( .DIN1(n771), .DIN2(g274), .Q(n1908) );
  nnd2s3 U1197 ( .DIN1(n1909), .DIN2(n862), .Q(n1907) );
  nnd2s3 U1198 ( .DIN1(n1910), .DIN2(n1911), .Q(g6322) );
  nnd2s3 U1199 ( .DIN1(n771), .DIN2(g273), .Q(n1911) );
  nnd2s3 U1200 ( .DIN1(n1909), .DIN2(n710), .Q(n1910) );
  nnd2s3 U1201 ( .DIN1(n1912), .DIN2(n1913), .Q(g6321) );
  nnd2s3 U1202 ( .DIN1(n771), .DIN2(g236), .Q(n1913) );
  nnd2s3 U1203 ( .DIN1(n1909), .DIN2(n783), .Q(n1912) );
  nnd2s3 U1204 ( .DIN1(n1914), .DIN2(n1915), .Q(g6320) );
  nnd2s3 U1205 ( .DIN1(n771), .DIN2(g235), .Q(n1915) );
  nnd2s3 U1206 ( .DIN1(n1909), .DIN2(n738), .Q(n1914) );
  nnd2s3 U1207 ( .DIN1(n1916), .DIN2(n1917), .Q(g6319) );
  nnd2s3 U1208 ( .DIN1(n771), .DIN2(g234), .Q(n1917) );
  nnd2s3 U1209 ( .DIN1(n1909), .DIN2(n833), .Q(n1916) );
  nnd2s3 U1210 ( .DIN1(n1918), .DIN2(n1919), .Q(g6318) );
  nnd2s3 U1211 ( .DIN1(n771), .DIN2(g233), .Q(n1919) );
  nnd2s3 U1212 ( .DIN1(n1909), .DIN2(n868), .Q(n1918) );
  nnd2s3 U1213 ( .DIN1(n1920), .DIN2(n1921), .Q(g6317) );
  nnd2s3 U1214 ( .DIN1(n771), .DIN2(g232), .Q(n1921) );
  nnd2s3 U1215 ( .DIN1(n1909), .DIN2(n844), .Q(n1920) );
  nnd2s3 U1216 ( .DIN1(n1922), .DIN2(n1923), .Q(g6316) );
  nnd2s3 U1217 ( .DIN1(n771), .DIN2(g231), .Q(n1923) );
  nnd2s3 U1218 ( .DIN1(n1909), .DIN2(n754), .Q(n1922) );
  nnd2s3 U1219 ( .DIN1(n1924), .DIN2(n1925), .Q(g6315) );
  nnd2s3 U1220 ( .DIN1(n771), .DIN2(g215), .Q(n1925) );
  nnd2s3 U1221 ( .DIN1(n1909), .DIN2(n753), .Q(n1924) );
  nnd2s3 U1222 ( .DIN1(n1926), .DIN2(n1927), .Q(g6314) );
  nnd2s3 U1223 ( .DIN1(n771), .DIN2(g214), .Q(n1927) );
  nnd2s3 U1224 ( .DIN1(n1909), .DIN2(n828), .Q(n1926) );
  nnd2s3 U1225 ( .DIN1(n1928), .DIN2(n1929), .Q(g6313) );
  nnd2s3 U1226 ( .DIN1(n771), .DIN2(g213), .Q(n1929) );
  or2s3 U1227 ( .DIN1(n771), .DIN2(n2245), .Q(n1928) );
  nnd2s3 U1228 ( .DIN1(n1930), .DIN2(n1931), .Q(g6312) );
  nnd2s3 U1229 ( .DIN1(n771), .DIN2(g212), .Q(n1931) );
  or2s3 U1230 ( .DIN1(n771), .DIN2(n2246), .Q(n1930) );
  nnd2s3 U1231 ( .DIN1(n1932), .DIN2(n1933), .Q(g6311) );
  nnd2s3 U1232 ( .DIN1(n771), .DIN2(g211), .Q(n1933) );
  or2s3 U1233 ( .DIN1(n771), .DIN2(n2247), .Q(n1932) );
  nnd2s3 U1234 ( .DIN1(g290), .DIN2(\DFF_342/net567 ), .Q(n1909) );
  nnd2s3 U1235 ( .DIN1(n1934), .DIN2(n799), .Q(g5746) );
  xor2s3 U1236 ( .DIN1(n1935), .DIN2(g7508), .Q(n1934) );
  nnd2s3 U1237 ( .DIN1(n2271), .DIN2(n1936), .Q(n1935) );
  nnd2s3 U1238 ( .DIN1(g5180), .DIN2(n1937), .Q(g5745) );
  nnd3s3 U1239 ( .DIN1(n2274), .DIN2(n2275), .DIN3(n2257), .Q(n1937) );
  nnd2s3 U1240 ( .DIN1(g5177), .DIN2(n1938), .Q(g5744) );
  nnd3s3 U1241 ( .DIN1(n2276), .DIN2(n2277), .DIN3(n2258), .Q(n1938) );
  nnd2s3 U1242 ( .DIN1(n1939), .DIN2(n1940), .Q(g5743) );
  xor2s3 U1244 ( .DIN1(n2259), .DIN2(n2260), .Q(n1941) );
  nnd2s3 U1245 ( .DIN1(n719), .DIN2(g141), .Q(n1939) );
  nnd2s3 U1246 ( .DIN1(n1942), .DIN2(n1943), .Q(g5742) );
  nnd2s3 U1247 ( .DIN1(n719), .DIN2(g145), .Q(n1943) );
  nnd4s2 U1249 ( .DIN1(n1486), .DIN2(n1502), .DIN3(n761), .DIN4(n709), .Q(
        g5740) );
  and3s3 U1250 ( .DIN1(n1513), .DIN2(n1494), .DIN3(n760), .Q(g5739) );
  and3s3 U1251 ( .DIN1(n1494), .DIN2(n739), .DIN3(n760), .Q(g5738) );
  and3s3 U1252 ( .DIN1(n1513), .DIN2(n709), .DIN3(n760), .Q(g5737) );
  nnd3s3 U1253 ( .DIN1(n827), .DIN2(n805), .DIN3(n761), .Q(n1725) );
  and3s3 U1254 ( .DIN1(n1791), .DIN2(n756), .DIN3(n1944), .Q(g5736) );
  nnd2s3 U1255 ( .DIN1(n1945), .DIN2(n1946), .Q(n1944) );
  or2s3 U1256 ( .DIN1(g5173), .DIN2(n1494), .Q(n1946) );
  nnd3s3 U1258 ( .DIN1(n709), .DIN2(n739), .DIN3(n761), .Q(n1791) );
  nor2s3 U1259 ( .DIN1(n1947), .DIN2(n735), .Q(g5735) );
  nor2s3 U1260 ( .DIN1(n1948), .DIN2(n651), .Q(g5733) );
  nor2s3 U1261 ( .DIN1(n1949), .DIN2(g5161), .Q(n1948) );
  xor2s3 U1262 ( .DIN1(g210), .DIN2(g1206), .Q(n1949) );
  nor2s3 U1263 ( .DIN1(n1950), .DIN2(n651), .Q(g5732) );
  nor2s3 U1264 ( .DIN1(n1951), .DIN2(g5160), .Q(n1950) );
  xor2s3 U1265 ( .DIN1(g205), .DIN2(g1202), .Q(n1951) );
  nor2s3 U1266 ( .DIN1(n1952), .DIN2(n651), .Q(g5731) );
  nor2s3 U1267 ( .DIN1(n1953), .DIN2(g5159), .Q(n1952) );
  xor2s3 U1268 ( .DIN1(g195), .DIN2(g1194), .Q(n1953) );
  nor2s3 U1269 ( .DIN1(n1954), .DIN2(n651), .Q(g5730) );
  nor2s3 U1270 ( .DIN1(n1955), .DIN2(g5158), .Q(n1954) );
  xor2s3 U1271 ( .DIN1(g186), .DIN2(g1198), .Q(n1955) );
  nnd2s3 U1272 ( .DIN1(n1956), .DIN2(n1957), .Q(g5187) );
  nnd3s3 U1273 ( .DIN1(n855), .DIN2(n837), .DIN3(n1415), .Q(n1957) );
  nnd2s3 U1274 ( .DIN1(n645), .DIN2(n646), .Q(n1956) );
  nnd2s3 U1275 ( .DIN1(n1958), .DIN2(n1959), .Q(g5186) );
  nnd2s3 U1276 ( .DIN1(g4668), .DIN2(n837), .Q(n1959) );
  nnd2s3 U1277 ( .DIN1(n1415), .DIN2(n645), .Q(n1958) );
  nnd3s3 U1278 ( .DIN1(n865), .DIN2(n837), .DIN3(n1960), .Q(g5185) );
  nnd2s3 U1279 ( .DIN1(n646), .DIN2(n855), .Q(n1960) );
  nnd2s3 U1280 ( .DIN1(n1961), .DIN2(n799), .Q(g5184) );
  xor2s3 U1281 ( .DIN1(n2271), .DIN2(n1936), .Q(n1961) );
  nnd2s3 U1282 ( .DIN1(n1962), .DIN2(n1963), .Q(g5183) );
  or3s3 U1283 ( .DIN1(g8219), .DIN2(n2272), .DIN3(n1936), .Q(n1963) );
  nnd2s3 U1284 ( .DIN1(n764), .DIN2(n774), .Q(n1962) );
  nnd2s3 U1285 ( .DIN1(n1964), .DIN2(n1965), .Q(g5182) );
  nnd4s2 U1286 ( .DIN1(n1458), .DIN2(n775), .DIN3(n774), .DIN4(n799), .Q(n1965) );
  nnd2s3 U1287 ( .DIN1(n2273), .DIN2(n764), .Q(n1964) );
  or3s3 U1288 ( .DIN1(n1458), .DIN2(n2272), .DIN3(n1936), .Q(g5181) );
  nor2s3 U1289 ( .DIN1(n2273), .DIN2(g8219), .Q(n1936) );
  nnd3s3 U1290 ( .DIN1(n2274), .DIN2(n2275), .DIN3(n2295), .Q(g5180) );
  and3s3 U1291 ( .DIN1(n699), .DIN2(n819), .DIN3(n1399), .Q(g5179) );
  nnd2s3 U1292 ( .DIN1(n1966), .DIN2(n1967), .Q(g5178) );
  nnd2s3 U1293 ( .DIN1(n1398), .DIN2(g8663), .Q(n1967) );
  or2s3 U1294 ( .DIN1(n2294), .DIN2(n2295), .Q(g8663) );
  nnd2s3 U1295 ( .DIN1(n699), .DIN2(g1724), .Q(n1966) );
  nnd3s3 U1296 ( .DIN1(n2276), .DIN2(n2277), .DIN3(n2294), .Q(g5177) );
  or5s3 U1297 ( .DIN1(n834), .DIN2(n839), .DIN3(n755), .DIN4(n769), .DIN5(
        n1968), .Q(g5175) );
  nnd4s2 U1298 ( .DIN1(n1482), .DIN2(n1506), .DIN3(n1480), .DIN4(n1492), .Q(
        n1968) );
  xor2s3 U1300 ( .DIN1(n739), .DIN2(n1494), .Q(n1969) );
  nnd4s2 U1302 ( .DIN1(n1396), .DIN2(\DFF_630/net855 ), .DIN3(n1456), .DIN4(
        n1970), .Q(g5172) );
  and3s3 U1303 ( .DIN1(\DFF_66/net291 ), .DIN2(\DFF_517/net742 ), .DIN3(
        \DFF_313/net538 ), .Q(n1970) );
  nor2s3 U1304 ( .DIN1(n1947), .DIN2(n1971), .Q(g5170) );
  nor2s3 U1305 ( .DIN1(n1972), .DIN2(n734), .Q(n1971) );
  nor2s3 U1306 ( .DIN1(n2280), .DIN2(g3857), .Q(n1972) );
  nor3s3 U1307 ( .DIN1(n2280), .DIN2(n2279), .DIN3(g3857), .Q(n1947) );
  xor2s3 U1308 ( .DIN1(n2280), .DIN2(g3857), .Q(g5169) );
  nor2s3 U1309 ( .DIN1(n1973), .DIN2(\DFF_391/net616 ), .Q(g5168) );
  nor2s3 U1310 ( .DIN1(n2293), .DIN2(n2292), .Q(n1973) );
  nor2s3 U1311 ( .DIN1(n717), .DIN2(n1974), .Q(g5167) );
  nor2s3 U1312 ( .DIN1(n1975), .DIN2(n716), .Q(n1974) );
  nor2s3 U1313 ( .DIN1(n2287), .DIN2(g3856), .Q(n1975) );
  or3s3 U1314 ( .DIN1(n2288), .DIN2(n2287), .DIN3(g3856), .Q(n1698) );
  xor2s3 U1315 ( .DIN1(n2287), .DIN2(g3856), .Q(g5166) );
  and3s3 U1316 ( .DIN1(n742), .DIN2(n859), .DIN3(n765), .Q(g5165) );
  nnd2s3 U1317 ( .DIN1(n1417), .DIN2(n766), .Q(n1706) );
  and3s3 U1318 ( .DIN1(n849), .DIN2(n766), .DIN3(n742), .Q(g5164) );
  nor2s3 U1319 ( .DIN1(n1457), .DIN2(n859), .Q(g5163) );
  and3s3 U1320 ( .DIN1(n865), .DIN2(n855), .DIN3(n1415), .Q(g4669) );
  and3s3 U1321 ( .DIN1(n1452), .DIN2(n646), .DIN3(n2282), .Q(g4668) );
  nnd2s3 U1322 ( .DIN1(n1399), .DIN2(n1976), .Q(g4665) );
  nnd2s3 U1323 ( .DIN1(n1398), .DIN2(n819), .Q(n1976) );
  nor2s3 U1324 ( .DIN1(g1401), .DIN2(\DFF_252/net477 ), .Q(g4664) );
  nor2s3 U1325 ( .DIN1(g1398), .DIN2(\DFF_218/net443 ), .Q(g4663) );
  nor2s3 U1326 ( .DIN1(g1395), .DIN2(\DFF_377/net602 ), .Q(g4661) );
  nor2s3 U1327 ( .DIN1(g1391), .DIN2(\DFF_402/net627 ), .Q(g4660) );
  nor6s3 U1328 ( .DIN1(n1977), .DIN2(n1978), .DIN3(n1979), .DIN4(n2286), 
        .DIN5(n2284), .DIN6(n2285), .Q(g4658) );
  nnd4s2 U1329 ( .DIN1(\DFF_635/net860 ), .DIN2(\DFF_422/net647 ), .DIN3(
        \DFF_63/net288 ), .DIN4(\DFF_412/net637 ), .Q(n1979) );
  nnd3s3 U1330 ( .DIN1(\DFF_518/net743 ), .DIN2(\DFF_527/net752 ), .DIN3(
        \DFF_140/net365 ), .Q(n1978) );
  nnd3s3 U1331 ( .DIN1(\DFF_260/net485 ), .DIN2(\DFF_24/net249 ), .DIN3(
        \DFF_180/net405 ), .Q(n1977) );
  nor6s3 U1332 ( .DIN1(n1980), .DIN2(n1981), .DIN3(n1982), .DIN4(n2291), 
        .DIN5(n2289), .DIN6(n2290), .Q(g4657) );
  nnd4s2 U1333 ( .DIN1(\DFF_564/net789 ), .DIN2(\DFF_84/net309 ), .DIN3(
        \DFF_200/net425 ), .DIN4(\DFF_314/net539 ), .Q(n1982) );
  nnd3s3 U1334 ( .DIN1(\DFF_155/net380 ), .DIN2(\DFF_597/net822 ), .DIN3(
        \DFF_619/net844 ), .Q(n1981) );
  nnd3s3 U1335 ( .DIN1(\DFF_521/net746 ), .DIN2(\DFF_101/net326 ), .DIN3(
        \DFF_20/net245 ), .Q(n1980) );
  nor2s3 U1336 ( .DIN1(g1269), .DIN2(g1268), .Q(g4656) );
  nnd2s3 U1337 ( .DIN1(n1427), .DIN2(n1983), .Q(g4655) );
  or2s3 U1338 ( .DIN1(n2293), .DIN2(n2292), .Q(n1983) );
  nnd2s3 U1339 ( .DIN1(n2292), .DIN2(n2293), .Q(n1427) );
  nor4s3 U1340 ( .DIN1(n1368), .DIN2(n875), .DIN3(n2101), .DIN4(n2052), .Q(
        g1015) );
  nor4s3 U1341 ( .DIN1(n1368), .DIN2(g6850), .DIN3(g6269), .DIN4(n2101), .Q(
        g1006) );
  or5s3 U1342 ( .DIN1(n663), .DIN2(n1984), .DIN3(n797), .DIN4(n778), .DIN5(
        n665), .Q(n1368) );
  nor2s3 U1343 ( .DIN1(n666), .DIN2(g7104), .Q(n1343) );
  and3s3 U1344 ( .DIN1(g43), .DIN2(g984), .DIN3(n1475), .Q(g7104) );
  nnd3s3 U1345 ( .DIN1(g43), .DIN2(g973), .DIN3(n667), .Q(n1239) );
  nnd3s3 U1346 ( .DIN1(g43), .DIN2(g976), .DIN3(n667), .Q(n1316) );
  or4s3 U1347 ( .DIN1(g962), .DIN2(g1871), .DIN3(g1870), .DIN4(n1985), .Q(
        n1984) );
  nnd4s2 U1348 ( .DIN1(\DFF_144/net369 ), .DIN2(\DFF_622/net847 ), .DIN3(
        \DFF_381/net606 ), .DIN4(\DFF_371/net596 ), .Q(n1985) );
  i1s3 U1349 ( .DIN(n963), .Q(n626) );
  i1s3 U1350 ( .DIN(n950), .Q(n627) );
  i1s3 U1351 ( .DIN(n927), .Q(n628) );
  i1s3 U1352 ( .DIN(n961), .Q(n629) );
  i1s3 U1353 ( .DIN(n948), .Q(n630) );
  i1s3 U1355 ( .DIN(n1017), .Q(n632) );
  i1s3 U1356 ( .DIN(n1021), .Q(n633) );
  i1s3 U1358 ( .DIN(n1018), .Q(n635) );
  i1s3 U1359 ( .DIN(n923), .Q(n636) );
  i1s3 U1360 ( .DIN(n920), .Q(n637) );
  i1s3 U1361 ( .DIN(n960), .Q(n638) );
  i1s3 U1362 ( .DIN(n949), .Q(n639) );
  i1s3 U1363 ( .DIN(n937), .Q(n640) );
  i1s3 U1364 ( .DIN(n945), .Q(n641) );
  i1s3 U1365 ( .DIN(n946), .Q(n642) );
  i1s3 U1366 ( .DIN(n1145), .Q(n643) );
  i1s3 U1367 ( .DIN(n1431), .Q(n644) );
  i1s3 U1368 ( .DIN(g5185), .Q(n645) );
  i1s3 U1369 ( .DIN(n1415), .Q(n646) );
  i1s3 U1370 ( .DIN(n2207), .Q(n647) );
  i1s3 U1371 ( .DIN(n2067), .Q(n648) );
  i1s3 U1372 ( .DIN(n1308), .Q(n649) );
  i1s3 U1373 ( .DIN(n1503), .Q(n650) );
  i1s3 U1374 ( .DIN(n2269), .Q(n651) );
  i1s3 U1375 ( .DIN(n1347), .Q(n652) );
  i1s3 U1376 ( .DIN(n2080), .Q(n653) );
  i1s3 U1377 ( .DIN(n1237), .Q(n654) );
  i1s3 U1378 ( .DIN(n1242), .Q(n655) );
  i1s3 U1379 ( .DIN(n1339), .Q(n656) );
  i1s3 U1380 ( .DIN(n1357), .Q(n657) );
  i1s3 U1381 ( .DIN(n1495), .Q(n658) );
  i1s3 U1382 ( .DIN(n1537), .Q(n659) );
  i1s3 U1383 ( .DIN(n1570), .Q(n660) );
  i1s3 U1384 ( .DIN(n1574), .Q(n661) );
  i1s3 U1385 ( .DIN(n2078), .Q(n662) );
  i1s3 U1386 ( .DIN(n1316), .Q(n663) );
  i1s3 U1387 ( .DIN(n1318), .Q(n664) );
  i1s3 U1388 ( .DIN(n1343), .Q(n665) );
  i1s3 U1389 ( .DIN(n1239), .Q(n666) );
  i1s3 U1390 ( .DIN(n1984), .Q(n667) );
  i1s3 U1391 ( .DIN(n2297), .Q(n668) );
  i1s3 U1392 ( .DIN(n2164), .Q(n669) );
  i1s3 U1393 ( .DIN(n2208), .Q(n670) );
  i1s3 U1394 ( .DIN(n1465), .Q(n671) );
  i1s3 U1395 ( .DIN(n2212), .Q(n672) );
  i1s3 U1396 ( .DIN(n1369), .Q(n673) );
  i1s3 U1397 ( .DIN(n2231), .Q(n674) );
  i1s3 U1398 ( .DIN(n2181), .Q(n675) );
  i1s3 U1399 ( .DIN(n2211), .Q(n676) );
  i1s3 U1400 ( .DIN(n2228), .Q(n677) );
  i1s3 U1401 ( .DIN(n1313), .Q(n678) );
  i1s3 U1402 ( .DIN(n1407), .Q(n679) );
  i1s3 U1403 ( .DIN(n2227), .Q(n680) );
  i1s3 U1404 ( .DIN(n2189), .Q(n681) );
  i1s3 U1405 ( .DIN(n2097), .Q(n682) );
  i1s3 U1406 ( .DIN(n1459), .Q(n683) );
  i1s3 U1407 ( .DIN(n2174), .Q(n684) );
  i1s3 U1408 ( .DIN(n1453), .Q(n685) );
  i1s3 U1409 ( .DIN(n2196), .Q(n686) );
  i1s3 U1410 ( .DIN(n1429), .Q(n687) );
  i1s3 U1411 ( .DIN(n1550), .Q(n688) );
  i1s3 U1412 ( .DIN(n1530), .Q(n689) );
  i1s3 U1413 ( .DIN(n1489), .Q(n690) );
  i1s3 U1414 ( .DIN(n1411), .Q(n691) );
  i1s3 U1415 ( .DIN(n1461), .Q(n692) );
  i1s3 U1416 ( .DIN(n2085), .Q(n693) );
  i1s3 U1417 ( .DIN(n2151), .Q(n694) );
  i1s3 U1418 ( .DIN(g999), .Q(n695) );
  i1s3 U1419 ( .DIN(n1811), .Q(n696) );
  i1s3 U1420 ( .DIN(n2194), .Q(n697) );
  i1s3 U1421 ( .DIN(n1419), .Q(n698) );
  i1s3 U1422 ( .DIN(n1398), .Q(n699) );
  i1s3 U1423 ( .DIN(n895), .Q(n700) );
  i1s3 U1424 ( .DIN(n1724), .Q(n701) );
  i1s3 U1425 ( .DIN(n1674), .Q(n702) );
  i1s3 U1426 ( .DIN(n1492), .Q(n703) );
  i1s3 U1427 ( .DIN(n2161), .Q(n704) );
  i1s3 U1428 ( .DIN(n2059), .Q(n705) );
  i1s3 U1429 ( .DIN(n2036), .Q(n706) );
  i1s3 U1430 ( .DIN(n1531), .Q(n707) );
  i1s3 U1431 ( .DIN(n1786), .Q(n708) );
  i1s3 U1432 ( .DIN(n1494), .Q(n709) );
  i1s3 U1433 ( .DIN(n2236), .Q(n710) );
  i1s3 U1434 ( .DIN(n1176), .Q(n711) );
  i1s3 U1435 ( .DIN(n1183), .Q(n712) );
  i1s3 U1436 ( .DIN(n1182), .Q(n713) );
  i1s3 U1437 ( .DIN(n1462), .Q(n714) );
  i1s3 U1438 ( .DIN(n2209), .Q(n715) );
  i1s3 U1439 ( .DIN(n2288), .Q(n716) );
  i1s3 U1440 ( .DIN(n1698), .Q(n717) );
  i1s3 U1441 ( .DIN(n2213), .Q(n718) );
  i1s3 U1443 ( .DIN(n2038), .Q(n720) );
  i1s3 U1444 ( .DIN(n2200), .Q(n721) );
  i1s3 U1445 ( .DIN(n1402), .Q(n722) );
  i1s3 U1446 ( .DIN(n1445), .Q(n723) );
  i1s3 U1447 ( .DIN(n2029), .Q(n724) );
  i1s3 U1448 ( .DIN(g9132), .Q(n725) );
  i1s3 U1449 ( .DIN(n1480), .Q(n726) );
  i1s3 U1450 ( .DIN(n2198), .Q(n727) );
  i1s3 U1451 ( .DIN(n1506), .Q(n728) );
  i1s3 U1452 ( .DIN(n2073), .Q(n729) );
  i1s3 U1453 ( .DIN(n1440), .Q(n730) );
  i1s3 U1454 ( .DIN(n1541), .Q(n731) );
  i1s3 U1455 ( .DIN(n2091), .Q(n732) );
  i1s3 U1456 ( .DIN(n2075), .Q(n733) );
  i1s3 U1457 ( .DIN(n2279), .Q(n734) );
  i1s3 U1458 ( .DIN(g4655), .Q(n735) );
  i1s3 U1459 ( .DIN(n1427), .Q(n736) );
  i1s3 U1460 ( .DIN(n2301), .Q(n737) );
  i1s3 U1461 ( .DIN(n2238), .Q(n738) );
  i1s3 U1462 ( .DIN(n1513), .Q(n739) );
  i1s3 U1463 ( .DIN(n2216), .Q(n740) );
  i1s3 U1464 ( .DIN(n2037), .Q(n741) );
  i1s3 U1465 ( .DIN(n1405), .Q(n742) );
  i1s3 U1466 ( .DIN(n1470), .Q(n743) );
  i1s3 U1467 ( .DIN(n2094), .Q(n744) );
  i1s3 U1468 ( .DIN(n1396), .Q(n745) );
  i1s3 U1469 ( .DIN(n1482), .Q(n746) );
  i1s3 U1470 ( .DIN(n1394), .Q(n747) );
  i1s3 U1471 ( .DIN(n2223), .Q(n748) );
  i1s3 U1472 ( .DIN(n2199), .Q(n749) );
  i1s3 U1473 ( .DIN(n2082), .Q(n750) );
  i1s3 U1474 ( .DIN(n2063), .Q(n751) );
  i1s3 U1475 ( .DIN(n2046), .Q(n752) );
  i1s3 U1476 ( .DIN(n2243), .Q(n753) );
  i1s3 U1477 ( .DIN(n2242), .Q(n754) );
  i1s3 U1478 ( .DIN(n1488), .Q(n755) );
  i1s3 U1479 ( .DIN(n2268), .Q(n756) );
  i1s3 U1480 ( .DIN(n2071), .Q(n757) );
  i1s3 U1481 ( .DIN(n1423), .Q(n758) );
  i1s3 U1482 ( .DIN(n2088), .Q(n759) );
  i1s3 U1483 ( .DIN(n1725), .Q(n760) );
  i1s3 U1484 ( .DIN(n1484), .Q(n761) );
  i1s3 U1486 ( .DIN(n1468), .Q(n763) );
  i1s3 U1487 ( .DIN(g5181), .Q(n764) );
  i1s3 U1488 ( .DIN(n1706), .Q(n765) );
  i1s3 U1489 ( .DIN(n1432), .Q(n766) );
  i1s3 U1490 ( .DIN(n1511), .Q(n767) );
  i1s3 U1491 ( .DIN(n2098), .Q(n768) );
  i1s3 U1492 ( .DIN(n1508), .Q(n769) );
  i1s3 U1493 ( .DIN(n2188), .Q(n770) );
  i1s3 U1496 ( .DIN(n1449), .Q(n773) );
  i1s3 U1497 ( .DIN(n2273), .Q(n774) );
  i1s3 U1498 ( .DIN(n1936), .Q(n775) );
  i1s3 U1499 ( .DIN(n2131), .Q(n776) );
  i1s3 U1500 ( .DIN(n2264), .Q(n777) );
  i1s3 U1501 ( .DIN(n1475), .Q(n778) );
  i1s3 U1502 ( .DIN(n2195), .Q(n779) );
  i1s3 U1503 ( .DIN(n1397), .Q(n780) );
  i1s3 U1504 ( .DIN(n2030), .Q(n781) );
  i1s3 U1505 ( .DIN(n2225), .Q(n782) );
  i1s3 U1506 ( .DIN(n2237), .Q(n783) );
  i1s3 U1507 ( .DIN(n2047), .Q(n784) );
  i1s3 U1508 ( .DIN(n2229), .Q(n785) );
  i1s3 U1509 ( .DIN(n1391), .Q(n786) );
  i1s3 U1510 ( .DIN(n1598), .Q(n787) );
  i1s3 U1511 ( .DIN(n2205), .Q(n788) );
  i1s3 U1512 ( .DIN(n2193), .Q(n789) );
  i1s3 U1513 ( .DIN(n2179), .Q(n790) );
  i1s3 U1514 ( .DIN(n2081), .Q(n791) );
  i1s3 U1515 ( .DIN(n919), .Q(n792) );
  i1s3 U1516 ( .DIN(n1496), .Q(n793) );
  i1s3 U1518 ( .DIN(n2042), .Q(n795) );
  i1s3 U1519 ( .DIN(n1481), .Q(n796) );
  i1s3 U1520 ( .DIN(n1401), .Q(n797) );
  i1s3 U1521 ( .DIN(n2214), .Q(n798) );
  i1s3 U1522 ( .DIN(n2272), .Q(n799) );
  i1s3 U1523 ( .DIN(n2197), .Q(n800) );
  i1s3 U1524 ( .DIN(n1469), .Q(n801) );
  i1s3 U1525 ( .DIN(n1473), .Q(n802) );
  i1s3 U1526 ( .DIN(n1409), .Q(n803) );
  i1s3 U1527 ( .DIN(n2178), .Q(n804) );
  i1s3 U1528 ( .DIN(n1502), .Q(n805) );
  i1s3 U1529 ( .DIN(n2192), .Q(n806) );
  i1s3 U1530 ( .DIN(n2230), .Q(n807) );
  i1s3 U1531 ( .DIN(n2086), .Q(n808) );
  i1s3 U1532 ( .DIN(n2074), .Q(n809) );
  i1s3 U1533 ( .DIN(n2175), .Q(n810) );
  i1s3 U1534 ( .DIN(n2224), .Q(n811) );
  i1s3 U1535 ( .DIN(n2191), .Q(n812) );
  i1s3 U1536 ( .DIN(n2093), .Q(n813) );
  i1s3 U1537 ( .DIN(n2070), .Q(n814) );
  i1s3 U1538 ( .DIN(n2215), .Q(n815) );
  i1s3 U1539 ( .DIN(n2172), .Q(n816) );
  i1s3 U1540 ( .DIN(n2190), .Q(n817) );
  i1s3 U1541 ( .DIN(n2173), .Q(n818) );
  i1s3 U1542 ( .DIN(n2283), .Q(n819) );
  i1s3 U1543 ( .DIN(n2204), .Q(n820) );
  i1s3 U1544 ( .DIN(n2201), .Q(n821) );
  i1s3 U1545 ( .DIN(n2064), .Q(n822) );
  i1s3 U1546 ( .DIN(n1433), .Q(n823) );
  i1s3 U1547 ( .DIN(n2055), .Q(n824) );
  i1s3 U1548 ( .DIN(n1390), .Q(n825) );
  i1s3 U1549 ( .DIN(n2083), .Q(n826) );
  i1s3 U1550 ( .DIN(n1486), .Q(n827) );
  i1s3 U1551 ( .DIN(n2244), .Q(n828) );
  i1s3 U1552 ( .DIN(n2180), .Q(n829) );
  i1s3 U1553 ( .DIN(n1403), .Q(n830) );
  i1s3 U1554 ( .DIN(n2053), .Q(n831) );
  i1s3 U1556 ( .DIN(n2239), .Q(n833) );
  i1s3 U1557 ( .DIN(n1490), .Q(n834) );
  i1s3 U1558 ( .DIN(n2203), .Q(n835) );
  i1s3 U1559 ( .DIN(n2154), .Q(n836) );
  i1s3 U1560 ( .DIN(n2270), .Q(n837) );
  i1s3 U1561 ( .DIN(n1460), .Q(n838) );
  i1s3 U1562 ( .DIN(n1477), .Q(n839) );
  i1s3 U1563 ( .DIN(n2060), .Q(n840) );
  i1s3 U1564 ( .DIN(n2048), .Q(n841) );
  i1s3 U1565 ( .DIN(n2218), .Q(n842) );
  i1s3 U1567 ( .DIN(n2241), .Q(n844) );
  i1s3 U1568 ( .DIN(n1454), .Q(n845) );
  i1s3 U1569 ( .DIN(n2051), .Q(n846) );
  i1s3 U1570 ( .DIN(n2210), .Q(n847) );
  i1s3 U1571 ( .DIN(n2217), .Q(n848) );
  i1s3 U1572 ( .DIN(n1417), .Q(n849) );
  i1s3 U1573 ( .DIN(n2077), .Q(n850) );
  i1s3 U1574 ( .DIN(n1446), .Q(n851) );
  i1s3 U1575 ( .DIN(n2226), .Q(n852) );
  i1s3 U1576 ( .DIN(n1996), .Q(n853) );
  i1s3 U1578 ( .DIN(n2282), .Q(n855) );
  i1s3 U1579 ( .DIN(n2090), .Q(n856) );
  i1s3 U1580 ( .DIN(n2202), .Q(n857) );
  i1s3 U1581 ( .DIN(n2076), .Q(n858) );
  i1s3 U1582 ( .DIN(n2281), .Q(n859) );
  i1s3 U1584 ( .DIN(n2263), .Q(n861) );
  i1s3 U1585 ( .DIN(n2235), .Q(n862) );
  i1s3 U1586 ( .DIN(n1421), .Q(n863) );
  i1s3 U1587 ( .DIN(n1463), .Q(n864) );
  i1s3 U1588 ( .DIN(n1452), .Q(n865) );
  i1s3 U1589 ( .DIN(n1444), .Q(n866) );
  i1s3 U1590 ( .DIN(n2068), .Q(n867) );
  i1s3 U1591 ( .DIN(n2240), .Q(n868) );
  i1s3 U1592 ( .DIN(n1422), .Q(n869) );
  i1s3 U1593 ( .DIN(n1395), .Q(n870) );
  i1s3 U1594 ( .DIN(n2206), .Q(n871) );
  i1s3 U1595 ( .DIN(n2130), .Q(n872) );
  i1s3 U1596 ( .DIN(n2222), .Q(n873) );
  i1s3 U1597 ( .DIN(n1441), .Q(n874) );
  i1s3 U1598 ( .DIN(g6289), .Q(n875) );
  i1s3 U1599 ( .DIN(g6291), .Q(n876) );
  i1s3 U1600 ( .DIN(g6303), .Q(n877) );
  i1s3 U1601 ( .DIN(g43), .Q(g6850) );
  i1s3 U1602 ( .DIN(g6307), .Q(n879) );
  i1s3 U1603 ( .DIN(n1549), .Q(n880) );
  i1s3 U1604 ( .DIN(g6308), .Q(n881) );
  i1s3 U1605 ( .DIN(g647), .Q(n882) );
  i1s3 U1606 ( .DIN(g648), .Q(n883) );
  i1s3 U1607 ( .DIN(g690), .Q(n884) );
  i1s3 U1608 ( .DIN(g694), .Q(n885) );
  i1s3 U1609 ( .DIN(g698), .Q(n886) );
  i1s3 U1610 ( .DIN(g702), .Q(n887) );
  i1s3 U1611 ( .DIN(g722), .Q(n888) );
  i1s3 U1612 ( .DIN(g723), .Q(n889) );
  i1s3 U1613 ( .DIN(g795), .Q(g3854) );
  i1s3 U1614 ( .DIN(g929), .Q(g3856) );
  i1s3 U1615 ( .DIN(g955), .Q(g3857) );
  and2s1 U1616 ( .DIN1(g751), .DIN2(n947), .Q(n941) );
  nnd2s1 U1617 ( .DIN1(g752), .DIN2(n947), .Q(n1043) );
  nnd2s1 U1618 ( .DIN1(g753), .DIN2(n947), .Q(n1081) );
  and2s1 U1619 ( .DIN1(g755), .DIN2(n947), .Q(n971) );
  and2s1 U1620 ( .DIN1(g754), .DIN2(n947), .Q(n995) );
  nnd2s2 U1621 ( .DIN1(g756), .DIN2(n947), .Q(n1105) );
  nnd2s2 U1622 ( .DIN1(g757), .DIN2(n947), .Q(n1147) );
  nnd2s2 U1623 ( .DIN1(g5729), .DIN2(n947), .Q(n1199) );
  nnd2s1 U1624 ( .DIN1(n1400), .DIN2(n1637), .Q(g7300) );
  nnd2s1 U1625 ( .DIN1(n1400), .DIN2(n1676), .Q(g7109) );
  nnd2s1 U1626 ( .DIN1(n1400), .DIN2(n1677), .Q(g7108) );
  nnd2s2 U1627 ( .DIN1(n1400), .DIN2(n1722), .Q(g6859) );
  nnd2s2 U1628 ( .DIN1(n1400), .DIN2(n1727), .Q(g6858) );
  nnd2s2 U1629 ( .DIN1(n1400), .DIN2(n1730), .Q(g6857) );
  nnd2s2 U1630 ( .DIN1(n1400), .DIN2(n1784), .Q(g6379) );
  nnd2s2 U1631 ( .DIN1(n1400), .DIN2(n1788), .Q(g6378) );
  nnd2s2 U1632 ( .DIN1(n1400), .DIN2(n1789), .Q(g6377) );
  nnd2s2 U1633 ( .DIN1(n1969), .DIN2(n1400), .Q(g5174) );
  and4s1 U1634 ( .DIN1(n1400), .DIN2(n1673), .DIN3(n1639), .DIN4(n756), .Q(
        g7110) );
  nnd2s2 U1635 ( .DIN1(n1400), .DIN2(n761), .Q(n1945) );
  nnd2s2 U1636 ( .DIN1(n1400), .DIN2(n739), .Q(g5173) );
  nnd2s1 U1637 ( .DIN1(n1441), .DIN2(n1238), .Q(n1585) );
  nnd3s1 U1638 ( .DIN1(n1238), .DIN2(n655), .DIN3(n1440), .Q(n1241) );
  nnd3s1 U1639 ( .DIN1(n1238), .DIN2(n656), .DIN3(n1459), .Q(n1338) );
  nnd3s1 U1640 ( .DIN1(n1238), .DIN2(n658), .DIN3(n1460), .Q(n1493) );
  nnd3s2 U1641 ( .DIN1(n1238), .DIN2(n660), .DIN3(n1462), .Q(n1566) );
  nnd3s2 U1642 ( .DIN1(n1238), .DIN2(n874), .DIN3(n1461), .Q(n1578) );
  nnd3s2 U1643 ( .DIN1(n657), .DIN2(n1339), .DIN3(n1238), .Q(n1355) );
  nnd3s2 U1644 ( .DIN1(n659), .DIN2(n1495), .DIN3(n1238), .Q(n1535) );
  nnd3s2 U1645 ( .DIN1(n661), .DIN2(n1570), .DIN3(n1238), .Q(n1569) );
  nnd4s1 U1646 ( .DIN1(n1238), .DIN2(n656), .DIN3(n1242), .DIN4(n683), .Q(
        n1312) );
  nnd4s1 U1647 ( .DIN1(n1238), .DIN2(n658), .DIN3(n1357), .DIN4(n838), .Q(
        n1392) );
  nnd4s1 U1648 ( .DIN1(n1238), .DIN2(n1574), .DIN3(n874), .DIN4(n692), .Q(
        n1573) );
  nnd4s1 U1649 ( .DIN1(n1238), .DIN2(n660), .DIN3(n1537), .DIN4(n714), .Q(
        n1587) );
  and3s1 U1650 ( .DIN1(n655), .DIN2(n730), .DIN3(n1238), .Q(n1231) );
  nnd2s1 U1651 ( .DIN1(n1504), .DIN2(n1611), .Q(n1610) );
  nnd2s1 U1652 ( .DIN1(n1504), .DIN2(n1651), .Q(n1650) );
  nnd2s1 U1653 ( .DIN1(n1504), .DIN2(n1941), .Q(n1940) );
  nnd2s1 U1654 ( .DIN1(n2260), .DIN2(n1504), .Q(n1942) );
  nnd2s1 U1655 ( .DIN1(n1622), .DIN2(n1504), .Q(n1621) );
  nnd2s1 U1656 ( .DIN1(n1626), .DIN2(n1504), .Q(n1625) );
  nnd2s1 U1657 ( .DIN1(n1655), .DIN2(n1504), .Q(n1654) );
  nnd2s2 U1658 ( .DIN1(n1663), .DIN2(n1504), .Q(n1662) );
  nnd2s2 U1659 ( .DIN1(n1667), .DIN2(n1504), .Q(n1666) );
  nnd3s2 U1660 ( .DIN1(n1617), .DIN2(n1612), .DIN3(n1504), .Q(n1616) );
  nnd3s2 U1661 ( .DIN1(n1646), .DIN2(n1623), .DIN3(n1504), .Q(n1645) );
  nnd3s2 U1662 ( .DIN1(n1658), .DIN2(n1652), .DIN3(n1504), .Q(n1657) );
  nnd3s2 U1663 ( .DIN1(n1720), .DIN2(n1664), .DIN3(n1504), .Q(n1719) );
  i1s3 U1664 ( .DIN(n1504), .Q(n719) );
  hi1s1 U1665 ( .DIN(n2302), .Q(n2303) );
  i1s3 U1666 ( .DIN(n2303), .Q(n2304) );
  ib1s9 U1667 ( .DIN(n2310), .Q(n2307) );
  ib1s9 U1668 ( .DIN(n2310), .Q(n2308) );
  ib1s5 U1669 ( .DIN(n1413), .Q(n860) );
  ib1s5 U1670 ( .DIN(n1412), .Q(n854) );
  ib1s5 U1671 ( .DIN(n1428), .Q(n843) );
  ib1s5 U1672 ( .DIN(n1855), .Q(n832) );
  ib1s5 U1673 ( .DIN(n1828), .Q(n794) );
  ib1s5 U1674 ( .DIN(n1414), .Q(n772) );
  ib1s5 U1675 ( .DIN(n1909), .Q(n771) );
  ib1s5 U1676 ( .DIN(n1882), .Q(n762) );
  ib1s5 U1677 ( .DIN(n1019), .Q(n634) );
  ib1s5 U1678 ( .DIN(n1020), .Q(n631) );
  and3s3 U1679 ( .DIN1(n1259), .DIN2(n786), .DIN3(n1185), .Q(n2305) );
  and3s3 U1680 ( .DIN1(n1259), .DIN2(n786), .DIN3(n1185), .Q(n2306) );
  i1s12 U1681 ( .DIN(n2310), .Q(n2309) );
  i1s12 U1682 ( .DIN(n633), .Q(n2310) );
  sdffs1 \DFF_637/Q_reg  ( .DIN(n843), .SDIN(g12), .SSEL(test_se), .CLK(CK), 
        .Q(test_so), .QN(n1431) );
  sdffs1 \DFF_636/Q_reg  ( .DIN(g7048), .SDIN(n2638), .SSEL(test_se), .CLK(CK), 
        .Q(g12) );
  sdffs1 \DFF_635/Q_reg  ( .DIN(g6879), .SDIN(n2637), .SSEL(test_se), .CLK(CK), 
        .Q(n2638), .QN(\DFF_635/net860 ) );
  sdffs1 \DFF_634/Q_reg  ( .DIN(g4373), .SDIN(g5158), .SSEL(test_se), .CLK(CK), 
        .Q(n2637), .QN(n1456) );
  sdffs1 \DFF_633/Q_reg  ( .DIN(g5730), .SDIN(n2636), .SSEL(test_se), .CLK(CK), 
        .Q(g5158) );
  sdffs1 \DFF_632/Q_reg  ( .DIN(g5186), .SDIN(n2635), .SSEL(test_se), .CLK(CK), 
        .Q(n2636), .QN(n1415) );
  sdffs1 \DFF_631/Q_reg  ( .DIN(g8676), .SDIN(g4370), .SSEL(test_se), .CLK(CK), 
        .Q(n2635), .QN(n2167) );
  sdffs1 \DFF_630/Q_reg  ( .DIN(g4371), .SDIN(n2634), .SSEL(test_se), .CLK(CK), 
        .Q(g4370), .QN(\DFF_630/net855 ) );
  sdffs1 \DFF_629/Q_reg  ( .DIN(g6351), .SDIN(n2633), .SSEL(test_se), .CLK(CK), 
        .Q(n2634), .QN(n2207) );
  sdffs1 \DFF_628/Q_reg  ( .DIN(g7771), .SDIN(n2632), .SSEL(test_se), .CLK(CK), 
        .Q(n2633), .QN(n2067) );
  sdffs1 \DFF_627/Q_reg  ( .DIN(g6843), .SDIN(n2631), .SSEL(test_se), .CLK(CK), 
        .Q(n2632), .QN(n2122) );
  sdffs1 \DFF_626/Q_reg  ( .DIN(g5742), .SDIN(n2269), .SSEL(test_se), .CLK(CK), 
        .Q(n2631), .QN(n2260) );
  sdffs1 \DFF_625/Q_reg  ( .DIN(g201), .SDIN(n2630), .SSEL(test_se), .CLK(CK), 
        .Q(n2269) );
  sdffs1 \DFF_624/Q_reg  ( .DIN(g7517), .SDIN(n2629), .SSEL(test_se), .CLK(CK), 
        .Q(n2630), .QN(n2080) );
  sdffs1 \DFF_623/Q_reg  ( .DIN(g7523), .SDIN(n2628), .SSEL(test_se), .CLK(CK), 
        .Q(n2629), .QN(n2078) );
  sdffs1 \DFF_622/Q_reg  ( .DIN(g1870), .SDIN(g435), .SSEL(test_se), .CLK(CK), 
        .Q(n2628), .QN(\DFF_622/net847 ) );
  sdffs1 \DFF_621/Q_reg  ( .DIN(g4650), .SDIN(n2627), .SSEL(test_se), .CLK(CK), 
        .Q(g435) );
  sdffs1 \DFF_620/Q_reg  ( .DIN(g7739), .SDIN(n2626), .SSEL(test_se), .CLK(CK), 
        .Q(n2627), .QN(n2278) );
  sdffs1 \DFF_619/Q_reg  ( .DIN(g6870), .SDIN(n2625), .SSEL(test_se), .CLK(CK), 
        .Q(n2626), .QN(\DFF_619/net844 ) );
  sdffs1 \DFF_618/Q_reg  ( .DIN(n2304), .SDIN(n2624), .SSEL(test_se), .CLK(CK), 
        .Q(n2625), .QN(n2128) );
  sdffs1 \DFF_617/Q_reg  ( .DIN(g7530), .SDIN(n2623), .SSEL(test_se), .CLK(CK), 
        .Q(n2624), .QN(n2164) );
  sdffs1 \DFF_615/Q_reg  ( .DIN(g6338), .SDIN(n2095), .SSEL(test_se), .CLK(CK), 
        .Q(n2623), .QN(n2220) );
  sdffs1 \DFF_614/Q_reg  ( .DIN(g7117), .SDIN(n2622), .SSEL(test_se), .CLK(CK), 
        .Q(n2095) );
  sdffs1 \DFF_613/Q_reg  ( .DIN(g6350), .SDIN(n2621), .SSEL(test_se), .CLK(CK), 
        .Q(n2622), .QN(n2208) );
  sdffs1 \DFF_612/Q_reg  ( .DIN(g9096), .SDIN(n2620), .SSEL(test_se), .CLK(CK), 
        .Q(n2621), .QN(n2024) );
  sdffs1 \DFF_611/Q_reg  ( .DIN(g6339), .SDIN(g3848), .SSEL(test_se), .CLK(CK), 
        .Q(n2620), .QN(n2219) );
  sdffs1 \DFF_610/Q_reg  ( .DIN(g7303), .SDIN(g1204), .SSEL(test_se), .CLK(CK), 
        .Q(g3848), .QN(n2261) );
  sdffs1 \DFF_609/Q_reg  ( .DIN(g1203), .SDIN(n2619), .SSEL(test_se), .CLK(CK), 
        .Q(g1204) );
  sdffs1 \DFF_608/Q_reg  ( .DIN(g5163), .SDIN(n2618), .SSEL(test_se), .CLK(CK), 
        .Q(n2619), .QN(n1465) );
  sdffs1 \DFF_607/Q_reg  ( .DIN(g6346), .SDIN(g162), .SSEL(test_se), .CLK(CK), 
        .Q(n2618), .QN(n2212) );
  sdffs1 \DFF_606/Q_reg  ( .DIN(g162), .SDIN(n2617), .SSEL(test_se), .CLK(CK), 
        .Q(g162), .QN(n2101) );
  sdffs1 \DFF_605/Q_reg  ( .DIN(g8671), .SDIN(n2616), .SSEL(test_se), .CLK(CK), 
        .Q(n2617), .QN(\DFF_605/net830 ) );
  sdffs1 \DFF_604/Q_reg  ( .DIN(g6327), .SDIN(n2615), .SSEL(test_se), .CLK(CK), 
        .Q(n2616), .QN(n2231) );
  sdffs1 \DFF_603/Q_reg  ( .DIN(n843), .SDIN(g673), .SSEL(test_se), .CLK(CK), 
        .Q(n2615), .QN(n2127) );
  sdffs1 \DFF_602/Q_reg  ( .DIN(g673), .SDIN(n2285), .SSEL(test_se), .CLK(CK), 
        .Q(g673), .QN(n2181) );
  sdffs1 \DFF_601/Q_reg  ( .DIN(g6886), .SDIN(g3852), .SSEL(test_se), .CLK(CK), 
        .Q(n2285) );
  sdffs1 \DFF_599/Q_reg  ( .DIN(g7301), .SDIN(g94), .SSEL(test_se), .CLK(CK), 
        .Q(g3852), .QN(n2267) );
  sdffs1 \DFF_598/Q_reg  ( .DIN(n2304), .SDIN(n2614), .SSEL(test_se), .CLK(CK), 
        .Q(g94) );
  sdffs1 \DFF_597/Q_reg  ( .DIN(g6872), .SDIN(n2613), .SSEL(test_se), .CLK(CK), 
        .Q(n2614), .QN(\DFF_597/net822 ) );
  sdffs1 \DFF_596/Q_reg  ( .DIN(g6347), .SDIN(g1311), .SSEL(test_se), .CLK(CK), 
        .Q(n2613), .QN(n2211) );
  sdffs1 \DFF_595/Q_reg  ( .DIN(g1310), .SDIN(n2612), .SSEL(test_se), .CLK(CK), 
        .Q(g1311) );
  sdffs1 \DFF_594/Q_reg  ( .DIN(g6330), .SDIN(n2611), .SSEL(test_se), .CLK(CK), 
        .Q(n2612), .QN(n2228) );
  sdffs1 \DFF_593/Q_reg  ( .DIN(g1159), .SDIN(n2610), .SSEL(test_se), .CLK(CK), 
        .Q(n2611), .QN(n1407) );
  sdffs1 \DFF_592/Q_reg  ( .DIN(g9108), .SDIN(n2609), .SSEL(test_se), .CLK(CK), 
        .Q(n2610), .QN(n2012) );
  sdffs1 \DFF_591/Q_reg  ( .DIN(g6331), .SDIN(g539), .SSEL(test_se), .CLK(CK), 
        .Q(n2609), .QN(n2227) );
  sdffs1 \DFF_590/Q_reg  ( .DIN(g3845), .SDIN(n2608), .SSEL(test_se), .CLK(CK), 
        .Q(g539) );
  sdffs1 \DFF_589/Q_reg  ( .DIN(g6369), .SDIN(n2607), .SSEL(test_se), .CLK(CK), 
        .Q(n2608), .QN(n2189) );
  sdffs1 \DFF_588/Q_reg  ( .DIN(g8227), .SDIN(g1253), .SSEL(test_se), .CLK(CK), 
        .Q(n2607), .QN(n1451) );
  sdffs1 \DFF_587/Q_reg  ( .DIN(n2298), .SDIN(n2097), .SSEL(test_se), .CLK(CK), 
        .Q(g1253) );
  sdffs1 \DFF_586/Q_reg  ( .DIN(g7115), .SDIN(g1393), .SSEL(test_se), .CLK(CK), 
        .Q(n2097) );
  sdffs1 \DFF_584/Q_reg  ( .DIN(g7505), .SDIN(g1193), .SSEL(test_se), .CLK(CK), 
        .Q(g1393) );
  sdffs1 \DFF_583/Q_reg  ( .DIN(g1192), .SDIN(g973), .SSEL(test_se), .CLK(CK), 
        .Q(g1193) );
  sdffs1 \DFF_582/Q_reg  ( .DIN(g8672), .SDIN(n2606), .SSEL(test_se), .CLK(CK), 
        .Q(g973) );
  sdffs1 \DFF_581/Q_reg  ( .DIN(g8959), .SDIN(g376), .SSEL(test_se), .CLK(CK), 
        .Q(n2606), .QN(n1459) );
  sdffs1 \DFF_580/Q_reg  ( .DIN(g4642), .SDIN(g677), .SSEL(test_se), .CLK(CK), 
        .Q(g376) );
  sdffs1 \DFF_579/Q_reg  ( .DIN(g677), .SDIN(n2290), .SSEL(test_se), .CLK(CK), 
        .Q(g677), .QN(n2174) );
  sdffs1 \DFF_578/Q_reg  ( .DIN(g6873), .SDIN(n2605), .SSEL(test_se), .CLK(CK), 
        .Q(n2290) );
  sdffs1 \DFF_577/Q_reg  ( .DIN(g6861), .SDIN(g7423), .SSEL(test_se), .CLK(CK), 
        .Q(n2605), .QN(n1474) );
  sdffs1 \DFF_576/Q_reg  ( .DIN(g7424), .SDIN(n2604), .SSEL(test_se), .CLK(CK), 
        .Q(g7423) );
  sdffs1 \DFF_575/Q_reg  ( .DIN(g7766), .SDIN(n2603), .SSEL(test_se), .CLK(CK), 
        .Q(n2604), .QN(n1453) );
  sdffs1 \DFF_574/Q_reg  ( .DIN(n1384), .SDIN(n2602), .SSEL(test_se), .CLK(CK), 
        .Q(n2603), .QN(n2149) );
  sdffs1 \DFF_573/Q_reg  ( .DIN(g6325), .SDIN(n2601), .SSEL(test_se), .CLK(CK), 
        .Q(n2602), .QN(n2233) );
  sdffs1 \DFF_572/Q_reg  ( .DIN(g6362), .SDIN(n2600), .SSEL(test_se), .CLK(CK), 
        .Q(n2601), .QN(n2196) );
  sdffs1 \DFF_571/Q_reg  ( .DIN(g9088), .SDIN(n1387), .SSEL(test_se), .CLK(CK), 
        .Q(n2600), .QN(n2032) );
  sdffs1 \DFF_570/Q_reg  ( .DIN(g9375), .SDIN(g2661), .SSEL(test_se), .CLK(CK), 
        .Q(n1387), .QN(n1429) );
  sdffs1 \DFF_569/Q_reg  ( .DIN(g6382), .SDIN(g1155), .SSEL(test_se), .CLK(CK), 
        .Q(g2661), .QN(g3863) );
  sdffs1 \DFF_568/Q_reg  ( .DIN(g1154), .SDIN(n2599), .SSEL(test_se), .CLK(CK), 
        .Q(g1155) );
  sdffs1 \DFF_567/Q_reg  ( .DIN(g7529), .SDIN(n2598), .SSEL(test_se), .CLK(CK), 
        .Q(n2599), .QN(n1424) );
  sdffs1 \DFF_566/Q_reg  ( .DIN(g1147), .SDIN(n2597), .SSEL(test_se), .CLK(CK), 
        .Q(n2598), .QN(n2134) );
  sdffs1 \DFF_565/Q_reg  ( .DIN(g9099), .SDIN(n2596), .SSEL(test_se), .CLK(CK), 
        .Q(n2597), .QN(n2021) );
  sdffs1 \DFF_564/Q_reg  ( .DIN(g6866), .SDIN(n2595), .SSEL(test_se), .CLK(CK), 
        .Q(n2596), .QN(\DFF_564/net789 ) );
  sdffs1 \DFF_563/Q_reg  ( .DIN(g9109), .SDIN(n2069), .SSEL(test_se), .CLK(CK), 
        .Q(n2595), .QN(n2011) );
  sdffs1 \DFF_562/Q_reg  ( .DIN(g7423), .SDIN(g5150), .SSEL(test_se), .CLK(CK), 
        .Q(n2069) );
  sdffs1 \DFF_561/Q_reg  ( .DIN(n772), .SDIN(g5153), .SSEL(test_se), .CLK(CK), 
        .Q(g5150), .QN(n1995) );
  sdffs1 \DFF_560/Q_reg  ( .DIN(g6841), .SDIN(n2594), .SSEL(test_se), .CLK(CK), 
        .Q(g5153), .QN(n1987) );
  sdffs1 \DFF_559/Q_reg  ( .DIN(g6862), .SDIN(n2593), .SSEL(test_se), .CLK(CK), 
        .Q(n2594), .QN(n1411) );
  sdffs1 \DFF_558/Q_reg  ( .DIN(g7522), .SDIN(n2085), .SSEL(test_se), .CLK(CK), 
        .Q(n2593), .QN(n1461) );
  sdffs1 \DFF_557/Q_reg  ( .DIN(g7309), .SDIN(g2673), .SSEL(test_se), .CLK(CK), 
        .Q(n2085) );
  sdffs1 \DFF_556/Q_reg  ( .DIN(g1894), .SDIN(g3846), .SSEL(test_se), .CLK(CK), 
        .Q(g2673) );
  sdffs1 \DFF_555/Q_reg  ( .DIN(g6383), .SDIN(n2151), .SSEL(test_se), .CLK(CK), 
        .Q(g3846), .QN(n2266) );
  sdffs1 \DFF_554/Q_reg  ( .DIN(n793), .SDIN(g999), .SSEL(test_se), .CLK(CK), 
        .Q(n2151) );
  sdffs1 \DFF_553/Q_reg  ( .DIN(g8865), .SDIN(g2844), .SSEL(test_se), .CLK(CK), 
        .Q(g999) );
  sdffs1 \DFF_550/Q_reg  ( .DIN(g1206), .SDIN(n2592), .SSEL(test_se), .CLK(CK), 
        .Q(g2844), .QN(\DFF_550/net775 ) );
  sdffs1 \DFF_549/Q_reg  ( .DIN(g6364), .SDIN(g205), .SSEL(test_se), .CLK(CK), 
        .Q(n2592), .QN(n2194) );
  sdffs1 \DFF_548/Q_reg  ( .DIN(g1202), .SDIN(g236), .SSEL(test_se), .CLK(CK), 
        .Q(g205) );
  sdffs1 \DFF_547/Q_reg  ( .DIN(g4649), .SDIN(n2591), .SSEL(test_se), .CLK(CK), 
        .Q(g236) );
  sdffs1 \DFF_546/Q_reg  ( .DIN(g6311), .SDIN(g8216), .SSEL(test_se), .CLK(CK), 
        .Q(n2591), .QN(n2247) );
  sdffs1 \DFF_545/Q_reg  ( .DIN(n700), .SDIN(n2590), .SSEL(test_se), .CLK(CK), 
        .Q(g8216), .QN(n1419) );
  sdffs1 \DFF_544/Q_reg  ( .DIN(n772), .SDIN(g395), .SSEL(test_se), .CLK(CK), 
        .Q(n2590), .QN(n2147) );
  sdffs1 \DFF_543/Q_reg  ( .DIN(g4646), .SDIN(n2589), .SSEL(test_se), .CLK(CK), 
        .Q(g395) );
  sdffs1 \DFF_542/Q_reg  ( .DIN(g4665), .SDIN(n2588), .SSEL(test_se), .CLK(CK), 
        .Q(n2589), .QN(n1398) );
  sdffs1 \DFF_541/Q_reg  ( .DIN(g9102), .SDIN(g4646), .SSEL(test_se), .CLK(CK), 
        .Q(n2588), .QN(n2018) );
  sdffs1 \DFF_540/Q_reg  ( .DIN(g6379), .SDIN(g1159), .SSEL(test_se), .CLK(CK), 
        .Q(g4646), .QN(n1492) );
  sdffs1 \DFF_539/Q_reg  ( .DIN(g1157), .SDIN(n2587), .SSEL(test_se), .CLK(CK), 
        .Q(g1159) );
  sdffs1 \DFF_538/Q_reg  ( .DIN(g3863), .SDIN(n2586), .SSEL(test_se), .CLK(CK), 
        .Q(n2587), .QN(n2171) );
  sdffs1 \DFF_537/Q_reg  ( .DIN(g8218), .SDIN(g1391), .SSEL(test_se), .CLK(CK), 
        .Q(n2586), .QN(n2002) );
  sdffs1 \DFF_536/Q_reg  ( .DIN(g1390), .SDIN(g1191), .SSEL(test_se), .CLK(CK), 
        .Q(g1391) );
  sdffs1 \DFF_535/Q_reg  ( .DIN(g6292), .SDIN(n2161), .SSEL(test_se), .CLK(CK), 
        .Q(g1191) );
  sdffs1 \DFF_534/Q_reg  ( .DIN(g7528), .SDIN(g1403), .SSEL(test_se), .CLK(CK), 
        .Q(n2161) );
  sdffs1 \DFF_533/Q_reg  ( .DIN(g1402), .SDIN(n2585), .SSEL(test_se), .CLK(CK), 
        .Q(g1403) );
  sdffs1 \DFF_532/Q_reg  ( .DIN(g7775), .SDIN(g1200), .SSEL(test_se), .CLK(CK), 
        .Q(n2585), .QN(n2059) );
  sdffs1 \DFF_531/Q_reg  ( .DIN(g1199), .SDIN(n2584), .SSEL(test_se), .CLK(CK), 
        .Q(g1200) );
  sdffs1 \DFF_530/Q_reg  ( .DIN(g6337), .SDIN(g3860), .SSEL(test_se), .CLK(CK), 
        .Q(n2584), .QN(n2221) );
  sdffs1 \DFF_529/Q_reg  ( .DIN(g4669), .SDIN(n2583), .SSEL(test_se), .CLK(CK), 
        .Q(g3860) );
  sdffs1 \DFF_528/Q_reg  ( .DIN(n1386), .SDIN(n2582), .SSEL(test_se), .CLK(CK), 
        .Q(n2583), .QN(n2153) );
  sdffs1 \DFF_527/Q_reg  ( .DIN(g6885), .SDIN(n2581), .SSEL(test_se), .CLK(CK), 
        .Q(n2582), .QN(\DFF_527/net752 ) );
  sdffs1 \DFF_526/Q_reg  ( .DIN(g9035), .SDIN(n2580), .SSEL(test_se), .CLK(CK), 
        .Q(n2581), .QN(n2036) );
  sdffs1 \DFF_525/Q_reg  ( .DIN(g7107), .SDIN(g3844), .SSEL(test_se), .CLK(CK), 
        .Q(n2580), .QN(n2100) );
  sdffs1 \DFF_524/Q_reg  ( .DIN(g7112), .SDIN(n2579), .SSEL(test_se), .CLK(CK), 
        .Q(g3844), .QN(n2265) );
  sdffs1 \DFF_523/Q_reg  ( .DIN(g7305), .SDIN(g201), .SSEL(test_se), .CLK(CK), 
        .Q(n2579), .QN(n2087) );
  sdffs1 \DFF_522/Q_reg  ( .DIN(g200), .SDIN(n2578), .SSEL(test_se), .CLK(CK), 
        .Q(g201) );
  sdffs1 \DFF_521/Q_reg  ( .DIN(g6876), .SDIN(g7424), .SSEL(test_se), .CLK(CK), 
        .Q(n2578), .QN(\DFF_521/net746 ) );
  sdffs1 \DFF_520/Q_reg  ( .DIN(g7425), .SDIN(n2577), .SSEL(test_se), .CLK(CK), 
        .Q(g7424) );
  sdffs1 \DFF_519/Q_reg  ( .DIN(g5165), .SDIN(n2576), .SSEL(test_se), .CLK(CK), 
        .Q(n2577), .QN(n2102) );
  sdffs1 \DFF_518/Q_reg  ( .DIN(g6884), .SDIN(g4373), .SSEL(test_se), .CLK(CK), 
        .Q(n2576), .QN(\DFF_518/net743 ) );
  sdffs1 \DFF_517/Q_reg  ( .DIN(g4372), .SDIN(g1871), .SSEL(test_se), .CLK(CK), 
        .Q(g4373), .QN(\DFF_517/net742 ) );
  sdffs1 \DFF_516/Q_reg  ( .DIN(n666), .SDIN(g4650), .SSEL(test_se), .CLK(CK), 
        .Q(g1871) );
  sdffs1 \DFF_515/Q_reg  ( .DIN(g5174), .SDIN(n2575), .SSEL(test_se), .CLK(CK), 
        .Q(g4650), .QN(n1494) );
  sdffs1 \DFF_514/Q_reg  ( .DIN(n2119), .SDIN(n2574), .SSEL(test_se), .CLK(CK), 
        .Q(n2575), .QN(n2054) );
  sdffs1 \DFF_513/Q_reg  ( .DIN(g7113), .SDIN(g595), .SSEL(test_se), .CLK(CK), 
        .Q(n2574), .QN(n2099) );
  sdffs1 \DFF_512/Q_reg  ( .DIN(g2844), .SDIN(g1911), .SSEL(test_se), .CLK(CK), 
        .Q(g595) );
  sdffs1 \DFF_511/Q_reg  ( .DIN(g6304), .SDIN(n2573), .SSEL(test_se), .CLK(CK), 
        .Q(g1911), .QN(n2057) );
  sdffs1 \DFF_510/Q_reg  ( .DIN(g5160), .SDIN(g125), .SSEL(test_se), .CLK(CK), 
        .Q(n2573), .QN(n1993) );
  sdffs1 \DFF_509/Q_reg  ( .DIN(g5155), .SDIN(n2572), .SSEL(test_se), .CLK(CK), 
        .Q(g125) );
  sdffs1 \DFF_508/Q_reg  ( .DIN(g6326), .SDIN(n2571), .SSEL(test_se), .CLK(CK), 
        .Q(n2572), .QN(n2232) );
  sdffs1 \DFF_507/Q_reg  ( .DIN(g6322), .SDIN(n2570), .SSEL(test_se), .CLK(CK), 
        .Q(n2571), .QN(n2236) );
  sdffs1 \DFF_506/Q_reg  ( .DIN(g9030), .SDIN(n2569), .SSEL(test_se), .CLK(CK), 
        .Q(n2570), .QN(n2041) );
  sdffs1 \DFF_505/Q_reg  ( .DIN(n687), .SDIN(g394), .SSEL(test_se), .CLK(CK), 
        .Q(n2569), .QN(n2138) );
  sdffs1 \DFF_504/Q_reg  ( .DIN(n769), .SDIN(g210), .SSEL(test_se), .CLK(CK), 
        .Q(g394) );
  sdffs1 \DFF_503/Q_reg  ( .DIN(g1206), .SDIN(g1398), .SSEL(test_se), .CLK(CK), 
        .Q(g210) );
  sdffs1 \DFF_502/Q_reg  ( .DIN(g1396), .SDIN(n2568), .SSEL(test_se), .CLK(CK), 
        .Q(g1398) );
  sdffs1 \DFF_501/Q_reg  ( .DIN(g7525), .SDIN(n2567), .SSEL(test_se), .CLK(CK), 
        .Q(n2568), .QN(n1462) );
  sdffs1 \DFF_500/Q_reg  ( .DIN(g6289), .SDIN(g476), .SSEL(test_se), .CLK(CK), 
        .Q(n2567), .QN(n1991) );
  sdffs1 \DFF_499/Q_reg  ( .DIN(g4646), .SDIN(n2566), .SSEL(test_se), .CLK(CK), 
        .Q(g476) );
  sdffs1 \DFF_498/Q_reg  ( .DIN(g6349), .SDIN(g5160), .SSEL(test_se), .CLK(CK), 
        .Q(n2566), .QN(n2209) );
  sdffs1 \DFF_497/Q_reg  ( .DIN(g5732), .SDIN(g146), .SSEL(test_se), .CLK(CK), 
        .Q(g5160) );
  sdffs1 \DFF_496/Q_reg  ( .DIN(g146), .SDIN(n2565), .SSEL(test_se), .CLK(CK), 
        .Q(g146), .QN(n2079) );
  sdffs1 \DFF_495/Q_reg  ( .DIN(g6841), .SDIN(n2564), .SSEL(test_se), .CLK(CK), 
        .Q(n2565), .QN(n2155) );
  sdffs1 \DFF_494/Q_reg  ( .DIN(g5167), .SDIN(n2563), .SSEL(test_se), .CLK(CK), 
        .Q(n2564), .QN(n2288) );
  sdffs1 \DFF_493/Q_reg  ( .DIN(g6345), .SDIN(n2562), .SSEL(test_se), .CLK(CK), 
        .Q(n2563), .QN(n2213) );
  sdffs1 \DFF_492/Q_reg  ( .DIN(g2663), .SDIN(g950), .SSEL(test_se), .CLK(CK), 
        .Q(n2562), .QN(n1504) );
  sdffs1 \DFF_491/Q_reg  ( .DIN(g8666), .SDIN(g1401), .SSEL(test_se), .CLK(CK), 
        .Q(g950) );
  sdffs1 \DFF_490/Q_reg  ( .DIN(g1399), .SDIN(n2561), .SSEL(test_se), .CLK(CK), 
        .Q(g1401) );
  sdffs1 \DFF_489/Q_reg  ( .DIN(g5161), .SDIN(n2560), .SSEL(test_se), .CLK(CK), 
        .Q(n2561), .QN(n1999) );
  sdffs1 \DFF_488/Q_reg  ( .DIN(n2304), .SDIN(g1312), .SSEL(test_se), .CLK(CK), 
        .Q(n2560), .QN(n2124) );
  sdffs1 \DFF_487/Q_reg  ( .DIN(g1311), .SDIN(g2663), .SSEL(test_se), .CLK(CK), 
        .Q(g1312) );
  sdffs1 \DFF_486/Q_reg  ( .DIN(g4656), .SDIN(n2559), .SSEL(test_se), .CLK(CK), 
        .Q(g2663) );
  sdffs1 \DFF_485/Q_reg  ( .DIN(g6843), .SDIN(n2558), .SSEL(test_se), .CLK(CK), 
        .Q(n2559), .QN(n2108) );
  sdffs1 \DFF_484/Q_reg  ( .DIN(g9032), .SDIN(g121), .SSEL(test_se), .CLK(CK), 
        .Q(n2558), .QN(n2038) );
  sdffs1 \DFF_483/Q_reg  ( .DIN(g5154), .SDIN(n2557), .SSEL(test_se), .CLK(CK), 
        .Q(g121) );
  sdffs1 \DFF_482/Q_reg  ( .DIN(n717), .SDIN(n2556), .SSEL(test_se), .CLK(CK), 
        .Q(n2557), .QN(n1457) );
  sdffs1 \DFF_481/Q_reg  ( .DIN(g6358), .SDIN(n2555), .SSEL(test_se), .CLK(CK), 
        .Q(n2556), .QN(n2200) );
  sdffs1 \DFF_480/Q_reg  ( .DIN(g7768), .SDIN(g1154), .SSEL(test_se), .CLK(CK), 
        .Q(n2555), .QN(n1430) );
  sdffs1 \DFF_479/Q_reg  ( .DIN(g1153), .SDIN(g543), .SSEL(test_se), .CLK(CK), 
        .Q(g1154) );
  sdffs1 \DFF_478/Q_reg  ( .DIN(g3846), .SDIN(n2554), .SSEL(test_se), .CLK(CK), 
        .Q(g543) );
  sdffs1 \DFF_477/Q_reg  ( .DIN(g1185), .SDIN(n2553), .SSEL(test_se), .CLK(CK), 
        .Q(n2554), .QN(n1402) );
  sdffs1 \DFF_476/Q_reg  ( .DIN(g7769), .SDIN(g1944), .SSEL(test_se), .CLK(CK), 
        .Q(n2553), .QN(n2066) );
  sdffs1 \DFF_475/Q_reg  ( .DIN(g6852), .SDIN(n2552), .SSEL(test_se), .CLK(CK), 
        .Q(g1944), .QN(n1445) );
  sdffs1 \DFF_474/Q_reg  ( .DIN(n793), .SDIN(n2551), .SSEL(test_se), .CLK(CK), 
        .Q(n2552), .QN(n2140) );
  sdffs1 \DFF_473/Q_reg  ( .DIN(g7119), .SDIN(n2550), .SSEL(test_se), .CLK(CK), 
        .Q(n2551), .QN(n1410) );
  sdffs1 \DFF_472/Q_reg  ( .DIN(g8874), .SDIN(g734), .SSEL(test_se), .CLK(CK), 
        .Q(n2550), .QN(n2072) );
  sdffs1 \DFF_471/Q_reg  ( .DIN(g734), .SDIN(g714), .SSEL(test_se), .CLK(CK), 
        .Q(g734), .QN(n2184) );
  sdffs1 \DFF_470/Q_reg  ( .DIN(g714), .SDIN(g1266), .SSEL(test_se), .CLK(CK), 
        .Q(g714), .QN(n2185) );
  sdffs1 \DFF_469/Q_reg  ( .DIN(g5739), .SDIN(g274), .SSEL(test_se), .CLK(CK), 
        .Q(g1266) );
  sdffs1 \DFF_468/Q_reg  ( .DIN(g4651), .SDIN(g373), .SSEL(test_se), .CLK(CK), 
        .Q(g274) );
  sdffs1 \DFF_467/Q_reg  ( .DIN(n726), .SDIN(g1395), .SSEL(test_se), .CLK(CK), 
        .Q(g373) );
  sdffs1 \DFF_466/Q_reg  ( .DIN(g1393), .SDIN(g1195), .SSEL(test_se), .CLK(CK), 
        .Q(g1395) );
  sdffs1 \DFF_465/Q_reg  ( .DIN(g6293), .SDIN(n2549), .SSEL(test_se), .CLK(CK), 
        .Q(g1195) );
  sdffs1 \DFF_464/Q_reg  ( .DIN(g9091), .SDIN(g1033), .SSEL(test_se), .CLK(CK), 
        .Q(n2549), .QN(n2029) );
  sdffs1 \DFF_463/Q_reg  ( .DIN(g9034), .SDIN(g4639), .SSEL(test_se), .CLK(CK), 
        .Q(g1033) );
  sdffs1 \DFF_462/Q_reg  ( .DIN(g7300), .SDIN(n2548), .SSEL(test_se), .CLK(CK), 
        .Q(g4639), .QN(n1480) );
  sdffs1 \DFF_461/Q_reg  ( .DIN(g7116), .SDIN(n2547), .SSEL(test_se), .CLK(CK), 
        .Q(n2548), .QN(n2096) );
  sdffs1 \DFF_460/Q_reg  ( .DIN(g6360), .SDIN(g4641), .SSEL(test_se), .CLK(CK), 
        .Q(n2547), .QN(n2198) );
  sdffs1 \DFF_459/Q_reg  ( .DIN(g7109), .SDIN(n2546), .SSEL(test_se), .CLK(CK), 
        .Q(g4641), .QN(n1506) );
  sdffs1 \DFF_458/Q_reg  ( .DIN(g8225), .SDIN(n2545), .SSEL(test_se), .CLK(CK), 
        .Q(n2546), .QN(n2073) );
  sdffs1 \DFF_457/Q_reg  ( .DIN(g9117), .SDIN(g5155), .SSEL(test_se), .CLK(CK), 
        .Q(n2545), .QN(n1440) );
  sdffs1 \DFF_456/Q_reg  ( .DIN(n793), .SDIN(n2544), .SSEL(test_se), .CLK(CK), 
        .Q(g5155), .QN(n1992) );
  sdffs1 \DFF_455/Q_reg  ( .DIN(n767), .SDIN(n2543), .SSEL(test_se), .CLK(CK), 
        .Q(n2544), .QN(n2120) );
  sdffs1 \DFF_454/Q_reg  ( .DIN(g6864), .SDIN(n2542), .SSEL(test_se), .CLK(CK), 
        .Q(n2543), .QN(n1420) );
  sdffs1 \DFF_453/Q_reg  ( .DIN(g5177), .SDIN(n2541), .SSEL(test_se), .CLK(CK), 
        .Q(n2542), .QN(n2258) );
  sdffs1 \DFF_452/Q_reg  ( .DIN(g1798), .SDIN(n2091), .SSEL(test_se), .CLK(CK), 
        .Q(n2541), .QN(n2254) );
  sdffs1 \DFF_451/Q_reg  ( .DIN(g7511), .SDIN(n2540), .SSEL(test_se), .CLK(CK), 
        .Q(n2091) );
  sdffs1 \DFF_450/Q_reg  ( .DIN(g9107), .SDIN(g5157), .SSEL(test_se), .CLK(CK), 
        .Q(n2540), .QN(n2013) );
  sdffs1 \DFF_449/Q_reg  ( .DIN(g99), .SDIN(n2539), .SSEL(test_se), .CLK(CK), 
        .Q(g5157), .QN(n1994) );
  sdffs1 \DFF_448/Q_reg  ( .DIN(g7521), .SDIN(n2538), .SSEL(test_se), .CLK(CK), 
        .Q(n2539), .QN(n2075) );
  sdffs1 \DFF_447/Q_reg  ( .DIN(g5170), .SDIN(n2537), .SSEL(test_se), .CLK(CK), 
        .Q(n2538), .QN(n2279) );
  sdffs1 \DFF_446/Q_reg  ( .DIN(n854), .SDIN(g478), .SSEL(test_se), .CLK(CK), 
        .Q(n2537), .QN(n2123) );
  sdffs1 \DFF_445/Q_reg  ( .DIN(g4648), .SDIN(n2293), .SSEL(test_se), .CLK(CK), 
        .Q(g478) );
  sdffs1 \DFF_444/Q_reg  ( .DIN(g5168), .SDIN(g1804), .SSEL(test_se), .CLK(CK), 
        .Q(n2293) );
  sdffs1 \DFF_443/Q_reg  ( .DIN(g1810), .SDIN(n2301), .SSEL(test_se), .CLK(CK), 
        .Q(g1804), .QN(n1383) );
  sdffs1 \DFF_442/Q_reg  ( .DIN(n2301), .SDIN(n2536), .SSEL(test_se), .CLK(CK), 
        .Q(n2301) );
  sdffs1 \DFF_441/Q_reg  ( .DIN(g6320), .SDIN(g4651), .SSEL(test_se), .CLK(CK), 
        .Q(n2536), .QN(n2238) );
  sdffs1 \DFF_440/Q_reg  ( .DIN(g5173), .SDIN(n2535), .SSEL(test_se), .CLK(CK), 
        .Q(g4651), .QN(n1513) );
  sdffs1 \DFF_439/Q_reg  ( .DIN(n1385), .SDIN(n2534), .SSEL(test_se), .CLK(CK), 
        .Q(n2535), .QN(n2157) );
  sdffs1 \DFF_438/Q_reg  ( .DIN(n2304), .SDIN(g108), .SSEL(test_se), .CLK(CK), 
        .Q(n2534), .QN(n2114) );
  sdffs1 \DFF_437/Q_reg  ( .DIN(g5147), .SDIN(n2533), .SSEL(test_se), .CLK(CK), 
        .Q(g108) );
  sdffs1 \DFF_436/Q_reg  ( .DIN(g9026), .SDIN(n2532), .SSEL(test_se), .CLK(CK), 
        .Q(n2533), .QN(n2045) );
  sdffs1 \DFF_435/Q_reg  ( .DIN(g9114), .SDIN(g1246), .SSEL(test_se), .CLK(CK), 
        .Q(n2532), .QN(n2006) );
  sdffs1 \DFF_434/Q_reg  ( .DIN(g1244), .SDIN(n2531), .SSEL(test_se), .CLK(CK), 
        .Q(g1246) );
  sdffs1 \DFF_433/Q_reg  ( .DIN(g6342), .SDIN(n2530), .SSEL(test_se), .CLK(CK), 
        .Q(n2531), .QN(n2216) );
  sdffs1 \DFF_432/Q_reg  ( .DIN(g9033), .SDIN(g785), .SSEL(test_se), .CLK(CK), 
        .Q(n2530), .QN(n2037) );
  sdffs1 \DFF_431/Q_reg  ( .DIN(g7100), .SDIN(n2529), .SSEL(test_se), .CLK(CK), 
        .Q(g785), .QN(n1405) );
  sdffs1 \DFF_430/Q_reg  ( .DIN(g6843), .SDIN(g1399), .SSEL(test_se), .CLK(CK), 
        .Q(n2529), .QN(n2137) );
  sdffs1 \DFF_429/Q_reg  ( .DIN(g7731), .SDIN(g1199), .SSEL(test_se), .CLK(CK), 
        .Q(g1399) );
  sdffs1 \DFF_428/Q_reg  ( .DIN(g6294), .SDIN(g233), .SSEL(test_se), .CLK(CK), 
        .Q(g1199) );
  sdffs1 \DFF_427/Q_reg  ( .DIN(n703), .SDIN(g213), .SSEL(test_se), .CLK(CK), 
        .Q(g233) );
  sdffs1 \DFF_426/Q_reg  ( .DIN(g4641), .SDIN(n2528), .SSEL(test_se), .CLK(CK), 
        .Q(g213) );
  sdffs1 \DFF_425/Q_reg  ( .DIN(n687), .SDIN(n2527), .SSEL(test_se), .CLK(CK), 
        .Q(n2528), .QN(n2121) );
  sdffs1 \DFF_424/Q_reg  ( .DIN(n2304), .SDIN(g377), .SSEL(test_se), .CLK(CK), 
        .Q(n2527), .QN(n2110) );
  sdffs1 \DFF_423/Q_reg  ( .DIN(g4643), .SDIN(n2526), .SSEL(test_se), .CLK(CK), 
        .Q(g377) );
  sdffs1 \DFF_422/Q_reg  ( .DIN(g6891), .SDIN(n2525), .SSEL(test_se), .CLK(CK), 
        .Q(n2526), .QN(\DFF_422/net647 ) );
  sdffs1 \DFF_421/Q_reg  ( .DIN(g9101), .SDIN(n2524), .SSEL(test_se), .CLK(CK), 
        .Q(n2525), .QN(n2019) );
  sdffs1 \DFF_420/Q_reg  ( .DIN(g9134), .SDIN(n2094), .SSEL(test_se), .CLK(CK), 
        .Q(n2524), .QN(n1470) );
  sdffs1 \DFF_419/Q_reg  ( .DIN(g7118), .SDIN(g4267), .SSEL(test_se), .CLK(CK), 
        .Q(n2094) );
  sdffs1 \DFF_418/Q_reg  ( .DIN(g9145), .SDIN(g4644), .SSEL(test_se), .CLK(CK), 
        .Q(g4267), .QN(n1396) );
  sdffs1 \DFF_417/Q_reg  ( .DIN(g6858), .SDIN(g1270), .SSEL(test_se), .CLK(CK), 
        .Q(g4644), .QN(n1482) );
  sdffs1 \DFF_416/Q_reg  ( .DIN(g1271), .SDIN(g1824), .SSEL(test_se), .CLK(CK), 
        .Q(g1270) );
  sdffs1 \DFF_415/Q_reg  ( .DIN(g1829), .SDIN(n2523), .SSEL(test_se), .CLK(CK), 
        .Q(g1824), .QN(n1394) );
  sdffs1 \DFF_414/Q_reg  ( .DIN(g5744), .SDIN(g1005), .SSEL(test_se), .CLK(CK), 
        .Q(n2523), .QN(n2294) );
  sdffs1 \DFF_413/Q_reg  ( .DIN(g1004), .SDIN(n2522), .SSEL(test_se), .CLK(CK), 
        .Q(g1005) );
  sdffs1 \DFF_412/Q_reg  ( .DIN(g6890), .SDIN(n2521), .SSEL(test_se), .CLK(CK), 
        .Q(n2522), .QN(\DFF_412/net637 ) );
  sdffs1 \DFF_411/Q_reg  ( .DIN(g5172), .SDIN(g953), .SSEL(test_se), .CLK(CK), 
        .Q(n2521), .QN(n2135) );
  sdffs1 \DFF_410/Q_reg  ( .DIN(g8669), .SDIN(n2520), .SSEL(test_se), .CLK(CK), 
        .Q(g953) );
  sdffs1 \DFF_409/Q_reg  ( .DIN(g6335), .SDIN(n2519), .SSEL(test_se), .CLK(CK), 
        .Q(n2520), .QN(n2223) );
  sdffs1 \DFF_408/Q_reg  ( .DIN(g2661), .SDIN(n2518), .SSEL(test_se), .CLK(CK), 
        .Q(n2519), .QN(g4667) );
  sdffs1 \DFF_407/Q_reg  ( .DIN(g2673), .SDIN(g195), .SSEL(test_se), .CLK(CK), 
        .Q(n2518), .QN(n2274) );
  sdffs1 \DFF_406/Q_reg  ( .DIN(g1194), .SDIN(g944), .SSEL(test_se), .CLK(CK), 
        .Q(g195) );
  sdffs1 \DFF_405/Q_reg  ( .DIN(g6372), .SDIN(g5146), .SSEL(test_se), .CLK(CK), 
        .Q(g944) );
  sdffs1 \DFF_404/Q_reg  ( .DIN(g94), .SDIN(n2517), .SSEL(test_se), .CLK(CK), 
        .Q(g5146), .QN(\DFF_404/net629 ) );
  sdffs1 \DFF_403/Q_reg  ( .DIN(g6359), .SDIN(n2516), .SSEL(test_se), .CLK(CK), 
        .Q(n2517), .QN(n2199) );
  sdffs1 \DFF_402/Q_reg  ( .DIN(g6296), .SDIN(n2515), .SSEL(test_se), .CLK(CK), 
        .Q(n2516), .QN(\DFF_402/net627 ) );
  sdffs1 \DFF_401/Q_reg  ( .DIN(g7762), .SDIN(g1192), .SSEL(test_se), .CLK(CK), 
        .Q(n2515), .QN(n2082) );
  sdffs1 \DFF_400/Q_reg  ( .DIN(g1191), .SDIN(n2514), .SSEL(test_se), .CLK(CK), 
        .Q(g1192) );
  sdffs1 \DFF_399/Q_reg  ( .DIN(n1384), .SDIN(n2513), .SSEL(test_se), .CLK(CK), 
        .Q(n2514), .QN(n2117) );
  sdffs1 \DFF_398/Q_reg  ( .DIN(g1824), .SDIN(g129), .SSEL(test_se), .CLK(CK), 
        .Q(n2513), .QN(n2250) );
  sdffs1 \DFF_397/Q_reg  ( .DIN(g5156), .SDIN(g1870), .SSEL(test_se), .CLK(CK), 
        .Q(g129) );
  sdffs1 \DFF_396/Q_reg  ( .DIN(n663), .SDIN(n2512), .SSEL(test_se), .CLK(CK), 
        .Q(g1870) );
  sdffs1 \DFF_395/Q_reg  ( .DIN(g8678), .SDIN(n2046), .SSEL(test_se), .CLK(CK), 
        .Q(n2512), .QN(n2063) );
  sdffs1 \DFF_394/Q_reg  ( .DIN(n2039), .SDIN(g706), .SSEL(test_se), .CLK(CK), 
        .Q(n2046) );
  sdffs1 \DFF_393/Q_reg  ( .DIN(g706), .SDIN(n2511), .SSEL(test_se), .CLK(CK), 
        .Q(g706), .QN(n2186) );
  sdffs1 \DFF_392/Q_reg  ( .DIN(g6315), .SDIN(n2510), .SSEL(test_se), .CLK(CK), 
        .Q(n2511), .QN(n2243) );
  sdffs1 \DFF_391/Q_reg  ( .DIN(g941), .SDIN(n2509), .SSEL(test_se), .CLK(CK), 
        .Q(n2510), .QN(\DFF_391/net616 ) );
  sdffs1 \DFF_390/Q_reg  ( .DIN(g6316), .SDIN(g4640), .SSEL(test_se), .CLK(CK), 
        .Q(n2509), .QN(n2242) );
  sdffs1 \DFF_388/Q_reg  ( .DIN(g7110), .SDIN(n2508), .SSEL(test_se), .CLK(CK), 
        .Q(g4640), .QN(n1488) );
  sdffs1 \DFF_387/Q_reg  ( .DIN(n1387), .SDIN(g1724), .SSEL(test_se), .CLK(CK), 
        .Q(n2508), .QN(n2166) );
  sdffs1 \DFF_386/Q_reg  ( .DIN(g5178), .SDIN(g556), .SSEL(test_se), .CLK(CK), 
        .Q(g1724) );
  sdffs1 \DFF_385/Q_reg  ( .DIN(g3847), .SDIN(g2662), .SSEL(test_se), .CLK(CK), 
        .Q(g556) );
  sdffs1 \DFF_384/Q_reg  ( .DIN(g6381), .SDIN(g103), .SSEL(test_se), .CLK(CK), 
        .Q(g2662), .QN(n2268) );
  sdffs1 \DFF_383/Q_reg  ( .DIN(g5157), .SDIN(n2507), .SSEL(test_se), .CLK(CK), 
        .Q(g103) );
  sdffs1 \DFF_382/Q_reg  ( .DIN(n854), .SDIN(n2506), .SSEL(test_se), .CLK(CK), 
        .Q(n2507), .QN(n2115) );
  sdffs1 \DFF_381/Q_reg  ( .DIN(n1401), .SDIN(n2505), .SSEL(test_se), .CLK(CK), 
        .Q(n2506), .QN(\DFF_381/net606 ) );
  sdffs1 \DFF_380/Q_reg  ( .DIN(g9389), .SDIN(g2644), .SSEL(test_se), .CLK(CK), 
        .Q(n2505), .QN(n2071) );
  sdffs1 \DFF_379/Q_reg  ( .DIN(g1798), .SDIN(n2504), .SSEL(test_se), .CLK(CK), 
        .Q(g2644), .QN(n1423) );
  sdffs1 \DFF_378/Q_reg  ( .DIN(g7770), .SDIN(n2503), .SSEL(test_se), .CLK(CK), 
        .Q(n2504), .QN(n1455) );
  sdffs1 \DFF_377/Q_reg  ( .DIN(g6297), .SDIN(g566), .SSEL(test_se), .CLK(CK), 
        .Q(n2503), .QN(\DFF_377/net602 ) );
  sdffs1 \DFF_376/Q_reg  ( .DIN(g3848), .SDIN(n2502), .SSEL(test_se), .CLK(CK), 
        .Q(g566) );
  sdffs1 \DFF_375/Q_reg  ( .DIN(n860), .SDIN(g1829), .SSEL(test_se), .CLK(CK), 
        .Q(n2502), .QN(n2105) );
  sdffs1 \DFF_374/Q_reg  ( .DIN(g1783), .SDIN(g5571), .SSEL(test_se), .CLK(CK), 
        .Q(g1829), .QN(n1382) );
  sdffs1 \DFF_373/Q_reg  ( .DIN(g1894), .SDIN(g1402), .SSEL(test_se), .CLK(CK), 
        .Q(g5571), .QN(\DFF_373/net598 ) );
  sdffs1 \DFF_372/Q_reg  ( .DIN(g6391), .SDIN(n2501), .SSEL(test_se), .CLK(CK), 
        .Q(g1402) );
  sdffs1 \DFF_371/Q_reg  ( .DIN(g2653), .SDIN(g296), .SSEL(test_se), .CLK(CK), 
        .Q(n2501), .QN(\DFF_371/net596 ) );
  sdffs1 \DFF_370/Q_reg  ( .DIN(g4643), .SDIN(g1310), .SSEL(test_se), .CLK(CK), 
        .Q(g296) );
  sdffs1 \DFF_369/Q_reg  ( .DIN(g1309), .SDIN(n2500), .SSEL(test_se), .CLK(CK), 
        .Q(g1310) );
  sdffs1 \DFF_368/Q_reg  ( .DIN(g7299), .SDIN(g4649), .SSEL(test_se), .CLK(CK), 
        .Q(n2500), .QN(n2088) );
  sdffs1 \DFF_367/Q_reg  ( .DIN(g5736), .SDIN(g855), .SSEL(test_se), .CLK(CK), 
        .Q(g4649), .QN(n1484) );
  sdffs1 \DFF_366/Q_reg  ( .DIN(g855), .SDIN(g3130), .SSEL(test_se), .CLK(CK), 
        .Q(g855), .QN(n1471) );
  sdffs1 \DFF_365/Q_reg  ( .DIN(g1198), .SDIN(g3855), .SSEL(test_se), .CLK(CK), 
        .Q(g3130), .QN(\DFF_365/net590 ) );
  sdffs1 \DFF_364/Q_reg  ( .DIN(g4316), .SDIN(g477), .SSEL(test_se), .CLK(CK), 
        .Q(g3855), .QN(n1468) );
  sdffs1 \DFF_363/Q_reg  ( .DIN(g4647), .SDIN(n2499), .SSEL(test_se), .CLK(CK), 
        .Q(g477) );
  sdffs1 \DFF_362/Q_reg  ( .DIN(g5181), .SDIN(n2498), .SSEL(test_se), .CLK(CK), 
        .Q(n2499), .QN(n1458) );
  sdffs1 \DFF_361/Q_reg  ( .DIN(n843), .SDIN(g1244), .SSEL(test_se), .CLK(CK), 
        .Q(n2498), .QN(n2113) );
  sdffs1 \DFF_360/Q_reg  ( .DIN(g2659), .SDIN(g949), .SSEL(test_se), .CLK(CK), 
        .Q(g1244) );
  sdffs1 \DFF_359/Q_reg  ( .DIN(g8665), .SDIN(n2497), .SSEL(test_se), .CLK(CK), 
        .Q(g949) );
  sdffs1 \DFF_358/Q_reg  ( .DIN(g9087), .SDIN(n2496), .SSEL(test_se), .CLK(CK), 
        .Q(n2497), .QN(n2033) );
  sdffs1 \DFF_357/Q_reg  ( .DIN(g9027), .SDIN(g7729), .SSEL(test_se), .CLK(CK), 
        .Q(n2496), .QN(n2044) );
  sdffs1 \DFF_356/Q_reg  ( .DIN(g7729), .SDIN(n2495), .SSEL(test_se), .CLK(CK), 
        .Q(g7729), .QN(n1990) );
  sdffs1 \DFF_354/Q_reg  ( .DIN(g7099), .SDIN(g6841), .SSEL(test_se), .CLK(CK), 
        .Q(n2495), .QN(n1432) );
  sdffs1 \DFF_353/Q_reg  ( .DIN(g9376), .SDIN(n2494), .SSEL(test_se), .CLK(CK), 
        .Q(g6841), .QN(n1511) );
  sdffs1 \DFF_352/Q_reg  ( .DIN(n854), .SDIN(n2493), .SSEL(test_se), .CLK(CK), 
        .Q(n2494), .QN(n2159) );
  sdffs1 \DFF_351/Q_reg  ( .DIN(g9098), .SDIN(g456), .SSEL(test_se), .CLK(CK), 
        .Q(n2493), .QN(n2022) );
  sdffs1 \DFF_350/Q_reg  ( .DIN(g4641), .SDIN(n2492), .SSEL(test_se), .CLK(CK), 
        .Q(g456) );
  sdffs1 \DFF_349/Q_reg  ( .DIN(g5166), .SDIN(n2491), .SSEL(test_se), .CLK(CK), 
        .Q(n2492), .QN(n2287) );
  sdffs1 \DFF_348/Q_reg  ( .DIN(g9095), .SDIN(g316), .SSEL(test_se), .CLK(CK), 
        .Q(n2491), .QN(n2025) );
  sdffs1 \DFF_347/Q_reg  ( .DIN(n827), .SDIN(n2490), .SSEL(test_se), .CLK(CK), 
        .Q(g316) );
  sdffs1 \DFF_346/Q_reg  ( .DIN(n854), .SDIN(n2489), .SSEL(test_se), .CLK(CK), 
        .Q(n2490), .QN(n2109) );
  sdffs1 \DFF_345/Q_reg  ( .DIN(g7114), .SDIN(g4645), .SSEL(test_se), .CLK(CK), 
        .Q(n2489), .QN(n2098) );
  sdffs1 \DFF_344/Q_reg  ( .DIN(g6857), .SDIN(n2488), .SSEL(test_se), .CLK(CK), 
        .Q(g4645), .QN(n1508) );
  sdffs1 \DFF_343/Q_reg  ( .DIN(g6370), .SDIN(g3096), .SSEL(test_se), .CLK(CK), 
        .Q(n2488), .QN(n2188) );
  sdffs1 \DFF_342/Q_reg  ( .DIN(g1194), .SDIN(n1385), .SSEL(test_se), .CLK(CK), 
        .Q(g3096), .QN(\DFF_342/net567 ) );
  sdffs1 \DFF_341/Q_reg  ( .DIN(n2296), .SDIN(g93), .SSEL(test_se), .CLK(CK), 
        .Q(n1385), .QN(n1414) );
  sdffs1 \DFF_340/Q_reg  ( .DIN(g5145), .SDIN(g1404), .SSEL(test_se), .CLK(CK), 
        .Q(g93) );
  sdffs1 \DFF_339/Q_reg  ( .DIN(g1403), .SDIN(g1004), .SSEL(test_se), .CLK(CK), 
        .Q(g1404) );
  sdffs1 \DFF_338/Q_reg  ( .DIN(n673), .SDIN(g890), .SSEL(test_se), .CLK(CK), 
        .Q(g1004) );
  sdffs1 \DFF_337/Q_reg  ( .DIN(g7102), .SDIN(g3845), .SSEL(test_se), .CLK(CK), 
        .Q(g890) );
  sdffs1 \DFF_336/Q_reg  ( .DIN(g6384), .SDIN(n2487), .SSEL(test_se), .CLK(CK), 
        .Q(g3845), .QN(n1449) );
  sdffs1 \DFF_335/Q_reg  ( .DIN(n1386), .SDIN(n2486), .SSEL(test_se), .CLK(CK), 
        .Q(n2487), .QN(n2141) );
  sdffs1 \DFF_334/Q_reg  ( .DIN(g5182), .SDIN(g2888), .SSEL(test_se), .CLK(CK), 
        .Q(n2486), .QN(n2273) );
  sdffs1 \DFF_333/Q_reg  ( .DIN(g7106), .SDIN(g290), .SSEL(test_se), .CLK(CK), 
        .Q(g2888), .QN(n2131) );
  sdffs1 \DFF_332/Q_reg  ( .DIN(g3096), .SDIN(g3850), .SSEL(test_se), .CLK(CK), 
        .Q(g290) );
  sdffs1 \DFF_331/Q_reg  ( .DIN(g7302), .SDIN(g199), .SSEL(test_se), .CLK(CK), 
        .Q(g3850), .QN(n2264) );
  sdffs1 \DFF_330/Q_reg  ( .DIN(n1418), .SDIN(n2485), .SSEL(test_se), .CLK(CK), 
        .Q(g199) );
  sdffs1 \DFF_329/Q_reg  ( .DIN(n2300), .SDIN(g2653), .SSEL(test_se), .CLK(CK), 
        .Q(n2485), .QN(n2248) );
  sdffs1 \DFF_328/Q_reg  ( .DIN(g7104), .SDIN(n2484), .SSEL(test_se), .CLK(CK), 
        .Q(g2653), .QN(n1475) );
  sdffs1 \DFF_327/Q_reg  ( .DIN(g6363), .SDIN(g516), .SSEL(test_se), .CLK(CK), 
        .Q(n2484), .QN(n2195) );
  sdffs1 \DFF_326/Q_reg  ( .DIN(g4650), .SDIN(n2483), .SSEL(test_se), .CLK(CK), 
        .Q(g516) );
  sdffs1 \DFF_325/Q_reg  ( .DIN(g9089), .SDIN(n2482), .SSEL(test_se), .CLK(CK), 
        .Q(n2483), .QN(n2031) );
  sdffs1 \DFF_324/Q_reg  ( .DIN(g2644), .SDIN(n2481), .SSEL(test_se), .CLK(CK), 
        .Q(n2482), .QN(n2253) );
  sdffs1 \DFF_323/Q_reg  ( .DIN(n860), .SDIN(g375), .SSEL(test_se), .CLK(CK), 
        .Q(n2481), .QN(n1397) );
  sdffs1 \DFF_322/Q_reg  ( .DIN(g4641), .SDIN(n2480), .SSEL(test_se), .CLK(CK), 
        .Q(g375) );
  sdffs1 \DFF_321/Q_reg  ( .DIN(g8675), .SDIN(g1157), .SSEL(test_se), .CLK(CK), 
        .Q(n2480), .QN(n2169) );
  sdffs1 \DFF_320/Q_reg  ( .DIN(g1156), .SDIN(n2479), .SSEL(test_se), .CLK(CK), 
        .Q(g1157) );
  sdffs1 \DFF_319/Q_reg  ( .DIN(g9090), .SDIN(n2478), .SSEL(test_se), .CLK(CK), 
        .Q(n2479), .QN(n2030) );
  sdffs1 \DFF_318/Q_reg  ( .DIN(g6333), .SDIN(n2477), .SSEL(test_se), .CLK(CK), 
        .Q(n2478), .QN(n2225) );
  sdffs1 \DFF_317/Q_reg  ( .DIN(g6321), .SDIN(n2476), .SSEL(test_se), .CLK(CK), 
        .Q(n2477), .QN(n2237) );
  sdffs1 \DFF_316/Q_reg  ( .DIN(g8873), .SDIN(n2475), .SSEL(test_se), .CLK(CK), 
        .Q(n2476), .QN(n2047) );
  sdffs1 \DFF_315/Q_reg  ( .DIN(g5183), .SDIN(n2474), .SSEL(test_se), .CLK(CK), 
        .Q(n2475), .QN(g8219) );
  sdffs1 \DFF_314/Q_reg  ( .DIN(g6877), .SDIN(g4371), .SSEL(test_se), .CLK(CK), 
        .Q(n2474), .QN(\DFF_314/net539 ) );
  sdffs1 \DFF_313/Q_reg  ( .DIN(g4267), .SDIN(g8217), .SSEL(test_se), .CLK(CK), 
        .Q(g4371), .QN(\DFF_313/net538 ) );
  sdffs1 \DFF_312/Q_reg  ( .DIN(g7111), .SDIN(n2473), .SSEL(test_se), .CLK(CK), 
        .Q(g8217) );
  sdffs1 \DFF_311/Q_reg  ( .DIN(g9097), .SDIN(g458), .SSEL(test_se), .CLK(CK), 
        .Q(n2473), .QN(n2023) );
  sdffs1 \DFF_310/Q_reg  ( .DIN(g4643), .SDIN(n2472), .SSEL(test_se), .CLK(CK), 
        .Q(g458) );
  sdffs1 \DFF_309/Q_reg  ( .DIN(g6329), .SDIN(g1156), .SSEL(test_se), .CLK(CK), 
        .Q(n2472), .QN(n2229) );
  sdffs1 \DFF_308/Q_reg  ( .DIN(g1944), .SDIN(n2471), .SSEL(test_se), .CLK(CK), 
        .Q(g1156) );
  sdffs1 \DFF_307/Q_reg  ( .DIN(n772), .SDIN(g1390), .SSEL(test_se), .CLK(CK), 
        .Q(n2471), .QN(n1391) );
  sdffs1 \DFF_306/Q_reg  ( .DIN(g8216), .SDIN(n2470), .SSEL(test_se), .CLK(CK), 
        .Q(g1390) );
  sdffs1 \DFF_304/Q_reg  ( .DIN(g9112), .SDIN(n2469), .SSEL(test_se), .CLK(CK), 
        .Q(n2470), .QN(n2008) );
  sdffs1 \DFF_303/Q_reg  ( .DIN(n843), .SDIN(n2468), .SSEL(test_se), .CLK(CK), 
        .Q(n2469), .QN(n2170) );
  sdffs1 \DFF_302/Q_reg  ( .DIN(g9028), .SDIN(g594), .SSEL(test_se), .CLK(CK), 
        .Q(n2468), .QN(n2043) );
  sdffs1 \DFF_301/Q_reg  ( .DIN(g4668), .SDIN(n2467), .SSEL(test_se), .CLK(CK), 
        .Q(g594) );
  sdffs1 \DFF_300/Q_reg  ( .DIN(n1416), .SDIN(n2466), .SSEL(test_se), .CLK(CK), 
        .Q(n2467), .QN(n1416) );
  sdffs1 \DFF_299/Q_reg  ( .DIN(g6353), .SDIN(n2465), .SSEL(test_se), .CLK(CK), 
        .Q(n2466), .QN(n2205) );
  sdffs1 \DFF_297/Q_reg  ( .DIN(n792), .SDIN(g371), .SSEL(test_se), .CLK(CK), 
        .Q(n2465), .QN(n1388) );
  sdffs1 \DFF_296/Q_reg  ( .DIN(g3130), .SDIN(n2464), .SSEL(test_se), .CLK(CK), 
        .Q(g371) );
  sdffs1 \DFF_295/Q_reg  ( .DIN(g6365), .SDIN(g665), .SSEL(test_se), .CLK(CK), 
        .Q(n2464), .QN(n2193) );
  sdffs1 \DFF_294/Q_reg  ( .DIN(g665), .SDIN(n2463), .SSEL(test_se), .CLK(CK), 
        .Q(g665), .QN(n2179) );
  sdffs1 \DFF_293/Q_reg  ( .DIN(g9113), .SDIN(n2462), .SSEL(test_se), .CLK(CK), 
        .Q(n2463), .QN(n2007) );
  sdffs1 \DFF_292/Q_reg  ( .DIN(g5743), .SDIN(n2461), .SSEL(test_se), .CLK(CK), 
        .Q(n2462), .QN(n2259) );
  sdffs1 \DFF_291/Q_reg  ( .DIN(g7733), .SDIN(g6843), .SSEL(test_se), .CLK(CK), 
        .Q(n2461), .QN(n2081) );
  sdffs1 \DFF_290/Q_reg  ( .DIN(g9374), .SDIN(n2460), .SSEL(test_se), .CLK(CK), 
        .Q(g6843), .QN(n1496) );
  sdffs1 \DFF_289/Q_reg  ( .DIN(g1014), .SDIN(g235), .SSEL(test_se), .CLK(CK), 
        .Q(n2460), .QN(n2052) );
  sdffs1 \DFF_288/Q_reg  ( .DIN(g4648), .SDIN(g215), .SSEL(test_se), .CLK(CK), 
        .Q(g235) );
  sdffs1 \DFF_287/Q_reg  ( .DIN(n839), .SDIN(g3191), .SSEL(test_se), .CLK(CK), 
        .Q(g215) );
  sdffs1 \DFF_286/Q_reg  ( .DIN(g1202), .SDIN(n2459), .SSEL(test_se), .CLK(CK), 
        .Q(g3191), .QN(\DFF_286/net511 ) );
  sdffs1 \DFF_285/Q_reg  ( .DIN(g9115), .SDIN(n2458), .SSEL(test_se), .CLK(CK), 
        .Q(n2459), .QN(n2005) );
  sdffs1 \DFF_284/Q_reg  ( .DIN(g9029), .SDIN(g98), .SSEL(test_se), .CLK(CK), 
        .Q(n2458), .QN(n2042) );
  sdffs1 \DFF_283/Q_reg  ( .DIN(g5146), .SDIN(g374), .SSEL(test_se), .CLK(CK), 
        .Q(g98) );
  sdffs1 \DFF_282/Q_reg  ( .DIN(g4640), .SDIN(g1147), .SSEL(test_se), .CLK(CK), 
        .Q(g374) );
  sdffs1 \DFF_281/Q_reg  ( .DIN(g1146), .SDIN(g8218), .SSEL(test_se), .CLK(CK), 
        .Q(g1147) );
  sdffs1 \DFF_280/Q_reg  ( .DIN(g8957), .SDIN(n2457), .SSEL(test_se), .CLK(CK), 
        .Q(g8218), .QN(n1401) );
  sdffs1 \DFF_279/Q_reg  ( .DIN(g6344), .SDIN(g436), .SSEL(test_se), .CLK(CK), 
        .Q(n2457), .QN(n2214) );
  sdffs1 \DFF_278/Q_reg  ( .DIN(g4651), .SDIN(n2272), .SSEL(test_se), .CLK(CK), 
        .Q(g436) );
  sdffs1 \DFF_277/Q_reg  ( .DIN(g4667), .SDIN(n2456), .SSEL(test_se), .CLK(CK), 
        .Q(n2272) );
  sdffs1 \DFF_276/Q_reg  ( .DIN(g8960), .SDIN(n2455), .SSEL(test_se), .CLK(CK), 
        .Q(n2456), .QN(n2058) );
  sdffs1 \DFF_275/Q_reg  ( .DIN(g6361), .SDIN(g1894), .SSEL(test_se), .CLK(CK), 
        .Q(n2455), .QN(n2197) );
  sdffs1 \DFF_274/Q_reg  ( .DIN(g1234), .SDIN(g859), .SSEL(test_se), .CLK(CK), 
        .Q(g1894) );
  sdffs1 \DFF_273/Q_reg  ( .DIN(g859), .SDIN(n2454), .SSEL(test_se), .CLK(CK), 
        .Q(g859), .QN(n1469) );
  sdffs1 \DFF_272/Q_reg  ( .DIN(n843), .SDIN(g150), .SSEL(test_se), .CLK(CK), 
        .Q(n2454), .QN(n2144) );
  sdffs1 \DFF_271/Q_reg  ( .DIN(g150), .SDIN(g5145), .SSEL(test_se), .CLK(CK), 
        .Q(g150), .QN(n2065) );
  sdffs1 \DFF_270/Q_reg  ( .DIN(g92), .SDIN(g1146), .SSEL(test_se), .CLK(CK), 
        .Q(g5145), .QN(\DFF_270/net495 ) );
  sdffs1 \DFF_269/Q_reg  ( .DIN(g2888), .SDIN(g293), .SSEL(test_se), .CLK(CK), 
        .Q(g1146) );
  sdffs1 \DFF_268/Q_reg  ( .DIN(g4640), .SDIN(n2453), .SSEL(test_se), .CLK(CK), 
        .Q(g293) );
  sdffs1 \DFF_267/Q_reg  ( .DIN(g7307), .SDIN(n2452), .SSEL(test_se), .CLK(CK), 
        .Q(n2453), .QN(n1473) );
  sdffs1 \DFF_266/Q_reg  ( .DIN(g1783), .SDIN(n2451), .SSEL(test_se), .CLK(CK), 
        .Q(n2452), .QN(n2252) );
  sdffs1 \DFF_265/Q_reg  ( .DIN(n2304), .SDIN(g661), .SSEL(test_se), .CLK(CK), 
        .Q(n2451), .QN(n1409) );
  sdffs1 \DFF_264/Q_reg  ( .DIN(g661), .SDIN(n2450), .SSEL(test_se), .CLK(CK), 
        .Q(g661), .QN(n2178) );
  sdffs1 \DFF_263/Q_reg  ( .DIN(n793), .SDIN(g158), .SSEL(test_se), .CLK(CK), 
        .Q(n2450), .QN(n2160) );
  sdffs1 \DFF_262/Q_reg  ( .DIN(g158), .SDIN(g4647), .SSEL(test_se), .CLK(CK), 
        .Q(g158), .QN(n1418) );
  sdffs1 \DFF_261/Q_reg  ( .DIN(g6378), .SDIN(n2449), .SSEL(test_se), .CLK(CK), 
        .Q(g4647), .QN(n1502) );
  sdffs1 \DFF_260/Q_reg  ( .DIN(g6889), .SDIN(n2448), .SSEL(test_se), .CLK(CK), 
        .Q(n2449), .QN(\DFF_260/net485 ) );
  sdffs1 \DFF_259/Q_reg  ( .DIN(g6366), .SDIN(g231), .SSEL(test_se), .CLK(CK), 
        .Q(n2448), .QN(n2192) );
  sdffs1 \DFF_258/Q_reg  ( .DIN(g4644), .SDIN(n2447), .SSEL(test_se), .CLK(CK), 
        .Q(g231) );
  sdffs1 \DFF_257/Q_reg  ( .DIN(g1829), .SDIN(g211), .SSEL(test_se), .CLK(CK), 
        .Q(n2447), .QN(n2251) );
  sdffs1 \DFF_256/Q_reg  ( .DIN(g4639), .SDIN(n2446), .SSEL(test_se), .CLK(CK), 
        .Q(g211) );
  sdffs1 \DFF_255/Q_reg  ( .DIN(g6328), .SDIN(g92), .SSEL(test_se), .CLK(CK), 
        .Q(n2446), .QN(n2230) );
  sdffs1 \DFF_254/Q_reg  ( .DIN(n854), .SDIN(n2445), .SSEL(test_se), .CLK(CK), 
        .Q(g92) );
  sdffs1 \DFF_253/Q_reg  ( .DIN(g7306), .SDIN(n2444), .SSEL(test_se), .CLK(CK), 
        .Q(n2445), .QN(n2086) );
  sdffs1 \DFF_252/Q_reg  ( .DIN(g6300), .SDIN(n2443), .SSEL(test_se), .CLK(CK), 
        .Q(n2444), .QN(\DFF_252/net477 ) );
  sdffs1 \DFF_251/Q_reg  ( .DIN(g8674), .SDIN(n2442), .SSEL(test_se), .CLK(CK), 
        .Q(n2443), .QN(n2074) );
  sdffs1 \DFF_250/Q_reg  ( .DIN(g646), .SDIN(g234), .SSEL(test_se), .CLK(CK), 
        .Q(n2442), .QN(n2175) );
  sdffs1 \DFF_249/Q_reg  ( .DIN(n805), .SDIN(g214), .SSEL(test_se), .CLK(CK), 
        .Q(g234) );
  sdffs1 \DFF_248/Q_reg  ( .DIN(n834), .SDIN(g2654), .SSEL(test_se), .CLK(CK), 
        .Q(g214) );
  sdffs1 \DFF_247/Q_reg  ( .DIN(g2654), .SDIN(n2441), .SSEL(test_se), .CLK(CK), 
        .Q(g2654), .QN(n2003) );
  sdffs1 \DFF_246/Q_reg  ( .DIN(g6334), .SDIN(g313), .SSEL(test_se), .CLK(CK), 
        .Q(n2441), .QN(n2224) );
  sdffs1 \DFF_245/Q_reg  ( .DIN(g4645), .SDIN(n2440), .SSEL(test_se), .CLK(CK), 
        .Q(g313) );
  sdffs1 \DFF_244/Q_reg  ( .DIN(g6367), .SDIN(n2439), .SSEL(test_se), .CLK(CK), 
        .Q(n2440), .QN(n2191) );
  sdffs1 \DFF_243/Q_reg  ( .DIN(g7758), .SDIN(n2438), .SSEL(test_se), .CLK(CK), 
        .Q(n2439), .QN(n2089) );
  sdffs1 \DFF_242/Q_reg  ( .DIN(g7756), .SDIN(g951), .SSEL(test_se), .CLK(CK), 
        .Q(n2438), .QN(n2093) );
  sdffs1 \DFF_241/Q_reg  ( .DIN(g8667), .SDIN(g7507), .SSEL(test_se), .CLK(CK), 
        .Q(g951) );
  sdffs1 \DFF_240/Q_reg  ( .DIN(g5184), .SDIN(g475), .SSEL(test_se), .CLK(CK), 
        .Q(g7507), .QN(n2271) );
  sdffs1 \DFF_239/Q_reg  ( .DIN(g4645), .SDIN(n2437), .SSEL(test_se), .CLK(CK), 
        .Q(g475) );
  sdffs1 \DFF_238/Q_reg  ( .DIN(g7516), .SDIN(g232), .SSEL(test_se), .CLK(CK), 
        .Q(n2437), .QN(n1464) );
  sdffs1 \DFF_237/Q_reg  ( .DIN(g4645), .SDIN(n2289), .SSEL(test_se), .CLK(CK), 
        .Q(g232) );
  sdffs1 \DFF_236/Q_reg  ( .DIN(g6874), .SDIN(g212), .SSEL(test_se), .CLK(CK), 
        .Q(n2289) );
  sdffs1 \DFF_235/Q_reg  ( .DIN(g4640), .SDIN(g145), .SSEL(test_se), .CLK(CK), 
        .Q(g212) );
  sdffs1 \DFF_234/Q_reg  ( .DIN(g5152), .SDIN(g5147), .SSEL(test_se), .CLK(CK), 
        .Q(g145) );
  sdffs1 \DFF_233/Q_reg  ( .DIN(g104), .SDIN(g954), .SSEL(test_se), .CLK(CK), 
        .Q(g5147), .QN(n1997) );
  sdffs1 \DFF_232/Q_reg  ( .DIN(g8670), .SDIN(n2436), .SSEL(test_se), .CLK(CK), 
        .Q(g954) );
  sdffs1 \DFF_231/Q_reg  ( .DIN(g6324), .SDIN(n2435), .SSEL(test_se), .CLK(CK), 
        .Q(n2436), .QN(n2234) );
  sdffs1 \DFF_230/Q_reg  ( .DIN(g7765), .SDIN(n2434), .SSEL(test_se), .CLK(CK), 
        .Q(n2435), .QN(n2070) );
  sdffs1 \DFF_229/Q_reg  ( .DIN(g1005), .SDIN(n2433), .SSEL(test_se), .CLK(CK), 
        .Q(n2434), .QN(n2050) );
  sdffs1 \DFF_228/Q_reg  ( .DIN(g6343), .SDIN(n2432), .SSEL(test_se), .CLK(CK), 
        .Q(n2433), .QN(n2215) );
  sdffs1 \DFF_226/Q_reg  ( .DIN(g5738), .SDIN(n2431), .SSEL(test_se), .CLK(CK), 
        .Q(n2432), .QN(n2172) );
  sdffs1 \DFF_225/Q_reg  ( .DIN(n687), .SDIN(n2430), .SSEL(test_se), .CLK(CK), 
        .Q(n2431), .QN(n2107) );
  sdffs1 \DFF_224/Q_reg  ( .DIN(g6368), .SDIN(n2429), .SSEL(test_se), .CLK(CK), 
        .Q(n2430), .QN(n2190) );
  sdffs1 \DFF_223/Q_reg  ( .DIN(g5737), .SDIN(g952), .SSEL(test_se), .CLK(CK), 
        .Q(n2429), .QN(n2173) );
  sdffs1 \DFF_222/Q_reg  ( .DIN(g8668), .SDIN(n2283), .SSEL(test_se), .CLK(CK), 
        .Q(g952) );
  sdffs1 \DFF_221/Q_reg  ( .DIN(g5179), .SDIN(n2428), .SSEL(test_se), .CLK(CK), 
        .Q(n2283) );
  sdffs1 \DFF_220/Q_reg  ( .DIN(g8870), .SDIN(g533), .SSEL(test_se), .CLK(CK), 
        .Q(n2428), .QN(n2049) );
  sdffs1 \DFF_219/Q_reg  ( .DIN(g3191), .SDIN(n2427), .SSEL(test_se), .CLK(CK), 
        .Q(g533) );
  sdffs1 \DFF_218/Q_reg  ( .DIN(g6298), .SDIN(n2426), .SSEL(test_se), .CLK(CK), 
        .Q(n2427), .QN(\DFF_218/net443 ) );
  sdffs1 \DFF_217/Q_reg  ( .DIN(g9116), .SDIN(g1197), .SSEL(test_se), .CLK(CK), 
        .Q(n2426), .QN(n2004) );
  sdffs1 \DFF_216/Q_reg  ( .DIN(g1196), .SDIN(n2284), .SSEL(test_se), .CLK(CK), 
        .Q(g1197) );
  sdffs1 \DFF_215/Q_reg  ( .DIN(g6887), .SDIN(n2425), .SSEL(test_se), .CLK(CK), 
        .Q(n2284) );
  sdffs1 \DFF_214/Q_reg  ( .DIN(g6354), .SDIN(n2424), .SSEL(test_se), .CLK(CK), 
        .Q(n2425), .QN(n2204) );
  sdffs1 \DFF_213/Q_reg  ( .DIN(g6357), .SDIN(g457), .SSEL(test_se), .CLK(CK), 
        .Q(n2424), .QN(n2201) );
  sdffs1 \DFF_212/Q_reg  ( .DIN(g4642), .SDIN(g317), .SSEL(test_se), .CLK(CK), 
        .Q(g457) );
  sdffs1 \DFF_211/Q_reg  ( .DIN(n761), .SDIN(n2423), .SSEL(test_se), .CLK(CK), 
        .Q(g317) );
  sdffs1 \DFF_210/Q_reg  ( .DIN(g8875), .SDIN(n2422), .SSEL(test_se), .CLK(CK), 
        .Q(n2423), .QN(n2064) );
  sdffs1 \DFF_209/Q_reg  ( .DIN(g9031), .SDIN(n2421), .SSEL(test_se), .CLK(CK), 
        .Q(n2422), .QN(n2040) );
  sdffs1 \DFF_208/Q_reg  ( .DIN(g8869), .SDIN(n2420), .SSEL(test_se), .CLK(CK), 
        .Q(n2421), .QN(n1433) );
  sdffs1 \DFF_207/Q_reg  ( .DIN(n860), .SDIN(n2419), .SSEL(test_se), .CLK(CK), 
        .Q(n2420), .QN(n2150) );
  sdffs1 \DFF_206/Q_reg  ( .DIN(g7774), .SDIN(g141), .SSEL(test_se), .CLK(CK), 
        .Q(n2419), .QN(n2055) );
  sdffs1 \DFF_205/Q_reg  ( .DIN(g5151), .SDIN(g1396), .SSEL(test_se), .CLK(CK), 
        .Q(g141) );
  sdffs1 \DFF_204/Q_reg  ( .DIN(g8217), .SDIN(g474), .SSEL(test_se), .CLK(CK), 
        .Q(g1396) );
  sdffs1 \DFF_203/Q_reg  ( .DIN(g4644), .SDIN(n2418), .SSEL(test_se), .CLK(CK), 
        .Q(g474) );
  sdffs1 \DFF_202/Q_reg  ( .DIN(g6863), .SDIN(n2417), .SSEL(test_se), .CLK(CK), 
        .Q(n2418), .QN(n1390) );
  sdffs1 \DFF_201/Q_reg  ( .DIN(g7513), .SDIN(n2416), .SSEL(test_se), .CLK(CK), 
        .Q(n2417), .QN(n2083) );
  sdffs1 \DFF_200/Q_reg  ( .DIN(g6867), .SDIN(g104), .SSEL(test_se), .CLK(CK), 
        .Q(n2416), .QN(\DFF_200/net425 ) );
  sdffs1 \DFF_199/Q_reg  ( .DIN(n843), .SDIN(g4648), .SSEL(test_se), .CLK(CK), 
        .Q(g104) );
  sdffs1 \DFF_198/Q_reg  ( .DIN(g6377), .SDIN(n2415), .SSEL(test_se), .CLK(CK), 
        .Q(g4648), .QN(n1486) );
  sdffs1 \DFF_197/Q_reg  ( .DIN(n843), .SDIN(n2414), .SSEL(test_se), .CLK(CK), 
        .Q(n2415), .QN(n2156) );
  sdffs1 \DFF_196/Q_reg  ( .DIN(n772), .SDIN(g1308), .SSEL(test_se), .CLK(CK), 
        .Q(n2414), .QN(n2103) );
  sdffs1 \DFF_195/Q_reg  ( .DIN(g6385), .SDIN(n2413), .SSEL(test_se), .CLK(CK), 
        .Q(g1308) );
  sdffs1 \DFF_194/Q_reg  ( .DIN(g7761), .SDIN(n2412), .SSEL(test_se), .CLK(CK), 
        .Q(n2413), .QN(n2084) );
  sdffs1 \DFF_193/Q_reg  ( .DIN(g9085), .SDIN(n2411), .SSEL(test_se), .CLK(CK), 
        .Q(n2412), .QN(n2035) );
  sdffs1 \DFF_192/Q_reg  ( .DIN(g6314), .SDIN(g5149), .SSEL(test_se), .CLK(CK), 
        .Q(n2411), .QN(n2244) );
  sdffs1 \DFF_191/Q_reg  ( .DIN(n2304), .SDIN(g5148), .SSEL(test_se), .CLK(CK), 
        .Q(g5149) );
  sdffs1 \DFF_190/Q_reg  ( .DIN(g109), .SDIN(g669), .SSEL(test_se), .CLK(CK), 
        .Q(g5148), .QN(n2000) );
  sdffs1 \DFF_189/Q_reg  ( .DIN(g669), .SDIN(n2410), .SSEL(test_se), .CLK(CK), 
        .Q(g669), .QN(n2180) );
  sdffs1 \DFF_188/Q_reg  ( .DIN(g6380), .SDIN(n2409), .SSEL(test_se), .CLK(CK), 
        .Q(n2410), .QN(n1403) );
  sdffs1 \DFF_187/Q_reg  ( .DIN(g4667), .SDIN(n2408), .SSEL(test_se), .CLK(CK), 
        .Q(n2409), .QN(n2275) );
  sdffs1 \DFF_186/Q_reg  ( .DIN(n767), .SDIN(n2053), .SSEL(test_se), .CLK(CK), 
        .Q(n2408), .QN(n2106) );
  sdffs1 \DFF_185/Q_reg  ( .DIN(g7518), .SDIN(g579), .SSEL(test_se), .CLK(CK), 
        .Q(n2053) );
  sdffs1 \DFF_184/Q_reg  ( .DIN(g3850), .SDIN(n2407), .SSEL(test_se), .CLK(CK), 
        .Q(g579) );
  sdffs1 \DFF_183/Q_reg  ( .DIN(g2672), .SDIN(n2406), .SSEL(test_se), .CLK(CK), 
        .Q(n2407), .QN(n2277) );
  sdffs1 \DFF_182/Q_reg  ( .DIN(g1804), .SDIN(n2405), .SSEL(test_se), .CLK(CK), 
        .Q(n2406), .QN(n2255) );
  sdffs1 \DFF_181/Q_reg  ( .DIN(g7510), .SDIN(n2404), .SSEL(test_se), .CLK(CK), 
        .Q(n2405), .QN(n2092) );
  sdffs1 \DFF_180/Q_reg  ( .DIN(g6882), .SDIN(n2403), .SSEL(test_se), .CLK(CK), 
        .Q(n2404), .QN(\DFF_180/net405 ) );
  sdffs1 \DFF_179/Q_reg  ( .DIN(g9106), .SDIN(n2402), .SSEL(test_se), .CLK(CK), 
        .Q(n2403), .QN(n2014) );
  sdffs1 \DFF_178/Q_reg  ( .DIN(g6312), .SDIN(g5152), .SSEL(test_se), .CLK(CK), 
        .Q(n2402), .QN(n2246) );
  sdffs1 \DFF_177/Q_reg  ( .DIN(n860), .SDIN(n2401), .SSEL(test_se), .CLK(CK), 
        .Q(g5152), .QN(n2001) );
  sdffs1 \DFF_176/Q_reg  ( .DIN(g9086), .SDIN(g7505), .SSEL(test_se), .CLK(CK), 
        .Q(n2401), .QN(n2034) );
  sdffs1 \DFF_175/Q_reg  ( .DIN(g1404), .SDIN(g5151), .SSEL(test_se), .CLK(CK), 
        .Q(g7505), .QN(\DFF_175/net400 ) );
  sdffs1 \DFF_174/Q_reg  ( .DIN(n1384), .SDIN(g5154), .SSEL(test_se), .CLK(CK), 
        .Q(g5151), .QN(n1998) );
  sdffs1 \DFF_173/Q_reg  ( .DIN(n1387), .SDIN(g517), .SSEL(test_se), .CLK(CK), 
        .Q(g5154), .QN(n1989) );
  sdffs1 \DFF_172/Q_reg  ( .DIN(g4651), .SDIN(g3159), .SSEL(test_se), .CLK(CK), 
        .Q(g517) );
  sdffs1 \DFF_171/Q_reg  ( .DIN(g1206), .SDIN(n2400), .SSEL(test_se), .CLK(CK), 
        .Q(g3159), .QN(\DFF_171/net396 ) );
  sdffs1 \DFF_170/Q_reg  ( .DIN(g6319), .SDIN(g4642), .SSEL(test_se), .CLK(CK), 
        .Q(n2400), .QN(n2239) );
  sdffs1 \DFF_169/Q_reg  ( .DIN(g7108), .SDIN(n2399), .SSEL(test_se), .CLK(CK), 
        .Q(g4642), .QN(n1490) );
  sdffs1 \DFF_168/Q_reg  ( .DIN(g5180), .SDIN(n2398), .SSEL(test_se), .CLK(CK), 
        .Q(n2399), .QN(n2257) );
  sdffs1 \DFF_167/Q_reg  ( .DIN(n1381), .SDIN(g7508), .SSEL(test_se), .CLK(CK), 
        .Q(n2398), .QN(n2158) );
  sdffs1 \DFF_166/Q_reg  ( .DIN(g5746), .SDIN(n2397), .SSEL(test_se), .CLK(CK), 
        .Q(g7508) );
  sdffs1 \DFF_165/Q_reg  ( .DIN(n843), .SDIN(g396), .SSEL(test_se), .CLK(CK), 
        .Q(n2397), .QN(n2104) );
  sdffs1 \DFF_164/Q_reg  ( .DIN(g4647), .SDIN(n2396), .SSEL(test_se), .CLK(CK), 
        .Q(g396) );
  sdffs1 \DFF_163/Q_reg  ( .DIN(g6355), .SDIN(n2395), .SSEL(test_se), .CLK(CK), 
        .Q(n2396), .QN(n2203) );
  sdffs1 \DFF_162/Q_reg  ( .DIN(n1381), .SDIN(n2270), .SSEL(test_se), .CLK(CK), 
        .Q(n2395), .QN(n2154) );
  sdffs1 \DFF_161/Q_reg  ( .DIN(g3863), .SDIN(n2394), .SSEL(test_se), .CLK(CK), 
        .Q(n2270) );
  sdffs1 \DFF_160/Q_reg  ( .DIN(g8867), .SDIN(n2291), .SSEL(test_se), .CLK(CK), 
        .Q(n2394), .QN(\DFF_160/net385 ) );
  sdffs1 \DFF_159/Q_reg  ( .DIN(g6875), .SDIN(n2393), .SSEL(test_se), .CLK(CK), 
        .Q(n2291) );
  sdffs1 \DFF_158/Q_reg  ( .DIN(g5169), .SDIN(n2392), .SSEL(test_se), .CLK(CK), 
        .Q(n2393), .QN(n2280) );
  sdffs1 \DFF_157/Q_reg  ( .DIN(n687), .SDIN(g186), .SSEL(test_se), .CLK(CK), 
        .Q(n2392), .QN(n2152) );
  sdffs1 \DFF_156/Q_reg  ( .DIN(g1198), .SDIN(n2391), .SSEL(test_se), .CLK(CK), 
        .Q(g186) );
  sdffs1 \DFF_155/Q_reg  ( .DIN(g6871), .SDIN(g7425), .SSEL(test_se), .CLK(CK), 
        .Q(n2391), .QN(\DFF_155/net380 ) );
  sdffs1 \DFF_154/Q_reg  ( .DIN(n2299), .SDIN(n2390), .SSEL(test_se), .CLK(CK), 
        .Q(g7425) );
  sdffs1 \DFF_153/Q_reg  ( .DIN(g8224), .SDIN(g99), .SSEL(test_se), .CLK(CK), 
        .Q(n2390), .QN(n1460) );
  sdffs1 \DFF_152/Q_reg  ( .DIN(n772), .SDIN(g4643), .SSEL(test_se), .CLK(CK), 
        .Q(g99) );
  sdffs1 \DFF_151/Q_reg  ( .DIN(g6859), .SDIN(g1810), .SSEL(test_se), .CLK(CK), 
        .Q(g4643), .QN(n1477) );
  sdffs1 \DFF_150/Q_reg  ( .DIN(g1817), .SDIN(g355), .SSEL(test_se), .CLK(CK), 
        .Q(g1810), .QN(n1380) );
  sdffs1 \DFF_149/Q_reg  ( .DIN(n739), .SDIN(n2389), .SSEL(test_se), .CLK(CK), 
        .Q(g355) );
  sdffs1 \DFF_148/Q_reg  ( .DIN(g6853), .SDIN(g685), .SSEL(test_se), .CLK(CK), 
        .Q(n2389), .QN(n2133) );
  sdffs1 \DFF_147/Q_reg  ( .DIN(g685), .SDIN(g174), .SSEL(test_se), .CLK(CK), 
        .Q(g685), .QN(n2177) );
  sdffs1 \DFF_146/Q_reg  ( .DIN(g174), .SDIN(n2388), .SSEL(test_se), .CLK(CK), 
        .Q(g174), .QN(n2060) );
  sdffs1 \DFF_145/Q_reg  ( .DIN(n687), .SDIN(n2387), .SSEL(test_se), .CLK(CK), 
        .Q(n2388), .QN(n2139) );
  sdffs1 \DFF_144/Q_reg  ( .DIN(g1871), .SDIN(n2386), .SSEL(test_se), .CLK(CK), 
        .Q(n2387), .QN(\DFF_144/net369 ) );
  sdffs1 \DFF_143/Q_reg  ( .DIN(g8871), .SDIN(n2385), .SSEL(test_se), .CLK(CK), 
        .Q(n2386), .QN(n2048) );
  sdffs1 \DFF_142/Q_reg  ( .DIN(g7512), .SDIN(g583), .SSEL(test_se), .CLK(CK), 
        .Q(n2385), .QN(n1472) );
  sdffs1 \DFF_141/Q_reg  ( .DIN(g3851), .SDIN(n2384), .SSEL(test_se), .CLK(CK), 
        .Q(g583) );
  sdffs1 \DFF_140/Q_reg  ( .DIN(g6883), .SDIN(g1185), .SSEL(test_se), .CLK(CK), 
        .Q(n2384), .QN(\DFF_140/net365 ) );
  sdffs1 \DFF_139/Q_reg  ( .DIN(g1155), .SDIN(n2383), .SSEL(test_se), .CLK(CK), 
        .Q(g1185) );
  sdffs1 \DFF_138/Q_reg  ( .DIN(g7773), .SDIN(n2382), .SSEL(test_se), .CLK(CK), 
        .Q(n2383), .QN(n2062) );
  sdffs1 \DFF_137/Q_reg  ( .DIN(g8226), .SDIN(n2381), .SSEL(test_se), .CLK(CK), 
        .Q(n2382), .QN(g7732) );
  sdffs1 \DFF_136/Q_reg  ( .DIN(g9094), .SDIN(n2380), .SSEL(test_se), .CLK(CK), 
        .Q(n2381), .QN(n2026) );
  sdffs1 \DFF_135/Q_reg  ( .DIN(g1817), .SDIN(n2379), .SSEL(test_se), .CLK(CK), 
        .Q(n2380), .QN(n2249) );
  sdffs1 \DFF_134/Q_reg  ( .DIN(g6340), .SDIN(n1986), .SSEL(test_se), .CLK(CK), 
        .Q(n2379), .QN(n2218) );
  sdffs1 \DFF_133/Q_reg  ( .DIN(g1270), .SDIN(n1384), .SSEL(test_se), .CLK(CK), 
        .Q(n1986) );
  sdffs1 \DFF_131/Q_reg  ( .DIN(g9360), .SDIN(n2378), .SSEL(test_se), .CLK(CK), 
        .Q(n1384), .QN(n1428) );
  sdffs1 \DFF_130/Q_reg  ( .DIN(g9104), .SDIN(n2377), .SSEL(test_se), .CLK(CK), 
        .Q(n2378), .QN(n2016) );
  sdffs1 \DFF_129/Q_reg  ( .DIN(g6313), .SDIN(g1268), .SSEL(test_se), .CLK(CK), 
        .Q(n2377), .QN(n2245) );
  sdffs1 \DFF_128/Q_reg  ( .DIN(g5175), .SDIN(n2376), .SSEL(test_se), .CLK(CK), 
        .Q(g1268) );
  sdffs1 \DFF_127/Q_reg  ( .DIN(n854), .SDIN(g5156), .SSEL(test_se), .CLK(CK), 
        .Q(n2376), .QN(n2129) );
  sdffs1 \DFF_126/Q_reg  ( .DIN(n854), .SDIN(g479), .SSEL(test_se), .CLK(CK), 
        .Q(g5156) );
  sdffs1 \DFF_125/Q_reg  ( .DIN(g4649), .SDIN(n2375), .SSEL(test_se), .CLK(CK), 
        .Q(g479) );
  sdffs1 \DFF_124/Q_reg  ( .DIN(g6317), .SDIN(g200), .SSEL(test_se), .CLK(CK), 
        .Q(n2375), .QN(n2241) );
  sdffs1 \DFF_123/Q_reg  ( .DIN(g199), .SDIN(n2374), .SSEL(test_se), .CLK(CK), 
        .Q(g200) );
  sdffs1 \DFF_122/Q_reg  ( .DIN(g6854), .SDIN(n2373), .SSEL(test_se), .CLK(CK), 
        .Q(n2374), .QN(n1454) );
  sdffs1 \DFF_121/Q_reg  ( .DIN(g8673), .SDIN(g109), .SSEL(test_se), .CLK(CK), 
        .Q(n2373), .QN(n2051) );
  sdffs1 \DFF_120/Q_reg  ( .DIN(n860), .SDIN(g1201), .SSEL(test_se), .CLK(CK), 
        .Q(g109) );
  sdffs1 \DFF_119/Q_reg  ( .DIN(g1200), .SDIN(n2372), .SSEL(test_se), .CLK(CK), 
        .Q(g1201) );
  sdffs1 \DFF_118/Q_reg  ( .DIN(g9100), .SDIN(n2371), .SSEL(test_se), .CLK(CK), 
        .Q(n2372), .QN(n2020) );
  sdffs1 \DFF_117/Q_reg  ( .DIN(g6348), .SDIN(g681), .SSEL(test_se), .CLK(CK), 
        .Q(n2371), .QN(n2210) );
  sdffs1 \DFF_116/Q_reg  ( .DIN(g681), .SDIN(n2370), .SSEL(test_se), .CLK(CK), 
        .Q(g681), .QN(n2176) );
  sdffs1 \DFF_115/Q_reg  ( .DIN(g9103), .SDIN(n2369), .SSEL(test_se), .CLK(CK), 
        .Q(n2370), .QN(n2017) );
  sdffs1 \DFF_114/Q_reg  ( .DIN(n767), .SDIN(n2368), .SSEL(test_se), .CLK(CK), 
        .Q(n2369), .QN(n2163) );
  sdffs1 \DFF_113/Q_reg  ( .DIN(g6341), .SDIN(n2367), .SSEL(test_se), .CLK(CK), 
        .Q(n2368), .QN(n2217) );
  sdffs1 \DFF_112/Q_reg  ( .DIN(g7101), .SDIN(g1309), .SSEL(test_se), .CLK(CK), 
        .Q(n2367), .QN(n1417) );
  sdffs1 \DFF_111/Q_reg  ( .DIN(g1308), .SDIN(n2366), .SSEL(test_se), .CLK(CK), 
        .Q(g1309) );
  sdffs1 \DFF_110/Q_reg  ( .DIN(g7524), .SDIN(g180), .SSEL(test_se), .CLK(CK), 
        .Q(n2366), .QN(n2077) );
  sdffs1 \DFF_109/Q_reg  ( .DIN(g5158), .SDIN(g133), .SSEL(test_se), .CLK(CK), 
        .Q(g180) );
  sdffs1 \DFF_108/Q_reg  ( .DIN(g5149), .SDIN(g113), .SSEL(test_se), .CLK(CK), 
        .Q(g133) );
  sdffs1 \DFF_107/Q_reg  ( .DIN(g5148), .SDIN(n2365), .SSEL(test_se), .CLK(CK), 
        .Q(g113) );
  sdffs1 \DFF_106/Q_reg  ( .DIN(n772), .SDIN(g354), .SSEL(test_se), .CLK(CK), 
        .Q(n2365), .QN(n2111) );
  sdffs1 \DFF_105/Q_reg  ( .DIN(n709), .SDIN(n2364), .SSEL(test_se), .CLK(CK), 
        .Q(g354) );
  sdffs1 \DFF_104/Q_reg  ( .DIN(g7515), .SDIN(g398), .SSEL(test_se), .CLK(CK), 
        .Q(n2364), .QN(n1393) );
  sdffs1 \DFF_103/Q_reg  ( .DIN(g4649), .SDIN(n2363), .SSEL(test_se), .CLK(CK), 
        .Q(g398) );
  sdffs1 \DFF_102/Q_reg  ( .DIN(g5571), .SDIN(n2362), .SSEL(test_se), .CLK(CK), 
        .Q(n2363), .QN(n2276) );
  sdffs1 \DFF_101/Q_reg  ( .DIN(g6868), .SDIN(g3077), .SSEL(test_se), .CLK(CK), 
        .Q(n2362), .QN(\DFF_101/net326 ) );
  sdffs1 \DFF_100/Q_reg  ( .DIN(g2654), .SDIN(g7730), .SSEL(test_se), .CLK(CK), 
        .Q(g3077), .QN(n1446) );
  sdffs1 \DFF_99/Q_reg  ( .DIN(g4658), .SDIN(n2361), .SSEL(test_se), .CLK(CK), 
        .Q(g7730) );
  sdffs1 \DFF_98/Q_reg  ( .DIN(g6392), .SDIN(n2360), .SSEL(test_se), .CLK(CK), 
        .Q(n2361), .QN(\DFF_98/net323 ) );
  sdffs1 \DFF_97/Q_reg  ( .DIN(g6332), .SDIN(n2359), .SSEL(test_se), .CLK(CK), 
        .Q(n2360), .QN(n2226) );
  sdffs1 \DFF_96/Q_reg  ( .DIN(g5745), .SDIN(g646), .SSEL(test_se), .CLK(CK), 
        .Q(n2359), .QN(n2295) );
  sdffs1 \DFF_95/Q_reg  ( .DIN(n1407), .SDIN(n2358), .SSEL(test_se), .CLK(CK), 
        .Q(g646) );
  sdffs1 \DFF_94/Q_reg  ( .DIN(g6841), .SDIN(g1012), .SSEL(test_se), .CLK(CK), 
        .Q(n2358), .QN(n2136) );
  sdffs1 \DFF_93/Q_reg  ( .DIN(g43), .SDIN(n2357), .SSEL(test_se), .CLK(CK), 
        .Q(g1012) );
  sdffs1 \DFF_92/Q_reg  ( .DIN(n772), .SDIN(g7504), .SSEL(test_se), .CLK(CK), 
        .Q(n2357), .QN(n2125) );
  sdffs1 \DFF_91/Q_reg  ( .DIN(g7308), .SDIN(n1996), .SSEL(test_se), .CLK(CK), 
        .Q(g7504) );
  sdffs1 \DFF_90/Q_reg  ( .DIN(n1525), .SDIN(g587), .SSEL(test_se), .CLK(CK), 
        .Q(n1996) );
  sdffs1 \DFF_89/Q_reg  ( .DIN(g3852), .SDIN(n1386), .SSEL(test_se), .CLK(CK), 
        .Q(g587) );
  sdffs1 \DFF_87/Q_reg  ( .DIN(g9373), .SDIN(g3847), .SSEL(test_se), .CLK(CK), 
        .Q(n1386), .QN(n1412) );
  sdffs1 \DFF_86/Q_reg  ( .DIN(g7304), .SDIN(n2356), .SSEL(test_se), .CLK(CK), 
        .Q(g3847), .QN(n2262) );
  sdffs1 \DFF_85/Q_reg  ( .DIN(g5187), .SDIN(n2355), .SSEL(test_se), .CLK(CK), 
        .Q(n2356), .QN(n2282) );
  sdffs1 \DFF_84/Q_reg  ( .DIN(g6878), .SDIN(n2354), .SSEL(test_se), .CLK(CK), 
        .Q(n2355), .QN(\DFF_84/net309 ) );
  sdffs1 \DFF_83/Q_reg  ( .DIN(n1381), .SDIN(n2353), .SSEL(test_se), .CLK(CK), 
        .Q(n2354), .QN(n2112) );
  sdffs1 \DFF_82/Q_reg  ( .DIN(g7759), .SDIN(n2352), .SSEL(test_se), .CLK(CK), 
        .Q(n2353), .QN(n2090) );
  sdffs1 \DFF_81/Q_reg  ( .DIN(g6356), .SDIN(n2351), .SSEL(test_se), .CLK(CK), 
        .Q(n2352), .QN(n2202) );
  sdffs1 \DFF_80/Q_reg  ( .DIN(g6855), .SDIN(n2350), .SSEL(test_se), .CLK(CK), 
        .Q(n2351), .QN(n2132) );
  sdffs1 \DFF_79/Q_reg  ( .DIN(g7519), .SDIN(g295), .SSEL(test_se), .CLK(CK), 
        .Q(n2350), .QN(n2076) );
  sdffs1 \DFF_78/Q_reg  ( .DIN(g4642), .SDIN(g730), .SSEL(test_se), .CLK(CK), 
        .Q(g295) );
  sdffs1 \DFF_77/Q_reg  ( .DIN(g730), .SDIN(g710), .SSEL(test_se), .CLK(CK), 
        .Q(g730), .QN(n2182) );
  sdffs1 \DFF_76/Q_reg  ( .DIN(g710), .SDIN(n2349), .SSEL(test_se), .CLK(CK), 
        .Q(g710), .QN(n2187) );
  sdffs1 \DFF_75/Q_reg  ( .DIN(n2304), .SDIN(n2348), .SSEL(test_se), .CLK(CK), 
        .Q(n2349), .QN(n2148) );
  sdffs1 \DFF_74/Q_reg  ( .DIN(g9092), .SDIN(g4316), .SSEL(test_se), .CLK(CK), 
        .Q(n2348), .QN(n2028) );
  sdffs1 \DFF_73/Q_reg  ( .DIN(g890), .SDIN(n2347), .SSEL(test_se), .CLK(CK), 
        .Q(g4316), .QN(n2281) );
  sdffs1 \DFF_72/Q_reg  ( .DIN(g9093), .SDIN(n1381), .SSEL(test_se), .CLK(CK), 
        .Q(n2347), .QN(n2027) );
  sdffs1 \DFF_71/Q_reg  ( .DIN(g9362), .SDIN(n2346), .SSEL(test_se), .CLK(CK), 
        .Q(n1381), .QN(n1413) );
  sdffs1 \DFF_70/Q_reg  ( .DIN(n860), .SDIN(g179), .SSEL(test_se), .CLK(CK), 
        .Q(n2346), .QN(n2165) );
  sdffs1 \DFF_69/Q_reg  ( .DIN(g5159), .SDIN(n2286), .SSEL(test_se), .CLK(CK), 
        .Q(g179) );
  sdffs1 \DFF_68/Q_reg  ( .DIN(g6888), .SDIN(g3851), .SSEL(test_se), .CLK(CK), 
        .Q(n2286) );
  sdffs1 \DFF_67/Q_reg  ( .DIN(g7527), .SDIN(g4372), .SSEL(test_se), .CLK(CK), 
        .Q(g3851), .QN(n2263) );
  sdffs1 \DFF_66/Q_reg  ( .DIN(g4370), .SDIN(n2345), .SSEL(test_se), .CLK(CK), 
        .Q(g4372), .QN(\DFF_66/net291 ) );
  sdffs1 \DFF_65/Q_reg  ( .DIN(n1385), .SDIN(g718), .SSEL(test_se), .CLK(CK), 
        .Q(n2345), .QN(n2116) );
  sdffs1 \DFF_64/Q_reg  ( .DIN(g718), .SDIN(n2344), .SSEL(test_se), .CLK(CK), 
        .Q(g718), .QN(n2183) );
  sdffs1 \DFF_63/Q_reg  ( .DIN(g6880), .SDIN(n2343), .SSEL(test_se), .CLK(CK), 
        .Q(n2344), .QN(\DFF_63/net288 ) );
  sdffs1 \DFF_62/Q_reg  ( .DIN(g6323), .SDIN(n2342), .SSEL(test_se), .CLK(CK), 
        .Q(n2343), .QN(n2235) );
  sdffs1 \DFF_61/Q_reg  ( .DIN(g1911), .SDIN(n2341), .SSEL(test_se), .CLK(CK), 
        .Q(n2342), .QN(n2056) );
  sdffs1 \DFF_60/Q_reg  ( .DIN(g9110), .SDIN(g137), .SSEL(test_se), .CLK(CK), 
        .Q(n2341), .QN(n2010) );
  sdffs1 \DFF_59/Q_reg  ( .DIN(g5150), .SDIN(g117), .SSEL(test_se), .CLK(CK), 
        .Q(g137) );
  sdffs1 \DFF_58/Q_reg  ( .DIN(g5153), .SDIN(g984), .SSEL(test_se), .CLK(CK), 
        .Q(g117) );
  sdffs1 \DFF_57/Q_reg  ( .DIN(g9133), .SDIN(g1014), .SSEL(test_se), .CLK(CK), 
        .Q(g984) );
  sdffs1 \DFF_56/Q_reg  ( .DIN(g1012), .SDIN(g1783), .SSEL(test_se), .CLK(CK), 
        .Q(g1014) );
  sdffs1 \DFF_55/Q_reg  ( .DIN(g3855), .SDIN(n2340), .SSEL(test_se), .CLK(CK), 
        .Q(g1783), .QN(n1379) );
  sdffs1 \DFF_54/Q_reg  ( .DIN(n772), .SDIN(g1817), .SSEL(test_se), .CLK(CK), 
        .Q(n2340), .QN(n2168) );
  sdffs1 \DFF_53/Q_reg  ( .DIN(g1824), .SDIN(g455), .SSEL(test_se), .CLK(CK), 
        .Q(g1817), .QN(n1421) );
  sdffs1 \DFF_52/Q_reg  ( .DIN(n755), .SDIN(g315), .SSEL(test_se), .CLK(CK), 
        .Q(g455) );
  sdffs1 \DFF_51/Q_reg  ( .DIN(g4647), .SDIN(n2339), .SSEL(test_se), .CLK(CK), 
        .Q(g315) );
  sdffs1 \DFF_50/Q_reg  ( .DIN(g1810), .SDIN(n2338), .SSEL(test_se), .CLK(CK), 
        .Q(n2339), .QN(n2256) );
  sdffs1 \DFF_49/Q_reg  ( .DIN(g7757), .SDIN(n2337), .SSEL(test_se), .CLK(CK), 
        .Q(n2338), .QN(n1463) );
  sdffs1 \DFF_48/Q_reg  ( .DIN(n2304), .SDIN(n2336), .SSEL(test_se), .CLK(CK), 
        .Q(n2337), .QN(n2142) );
  sdffs1 \DFF_47/Q_reg  ( .DIN(g9105), .SDIN(n2335), .SSEL(test_se), .CLK(CK), 
        .Q(n2336), .QN(n2015) );
  sdffs1 \DFF_46/Q_reg  ( .DIN(n860), .SDIN(g1269), .SSEL(test_se), .CLK(CK), 
        .Q(n2335), .QN(n2118) );
  sdffs1 \DFF_45/Q_reg  ( .DIN(g5740), .SDIN(n2334), .SSEL(test_se), .CLK(CK), 
        .Q(g1269) );
  sdffs1 \DFF_44/Q_reg  ( .DIN(g5185), .SDIN(n2333), .SSEL(test_se), .CLK(CK), 
        .Q(n2334), .QN(n1452) );
  sdffs1 \DFF_43/Q_reg  ( .DIN(n854), .SDIN(n2332), .SSEL(test_se), .CLK(CK), 
        .Q(n2333), .QN(n1444) );
  sdffs1 \DFF_42/Q_reg  ( .DIN(g7772), .SDIN(n2331), .SSEL(test_se), .CLK(CK), 
        .Q(n2332), .QN(n2068) );
  sdffs1 \DFF_41/Q_reg  ( .DIN(g6318), .SDIN(n2330), .SSEL(test_se), .CLK(CK), 
        .Q(n2331), .QN(n2240) );
  sdffs1 \DFF_40/Q_reg  ( .DIN(g1312), .SDIN(g1798), .SSEL(test_se), .CLK(CK), 
        .Q(n2330), .QN(n1422) );
  sdffs1 \DFF_39/Q_reg  ( .DIN(g1804), .SDIN(n2329), .SSEL(test_se), .CLK(CK), 
        .Q(g1798), .QN(n1395) );
  sdffs1 \DFF_38/Q_reg  ( .DIN(n860), .SDIN(n2328), .SSEL(test_se), .CLK(CK), 
        .Q(n2329), .QN(n2145) );
  sdffs1 \DFF_37/Q_reg  ( .DIN(g6352), .SDIN(g1205), .SSEL(test_se), .CLK(CK), 
        .Q(n2328), .QN(n2206) );
  sdffs1 \DFF_36/Q_reg  ( .DIN(g1204), .SDIN(n2327), .SSEL(test_se), .CLK(CK), 
        .Q(g1205) );
  sdffs1 \DFF_35/Q_reg  ( .DIN(n860), .SDIN(n2302), .SSEL(test_se), .CLK(CK), 
        .Q(n2327), .QN(n2126) );
  sdffs1 \DFF_33/Q_reg  ( .DIN(g9036), .SDIN(g294), .SSEL(test_se), .CLK(CK), 
        .Q(n2326), .QN(n2061) );
  sdffs1 \DFF_32/Q_reg  ( .DIN(n728), .SDIN(g2659), .SSEL(test_se), .CLK(CK), 
        .Q(g294) );
  sdffs1 \DFF_31/Q_reg  ( .DIN(g5571), .SDIN(n2325), .SSEL(test_se), .CLK(CK), 
        .Q(g2659), .QN(n1400) );
  sdffs1 \DFF_30/Q_reg  ( .DIN(g7767), .SDIN(g393), .SSEL(test_se), .CLK(CK), 
        .Q(n2325), .QN(n2130) );
  sdffs1 \DFF_29/Q_reg  ( .DIN(g4644), .SDIN(n2324), .SSEL(test_se), .CLK(CK), 
        .Q(g393) );
  sdffs1 \DFF_28/Q_reg  ( .DIN(n767), .SDIN(g2672), .SSEL(test_se), .CLK(CK), 
        .Q(n2324), .QN(n2146) );
  sdffs1 \DFF_27/Q_reg  ( .DIN(g3863), .SDIN(g7506), .SSEL(test_se), .CLK(CK), 
        .Q(g2672), .QN(n1399) );
  sdffs1 \DFF_26/Q_reg  ( .DIN(g6386), .SDIN(n2323), .SSEL(test_se), .CLK(CK), 
        .Q(g7506) );
  sdffs1 \DFF_25/Q_reg  ( .DIN(g6865), .SDIN(n2322), .SSEL(test_se), .CLK(CK), 
        .Q(n2323), .QN(n1408) );
  sdffs1 \DFF_24/Q_reg  ( .DIN(g6881), .SDIN(n2321), .SSEL(test_se), .CLK(CK), 
        .Q(n2322), .QN(\DFF_24/net249 ) );
  sdffs1 \DFF_23/Q_reg  ( .DIN(g6336), .SDIN(n2320), .SSEL(test_se), .CLK(CK), 
        .Q(n2321), .QN(n2222) );
  sdffs1 \DFF_22/Q_reg  ( .DIN(g6291), .SDIN(n2319), .SSEL(test_se), .CLK(CK), 
        .Q(n2320), .QN(n1988) );
  sdffs1 \DFF_21/Q_reg  ( .DIN(g6371), .SDIN(n2318), .SSEL(test_se), .CLK(CK), 
        .Q(n2319), .QN(g6895) );
  sdffs1 \DFF_20/Q_reg  ( .DIN(g6869), .SDIN(n2317), .SSEL(test_se), .CLK(CK), 
        .Q(n2318), .QN(\DFF_20/net245 ) );
  sdffs1 \DFF_19/Q_reg  ( .DIN(n1385), .SDIN(g292), .SSEL(test_se), .CLK(CK), 
        .Q(n2317), .QN(n2143) );
  sdffs1 \DFF_18/Q_reg  ( .DIN(g4639), .SDIN(g535), .SSEL(test_se), .CLK(CK), 
        .Q(g292) );
  sdffs1 \DFF_17/Q_reg  ( .DIN(g3844), .SDIN(g5159), .SSEL(test_se), .CLK(CK), 
        .Q(g535) );
  sdffs1 \DFF_16/Q_reg  ( .DIN(g5731), .SDIN(g454), .SSEL(test_se), .CLK(CK), 
        .Q(g5159) );
  sdffs1 \DFF_15/Q_reg  ( .DIN(g4639), .SDIN(n2316), .SSEL(test_se), .CLK(CK), 
        .Q(g454) );
  sdffs1 \DFF_14/Q_reg  ( .DIN(g7520), .SDIN(g314), .SSEL(test_se), .CLK(CK), 
        .Q(n2316), .QN(n1441) );
  sdffs1 \DFF_13/Q_reg  ( .DIN(g4646), .SDIN(n2315), .SSEL(test_se), .CLK(CK), 
        .Q(g314) );
  sdffs1 \DFF_12/Q_reg  ( .DIN(g9111), .SDIN(g976), .SSEL(test_se), .CLK(CK), 
        .Q(n2315), .QN(n2009) );
  sdffs1 \DFF_11/Q_reg  ( .DIN(g8864), .SDIN(n2314), .SSEL(test_se), .CLK(CK), 
        .Q(g976) );
  sdffs1 \DFF_10/Q_reg  ( .DIN(g5735), .SDIN(g1153), .SSEL(test_se), .CLK(CK), 
        .Q(n2314), .QN(n2292) );
  sdffs1 \DFF_9/Q_reg  ( .DIN(g6856), .SDIN(g5161), .SSEL(test_se), .CLK(CK), 
        .Q(g1153) );
  sdffs1 \DFF_7/Q_reg  ( .DIN(g5733), .SDIN(n2313), .SSEL(test_se), .CLK(CK), 
        .Q(g5161) );
  sdffs1 \DFF_6/Q_reg  ( .DIN(n2304), .SDIN(g948), .SSEL(test_se), .CLK(CK), 
        .Q(n2313), .QN(n2162) );
  sdffs1 \DFF_5/Q_reg  ( .DIN(g8664), .SDIN(g452), .SSEL(test_se), .CLK(CK), 
        .Q(g948) );
  sdffs1 \DFF_4/Q_reg  ( .DIN(g3159), .SDIN(g273), .SSEL(test_se), .CLK(CK), 
        .Q(g452) );
  sdffs1 \DFF_3/Q_reg  ( .DIN(g4650), .SDIN(g312), .SSEL(test_se), .CLK(CK), 
        .Q(g273) );
  sdffs1 \DFF_2/Q_reg  ( .DIN(n746), .SDIN(g1271), .SSEL(test_se), .CLK(CK), 
        .Q(g312) );
  sdffs1 \DFF_1/Q_reg  ( .DIN(n2297), .SDIN(g397), .SSEL(test_se), .CLK(CK), 
        .Q(g1271) );
  sdffs1 \DFF_0/Q_reg  ( .DIN(g4648), .SDIN(test_si), .SSEL(test_se), .CLK(CK), 
        .Q(g397) );
  sdffs1 \DFF_34/Q_reg  ( .DIN(g9372), .SDIN(n2326), .SSEL(test_se), .CLK(CK), 
        .Q(n2302) );
  nor2s1 troj1_0U1 ( .DIN1(troj1_0n1), .DIN2(troj1_0n2), .Q(Trigger_en1_0) );
  nnd4s1 troj1_0U2 ( .DIN1(n1522), .DIN2(n1309), .DIN3(n1954), .DIN4(troj1_0n3), .Q(troj1_0n2) );
  and4s1 troj1_0U3 ( .DIN1(n1092), .DIN2(g7528), .DIN3(g5163), .DIN4(troj1_0n4), .Q(troj1_0n3) );
  i1s1 troj1_0U4 ( .DIN(g6354), .Q(troj1_0n4) );
  or5s1 troj1_0U5 ( .DIN1(g9105), .DIN2(g7109), .DIN3(n1377), .DIN4(n1310), .DIN5(troj1_0n5),         .Q(troj1_0n1) );
  nnd2s1 troj1_0U6 ( .DIN1(troj1_0n6), .DIN2(troj1_0n7), .Q(troj1_0n5) );
  nor2s1 troj1_0U7 ( .DIN1(n782), .DIN2(n680), .Q(troj1_0n7) );
  nor2s1 troj1_0U8 ( .DIN1(n650), .DIN2(n1554), .Q(troj1_0n6) );
    xor2s1 trojan1_0  (.DIN1(tempg9027), .DIN2(Trigger_en1_0), .Q(g9027) );
  nor5s1 troj1_1U1 ( .DIN1(troj1_1n1), .DIN2(troj1_1n2), .DIN3(g9086), .DIN4(n1363), .DIN5(n1348),         .Q(Trigger_en1_1) );
  i1s1 troj1_1U2 ( .DIN(troj1_1n3), .Q(troj1_1n2) );
  nor4s1 troj1_1U3 ( .DIN1(n751), .DIN2(n738), .DIN3(n1879), .DIN4(n1643), .Q(troj1_1n3) );
  nnd4s1 troj1_1U4 ( .DIN1(n1126), .DIN2(g6877), .DIN3(troj1_1n4), .DIN4(troj1_1n5), .Q(troj1_1n1) );
  and3s1 troj1_1U5 ( .DIN1(n1691), .DIN2(n1671), .DIN3(n660), .Q(troj1_1n5) );
  nor2s1 troj1_1U6 ( .DIN1(g8678), .DIN2(g6857), .Q(troj1_1n4) );
    xor2s1 trojan1_1  (.DIN1(tempg9112), .DIN2(Trigger_en1_1), .Q(g9112) );

endmodule

