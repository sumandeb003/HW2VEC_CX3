module c6288 (N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426,
N443, N460, N477, N494, N511, N528, N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288);

input N1, N18, N35, N52, N69, N86, N103, N120, N137, N154, N171, N188, N205, N222, N239, N256, N273, N290, N307, N324, N341, N358, N375, N392, N409, N426, N443, N460, N477, N494, N511, N528;

output N545, N1581, N1901, N2223, N2548, N2877, N3211, N3552, N3895, N4241, N4591, N4946, N5308, N5672, N5971, N6123, N6150, N6160, N6170, N6180, N6190, N6200, N6210, N6220, N6230, N6240, N6250, N6260, N6270, N6280, N6287, N6288;

wire N546, N549, N552, N555, N558, N561, N564, N567, N570, N573, N576, N579, N582, N585, N588, N591, N594, N597, N600, N603, N606, N609, N612, N615, N618, N621, N624, N627, N630, N633, N636, N639, N642, N645, N648, N651, N654, N657, N660, N663, N666, N669, N672, N675, N678, N681, N684, N687, N690, N693, N696, N699, N702, N705, N708, N711, N714, N717, N720, N723, N726, N729, N732, N735, N738, N741, N744, N747, N750, N753, N756, N759, N762, N765, N768, N771, N774, N777, N780, N783, N786, N789, N792, N795, N798, N801, N804, N807, N810, N813, N816, N819, N822, N825, N828, N831, N834, N837, N840, N843, N846, N849, N852, N855, N858, N861, N864, N867, N870, N873, N876, N879, N882, N885, N888, N891, N894, N897, N900, N903, N906, N909, N912, N915, N918, N921, N924, N927, N930, N933, N936, N939, N942, N945, N948, N951, N954, N957, N960, N963, N966, N969, N972, N975, N978, N981, N984, N987, N990, N993, N996, N999, N1002, N1005, N1008, N1011, N1014, N1017, N1020, N1023, N1026, N1029, N1032, N1035, N1038, N1041, N1044, N1047, N1050, N1053, N1056, N1059, N1062, N1065, N1068, N1071, N1074, N1077, N1080, N1083, N1086, N1089, N1092, N1095, N1098, N1101, N1104, N1107, N1110, N1113, N1116, N1119, N1122, N1125, N1128, N1131, N1134, N1137, N1140, N1143, N1146, N1149, N1152, N1155, N1158, N1161, N1164, N1167, N1170, N1173, N1176, N1179, N1182, N1185, N1188, N1191, N1194, N1197, N1200, N1203, N1206, N1209, N1212, N1215, N1218, N1221, N1224, N1227, N1230, N1233, N1236, N1239, N1242, N1245, N1248, N1251, N1254, N1257, N1260, N1263, N1266, N1269, N1272, N1275, N1278, N1281, N1284, N1287, N1290, N1293, N1296, N1299, N1302, N1305, N1308, N1311, N1315, N1319, N1323, N1327, N1331, N1335, N1339, N1343, N1347, N1351, N1355, N1359, N1363, N1367, N1371, N1372, N1373, N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383, N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1404, N1407, N1410, N1413, N1416, N1419, N1422, N1425, N1428, N1431, N1434, N1437, N1440, N1443, N1446, N1450, N1454, N1458, N1462, N1466, N1470, N1474, N1478, N1482, N1486, N1490, N1494, N1498, N1502, N1506, N1507, N1508, N1511, N1512, N1513, N1516, N1517, N1518, N1521, N1522, N1523, N1526, N1527, N1528, N1531, N1532, N1533, N1536, N1537, N1538, N1541, N1542, N1543, N1546, N1547, N1548, N1551, N1552, N1553, N1556, N1557, N1558, N1561, N1562, N1563, N1566, N1567, N1568, N1571, N1572, N1573, N1576, N1577, N1578, N1582, N1585, N1588, N1591, N1594, N1597, N1600, N1603, N1606, N1609, N1612, N1615, N1618, N1621, N1624, N1628, N1632, N1636, N1640, N1644, N1648, N1652, N1656, N1660, N1664, N1668, N1672, N1676, N1680, N1684, N1685, N1686, N1687, N1688, N1689, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1697, N1698, N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708, N1709, N1710, N1711, N1712, N1713, N1714, N1717, N1720, N1723, N1726, N1729, N1732, N1735, N1738, N1741, N1744, N1747, N1750, N1753, N1756, N1759, N1763, N1767, N1771, N1775, N1779, N1783, N1787, N1791, N1795, N1799, N1803, N1807, N1811, N1815, N1819, N1820, N1821, N1824, N1825, N1826, N1829, N1830, N1831, N1834, N1835, N1836, N1839, N1840, N1841, N1844, N1845, N1846, N1849, N1850, N1851, N1854, N1855, N1856, N1859, N1860, N1861, N1864, N1865, N1866, N1869, N1870, N1871, N1874, N1875, N1876, N1879, N1880, N1881, N1884, N1885, N1886, N1889, N1890, N1891, N1894, N1897, N1902, N1905, N1908, N1911, N1914, N1917, N1920, N1923, N1926, N1929, N1932, N1935, N1938, N1941, N1945, N1946, N1947, N1951, N1955, N1959, N1963, N1967, N1971, N1975, N1979, N1983, N1987, N1991, N1995, N1999, N2000, N2001, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012, N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022, N2023, N2024, N2025, N2026, N2027, N2028, N2029, N2030, N2033, N2037, N2040, N2043, N2046, N2049, N2052, N2055, N2058, N2061, N2064, N2067, N2070, N2073, N2076, N2080, N2081, N2082, N2085, N2089, N2093, N2097, N2101, N2105, N2109, N2113, N2117, N2121, N2125, N2129, N2133, N2137, N2138, N2139, N2142, N2145, N2149, N2150, N2151, N2154, N2155, N2156, N2159, N2160, N2161, N2164, N2165, N2166, N2169, N2170, N2171, N2174, N2175, N2176, N2179, N2180, N2181, N2184, N2185, N2186, N2189, N2190, N2191, N2194, N2195, N2196, N2199, N2200, N2201, N2204, N2205, N2206, N2209, N2210, N2211, N2214, N2217, N2221, N2222, N2224, N2227, N2230, N2233, N2236, N2239, N2242, N2245, N2248, N2251, N2254, N2257, N2260, N2264, N2265, N2266, N2269, N2273, N2277, N2281, N2285, N2289, N2293, N2297, N2301, N2305, N2309, N2313, N2317, N2318, N2319, N2322, N2326, N2327, N2328, N2329, N2330, N2331, N2332, N2333, N2334, N2335, N2336, N2337, N2338, N2339, N2340, N2341, N2342, N2343, N2344, N2345, N2346, N2347, N2348, N2349, N2350, N2353, N2357, N2358, N2359, N2362, N2365, N2368, N2371, N2374, N2377, N2380, N2383, N2386, N2389, N2392, N2395, N2398, N2402, N2403, N2404, N2407, N2410, N2414, N2418, N2422, N2426, N2430, N2434, N2438, N2442, N2446, N2450, N2454, N2458, N2462, N2463, N2464, N2467, N2470, N2474, N2475, N2476, N2477, N2478, N2481, N2482, N2483, N2486, N2487, N2488, N2491, N2492, N2493, N2496, N2497, N2498, N2501, N2502, N2503, N2506, N2507, N2508, N2511, N2512, N2513, N2516, N2517, N2518, N2521, N2522, N2523, N2526, N2527, N2528, N2531, N2532, N2533, N2536, N2539, N2543, N2544, N2545, N2549, N2552, N2555, N2558, N2561, N2564, N2567, N2570, N2573, N2576, N2579, N2582, N2586, N2587, N2588, N2591, N2595, N2599, N2603, N2607, N2611, N2615, N2619, N2623, N2627, N2631, N2635, N2639, N2640, N2641, N2644, N2648, N2649, N2650, N2653, N2654, N2655, N2656, N2657, N2658, N2659, N2660, N2661, N2662, N2663, N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673, N2674, N2675, N2678, N2682, N2683, N2684, N2687, N2690, N2694, N2697, N2700, N2703, N2706, N2709, N2712, N2715, N2718, N2721, N2724, N2727, N2731, N2732, N2733, N2736, N2739, N2743, N2744, N2745, N2749, N2753, N2757, N2761, N2765, N2769, N2773, N2777, N2781, N2785, N2789, N2790, N2791, N2794, N2797, N2801, N2802, N2803, N2806, N2807, N2808, N2811, N2812, N2813, N2816, N2817, N2818, N2821, N2822, N2823, N2826, N2827, N2828, N2831, N2832, N2833, N2836, N2837, N2838, N2841, N2842, N2843, N2846, N2847, N2848, N2851, N2852, N2853, N2856, N2857, N2858, N2861, N2864, N2868, N2869, N2870, N2873, N2878, N2881, N2884, N2887, N2890, N2893, N2896, N2899, N2902, N2905, N2908, N2912, N2913, N2914, N2917, N2921, N2922, N2923, N2926, N2930, N2934, N2938, N2942, N2946, N2950, N2954, N2958, N2962, N2966, N2967, N2968, N2971, N2975, N2976, N2977, N2980, N2983, N2987, N2988, N2989, N2990, N2991, N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001, N3002, N3003, N3004, N3005, N3006, N3007, N3010, N3014, N3015, N3016, N3019, N3022, N3026, N3027, N3028, N3031, N3034, N3037, N3040, N3043, N3046, N3049, N3052, N3055, N3058, N3062, N3063, N3064, N3067, N3070, N3074, N3075, N3076, N3079, N3083, N3087, N3091, N3095, N3099, N3103, N3107, N3111, N3115, N3119, N3120, N3121, N3124, N3127, N3131, N3132, N3133, N3136, N3140, N3141, N3142, N3145, N3146, N3147, N3150, N3151, N3152, N3155, N3156, N3157, N3160, N3161, N3162, N3165, N3166, N3167, N3170, N3171, N3172, N3175, N3176, N3177, N3180, N3181, N3182, N3185, N3186, N3187, N3190, N3193, N3197, N3198, N3199, N3202, N3206, N3207, N3208, N3212, N3215, N3218, N3221, N3224, N3227, N3230, N3233, N3236, N3239, N3243, N3244, N3245, N3248, N3252, N3253, N3254, N3257, N3260, N3264, N3268, N3272, N3276, N3280, N3284, N3288, N3292, N3296, N3300, N3301, N3302, N3305, N3309, N3310, N3311, N3314, N3317, N3321, N3322, N3323, N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334, N3335, N3336, N3337, N3338, N3339, N3340, N3341, N3344, N3348, N3349, N3350, N3353, N3356, N3360, N3361, N3362, N3365, N3368, N3371, N3374, N3377, N3380, N3383, N3386, N3389, N3392, N3396, N3397, N3398, N3401, N3404, N3408, N3409, N3410, N3413, N3417, N3421, N3425, N3429, N3433, N3437, N3441, N3445, N3449, N3453, N3454, N3455, N3458, N3461, N3465, N3466, N3467, N3470, N3474, N3475, N3476, N3479, N3480, N3481, N3484, N3485, N3486, N3489, N3490, N3491, N3494, N3495, N3496, N3499, N3500, N3501, N3504, N3505, N3506, N3509, N3510, N3511, N3514, N3515, N3516, N3519, N3520, N3521, N3524, N3527, N3531, N3532, N3533, N3536, N3540, N3541, N3542, N3545, N3548, N3553, N3556, N3559, N3562, N3565, N3568, N3571, N3574, N3577, N3581, N3582, N3583, N3586, N3590, N3591, N3592, N3595, N3598, N3602, N3603, N3604, N3608, N3612, N3616, N3620, N3624, N3628, N3632, N3636, N3637, N3638, N3641, N3645, N3646, N3647, N3650, N3653, N3657, N3658, N3659, N3662, N3663, N3664, N3665, N3666, N3667, N3668, N3669, N3670, N3671, N3672, N3673, N3674, N3675, N3676, N3677, N3678, N3681, N3685, N3686, N3687, N3690, N3693, N3697, N3698, N3699, N3702, N3706, N3709, N3712, N3715, N3718, N3721, N3724, N3727, N3730, N3734, N3735, N3736, N3739, N3742, N3746, N3747, N3748, N3751, N3755, N3756, N3757, N3760, N3764, N3768, N3772, N3776, N3780, N3784, N3788, N3792, N3793, N3794, N3797, N3800, N3804, N3805, N3806, N3809, N3813, N3814, N3815, N3818, N3821, N3825, N3826, N3827, N3830, N3831, N3832, N3835, N3836, N3837, N3840, N3841, N3842, N3845, N3846, N3847, N3850, N3851, N3852, N3855, N3856, N3857, N3860, N3861, N3862, N3865, N3868, N3872, N3873, N3874, N3877, N3881, N3882, N3883, N3886, N3889, N3893, N3894, N3896, N3899, N3902, N3905, N3908, N3911, N3914, N3917, N3921, N3922, N3923, N3926, N3930, N3931, N3932, N3935, N3938, N3942, N3943, N3944, N3947, N3951, N3955, N3959, N3963, N3967, N3971, N3975, N3976, N3977, N3980, N3984, N3985, N3986, N3989, N3992, N3996, N3997, N3998, N4001, N4005, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014, N4015, N4016, N4017, N4018, N4019, N4022, N4026, N4027, N4028, N4031, N4034, N4038, N4039, N4040, N4043, N4047, N4048, N4049, N4052, N4055, N4058, N4061, N4064, N4067, N4070, N4073, N4077, N4078, N4079, N4082, N4085, N4089, N4090, N4091, N4094, N4098, N4099, N4100, N4103, N4106, N4110, N4114, N4118, N4122, N4126, N4130, N4134, N4138, N4139, N4140, N4143, N4146, N4150, N4151, N4152, N4155, N4159, N4160, N4161, N4164, N4167, N4171, N4172, N4173, N4174, N4175, N4178, N4179, N4180, N4183, N4184, N4185, N4188, N4189, N4190, N4193, N4194, N4195, N4198, N4199, N4200, N4203, N4204, N4205, N4208, N4211, N4215, N4216, N4217, N4220, N4224, N4225, N4226, N4229, N4232, N4236, N4237, N4238, N4242, N4245, N4248, N4251, N4254, N4257, N4260, N4264, N4265, N4266, N4269, N4273, N4274, N4275, N4278, N4281, N4285, N4286, N4287, N4290, N4294, N4298, N4302, N4306, N4310, N4314, N4318, N4319, N4320, N4323, N4327, N4328, N4329, N4332, N4335, N4339, N4340, N4341, N4344, N4348, N4349, N4350, N4353, N4354, N4355, N4356, N4357, N4358, N4359, N4360, N4361, N4362, N4363, N4364, N4365, N4368, N4372, N4373, N4374, N4377, N4380, N4384, N4385, N4386, N4389, N4393, N4394, N4395, N4398, N4401, N4405, N4408, N4411, N4414, N4417, N4420, N4423, N4427, N4428, N4429, N4432, N4435, N4439, N4440, N4441, N4444, N4448, N4449, N4450, N4453, N4456, N4460, N4461, N4462, N4466, N4470, N4474, N4478, N4482, N4486, N4487, N4488, N4491, N4494, N4498, N4499, N4500, N4503, N4507, N4508, N4509, N4512, N4515, N4519, N4520, N4521, N4524, N4525, N4526, N4529, N4530, N4531, N4534, N4535, N4536, N4539, N4540, N4541, N4544, N4545, N4546, N4549, N4550, N4551, N4554, N4557, N4561, N4562, N4563, N4566, N4570, N4571, N4572, N4575, N4578, N4582, N4583, N4584, N4587, N4592, N4595, N4598, N4601, N4604, N4607, N4611, N4612, N4613, N4616, N4620, N4621, N4622, N4625, N4628, N4632, N4633, N4634, N4637, N4641, N4642, N4643, N4646, N4650, N4654, N4658, N4662, N4666, N4667, N4668, N4671, N4675, N4676, N4677, N4680, N4683, N4687, N4688, N4689, N4692, N4696, N4697, N4698, N4701, N4704, N4708, N4709, N4710, N4711, N4712, N4713, N4714, N4715, N4716, N4717, N4718, N4721, N4725, N4726, N4727, N4730, N4733, N4737, N4738, N4739, N4742, N4746, N4747, N4748, N4751, N4754, N4758, N4759, N4760, N4763, N4766, N4769, N4772, N4775, N4779, N4780, N4781, N4784, N4787, N4791, N4792, N4793, N4796, N4800, N4801, N4802, N4805, N4808, N4812, N4813, N4814, N4817, N4821, N4825, N4829, N4833, N4837, N4838, N4839, N4842, N4845, N4849, N4850, N4851, N4854, N4858, N4859, N4860, N4863, N4866, N4870, N4871, N4872, N4875, N4879, N4880, N4881, N4884, N4885, N4886, N4889, N4890, N4891, N4894, N4895, N4896, N4899, N4900, N4901, N4904, N4907, N4911, N4912, N4913, N4916, N4920, N4921, N4922, N4925, N4928, N4932, N4933, N4934, N4937, N4941, N4942, N4943, N4947, N4950, N4953, N4956, N4959, N4963, N4964, N4965, N4968, N4972, N4973, N4974, N4977, N4980, N4984, N4985, N4986, N4989, N4993, N4994, N4995, N4998, N5001, N5005, N5009, N5013, N5017, N5021, N5022, N5023, N5026, N5030, N5031, N5032, N5035, N5038, N5042, N5043, N5044, N5047, N5051, N5052, N5053, N5056, N5059, N5063, N5064, N5065, N5066, N5067, N5068, N5069, N5070, N5071, N5072, N5073, N5076, N5080, N5081, N5082, N5085, N5088, N5092, N5093, N5094, N5097, N5101, N5102, N5103, N5106, N5109, N5113, N5114, N5115, N5118, N5121, N5124, N5127, N5130, N5134, N5135, N5136, N5139, N5142, N5146, N5147, N5148, N5151, N5155, N5156, N5157, N5160, N5163, N5167, N5168, N5169, N5172, N5176, N5180, N5184, N5188, N5192, N5193, N5194, N5197, N5200, N5204, N5205, N5206, N5209, N5213, N5214, N5215, N5218, N5221, N5225, N5226, N5227, N5230, N5234, N5235, N5236, N5239, N5240, N5241, N5244, N5245, N5246, N5249, N5250, N5251, N5254, N5255, N5256, N5259, N5262, N5266, N5267, N5268, N5271, N5275, N5276, N5277, N5280, N5283, N5287, N5288, N5289, N5292, N5296, N5297, N5298, N5301, N5304, N5309, N5312, N5315, N5318, N5322, N5323, N5324, N5327, N5331, N5332, N5333, N5336, N5339, N5343, N5344, N5345, N5348, N5352, N5353, N5354, N5357, N5360, N5364, N5365, N5366, N5370, N5374, N5378, N5379, N5380, N5383, N5387, N5388, N5389, N5392, N5395, N5399, N5400, N5401, N5404, N5408, N5409, N5410, N5413, N5416, N5420, N5421, N5422, N5425, N5426, N5427, N5428, N5429, N5430, N5431, N5434, N5438, N5439, N5440, N5443, N5446, N5450, N5451, N5452, N5455, N5459, N5460, N5461, N5464, N5467, N5471, N5472, N5473, N5476, N5480, N5483, N5486, N5489, N5493, N5494, N5495, N5498, N5501, N5505, N5506, N5507, N5510, N5514, N5515, N5516, N5519, N5522, N5526, N5527, N5528, N5531, N5535, N5536, N5537, N5540, N5544, N5548, N5552, N5553, N5554, N5557, N5560, N5564, N5565, N5566, N5569, N5573, N5574, N5575, N5578, N5581, N5585, N5586, N5587, N5590, N5594, N5595, N5596, N5599, N5602, N5606, N5607, N5608, N5611, N5612, N5613, N5616, N5617, N5618, N5621, N5624, N5628, N5629, N5630, N5633, N5637, N5638, N5639, N5642, N5645, N5649, N5650, N5651, N5654, N5658, N5659, N5660, N5663, N5666, N5670, N5671, N5673, N5676, N5679, N5683, N5684, N5685, N5688, N5692, N5693, N5694, N5697, N5700, N5704, N5705, N5706, N5709, N5713, N5714, N5715, N5718, N5721, N5725, N5726, N5727, N5730, N5734, N5738, N5739, N5740, N5743, N5747, N5748, N5749, N5752, N5755, N5759, N5760, N5761, N5764, N5768, N5769, N5770, N5773, N5776, N5780, N5781, N5782, N5785, N5786, N5787, N5788, N5789, N5792, N5796, N5797, N5798, N5801, N5804, N5808, N5809, N5810, N5813, N5817, N5818, N5819, N5822, N5825, N5829, N5830, N5831, N5834, N5837, N5840, N5844, N5845, N5846, N5849, N5852, N5856, N5857, N5858, N5861, N5865, N5866, N5867, N5870, N5873, N5877, N5878, N5879, N5882, N5886, N5890, N5891, N5892, N5895, N5898, N5902, N5903, N5904, N5907, N5911, N5912, N5913, N5916, N5919, N5923, N5924, N5925, N5928, N5929, N5930, N5933, N5934, N5935, N5938, N5941, N5945, N5946, N5947, N5950, N5954, N5955, N5956, N5959, N5962, N5966, N5967, N5968, N5972, N5975, N5979, N5980, N5981, N5984, N5988, N5989, N5990, N5993, N5996, N6000, N6001, N6002, N6005, N6009, N6010, N6011, N6014, N6018, N6019, N6020, N6023, N6026, N6030, N6031, N6032, N6035, N6036, N6037, N6040, N6044, N6045, N6046, N6049, N6052, N6056, N6057, N6058, N6061, N6064, N6068, N6069, N6070, N6073, N6076, N6080, N6081, N6082, N6085, N6089, N6090, N6091, N6094, N6097, N6101, N6102, N6103, N6106, N6107, N6108, N6111, N6114, N6118, N6119, N6120, N6124, N6128, N6129, N6130, N6133, N6134, N6135, N6138, N6141, N6145, N6146, N6147, N6151, N6155, N6156, N6157, N6161, N6165, N6166, N6167, N6171, N6175, N6176, N6177, N6181, N6185, N6186, N6187, N6191, N6195, N6196, N6197, N6201, N6205, N6206, N6207, N6211, N6215, N6216, N6217, N6221, N6225, N6226, N6227, N6231, N6235, N6236, N6237, N6241, N6245, N6246, N6247, N6251, N6255, N6256, N6257, N6261, N6265, N6266, N6267, N6271, N6275, N6276, N6277, N6281, N6285, N6286;


wire Trigger_en65_0,  troj65_0n1,  troj65_0n2,  troj65_0n3,  troj65_0n4,  troj65_0n5,  troj65_0n6,  troj65_0n7,  troj65_0n8,  tempN6265;

and2s1 U1 (.Q(N545), .DIN1(N1), .DIN2(N273));
and2s1 U2 (.Q(N546), .DIN1(N1), .DIN2(N290));
and2s1 U3 (.Q(N549), .DIN1(N1), .DIN2(N307));
and2s1 U4 (.Q(N552), .DIN1(N1), .DIN2(N324));
and2s1 U5 (.Q(N555), .DIN1(N1), .DIN2(N341));
and2s1 U6 (.Q(N558), .DIN1(N1), .DIN2(N358));
and2s1 U7 (.Q(N561), .DIN1(N1), .DIN2(N375));
and2s1 U8 (.Q(N564), .DIN1(N1), .DIN2(N392));
and2s1 U9 (.Q(N567), .DIN1(N1), .DIN2(N409));
and2s1 U10 (.Q(N570), .DIN1(N1), .DIN2(N426));
and2s1 U11 (.Q(N573), .DIN1(N1), .DIN2(N443));
and2s1 U12 (.Q(N576), .DIN1(N1), .DIN2(N460));
and2s1 U13 (.Q(N579), .DIN1(N1), .DIN2(N477));
and2s1 U14 (.Q(N582), .DIN1(N1), .DIN2(N494));
and2s1 U15 (.Q(N585), .DIN1(N1), .DIN2(N511));
and2s1 U16 (.Q(N588), .DIN1(N1), .DIN2(N528));
and2s1 U17 (.Q(N591), .DIN1(N18), .DIN2(N273));
and2s1 U18 (.Q(N594), .DIN1(N18), .DIN2(N290));
and2s1 U19 (.Q(N597), .DIN1(N18), .DIN2(N307));
and2s1 U20 (.Q(N600), .DIN1(N18), .DIN2(N324));
and2s1 U21 (.Q(N603), .DIN1(N18), .DIN2(N341));
and2s1 U22 (.Q(N606), .DIN1(N18), .DIN2(N358));
and2s1 U23 (.Q(N609), .DIN1(N18), .DIN2(N375));
and2s1 U24 (.Q(N612), .DIN1(N18), .DIN2(N392));
and2s1 U25 (.Q(N615), .DIN1(N18), .DIN2(N409));
and2s1 U26 (.Q(N618), .DIN1(N18), .DIN2(N426));
and2s1 U27 (.Q(N621), .DIN1(N18), .DIN2(N443));
and2s1 U28 (.Q(N624), .DIN1(N18), .DIN2(N460));
and2s1 U29 (.Q(N627), .DIN1(N18), .DIN2(N477));
and2s1 U30 (.Q(N630), .DIN1(N18), .DIN2(N494));
and2s1 U31 (.Q(N633), .DIN1(N18), .DIN2(N511));
and2s1 U32 (.Q(N636), .DIN1(N18), .DIN2(N528));
and2s1 U33 (.Q(N639), .DIN1(N35), .DIN2(N273));
and2s1 U34 (.Q(N642), .DIN1(N35), .DIN2(N290));
and2s1 U35 (.Q(N645), .DIN1(N35), .DIN2(N307));
and2s1 U36 (.Q(N648), .DIN1(N35), .DIN2(N324));
and2s1 U37 (.Q(N651), .DIN1(N35), .DIN2(N341));
and2s1 U38 (.Q(N654), .DIN1(N35), .DIN2(N358));
and2s1 U39 (.Q(N657), .DIN1(N35), .DIN2(N375));
and2s1 U40 (.Q(N660), .DIN1(N35), .DIN2(N392));
and2s1 U41 (.Q(N663), .DIN1(N35), .DIN2(N409));
and2s1 U42 (.Q(N666), .DIN1(N35), .DIN2(N426));
and2s1 U43 (.Q(N669), .DIN1(N35), .DIN2(N443));
and2s1 U44 (.Q(N672), .DIN1(N35), .DIN2(N460));
and2s1 U45 (.Q(N675), .DIN1(N35), .DIN2(N477));
and2s1 U46 (.Q(N678), .DIN1(N35), .DIN2(N494));
and2s1 U47 (.Q(N681), .DIN1(N35), .DIN2(N511));
and2s1 U48 (.Q(N684), .DIN1(N35), .DIN2(N528));
and2s1 U49 (.Q(N687), .DIN1(N52), .DIN2(N273));
and2s1 U50 (.Q(N690), .DIN1(N52), .DIN2(N290));
and2s1 U51 (.Q(N693), .DIN1(N52), .DIN2(N307));
and2s1 U52 (.Q(N696), .DIN1(N52), .DIN2(N324));
and2s1 U53 (.Q(N699), .DIN1(N52), .DIN2(N341));
and2s1 U54 (.Q(N702), .DIN1(N52), .DIN2(N358));
and2s1 U55 (.Q(N705), .DIN1(N52), .DIN2(N375));
and2s1 U56 (.Q(N708), .DIN1(N52), .DIN2(N392));
and2s1 U57 (.Q(N711), .DIN1(N52), .DIN2(N409));
and2s1 U58 (.Q(N714), .DIN1(N52), .DIN2(N426));
and2s1 U59 (.Q(N717), .DIN1(N52), .DIN2(N443));
and2s1 U60 (.Q(N720), .DIN1(N52), .DIN2(N460));
and2s1 U61 (.Q(N723), .DIN1(N52), .DIN2(N477));
and2s1 U62 (.Q(N726), .DIN1(N52), .DIN2(N494));
and2s1 U63 (.Q(N729), .DIN1(N52), .DIN2(N511));
and2s1 U64 (.Q(N732), .DIN1(N52), .DIN2(N528));
and2s1 U65 (.Q(N735), .DIN1(N69), .DIN2(N273));
and2s1 U66 (.Q(N738), .DIN1(N69), .DIN2(N290));
and2s1 U67 (.Q(N741), .DIN1(N69), .DIN2(N307));
and2s1 U68 (.Q(N744), .DIN1(N69), .DIN2(N324));
and2s1 U69 (.Q(N747), .DIN1(N69), .DIN2(N341));
and2s1 U70 (.Q(N750), .DIN1(N69), .DIN2(N358));
and2s1 U71 (.Q(N753), .DIN1(N69), .DIN2(N375));
and2s1 U72 (.Q(N756), .DIN1(N69), .DIN2(N392));
and2s1 U73 (.Q(N759), .DIN1(N69), .DIN2(N409));
and2s1 U74 (.Q(N762), .DIN1(N69), .DIN2(N426));
and2s1 U75 (.Q(N765), .DIN1(N69), .DIN2(N443));
and2s1 U76 (.Q(N768), .DIN1(N69), .DIN2(N460));
and2s1 U77 (.Q(N771), .DIN1(N69), .DIN2(N477));
and2s1 U78 (.Q(N774), .DIN1(N69), .DIN2(N494));
and2s1 U79 (.Q(N777), .DIN1(N69), .DIN2(N511));
and2s1 U80 (.Q(N780), .DIN1(N69), .DIN2(N528));
and2s1 U81 (.Q(N783), .DIN1(N86), .DIN2(N273));
and2s1 U82 (.Q(N786), .DIN1(N86), .DIN2(N290));
and2s1 U83 (.Q(N789), .DIN1(N86), .DIN2(N307));
and2s1 U84 (.Q(N792), .DIN1(N86), .DIN2(N324));
and2s1 U85 (.Q(N795), .DIN1(N86), .DIN2(N341));
and2s1 U86 (.Q(N798), .DIN1(N86), .DIN2(N358));
and2s1 U87 (.Q(N801), .DIN1(N86), .DIN2(N375));
and2s1 U88 (.Q(N804), .DIN1(N86), .DIN2(N392));
and2s1 U89 (.Q(N807), .DIN1(N86), .DIN2(N409));
and2s1 U90 (.Q(N810), .DIN1(N86), .DIN2(N426));
and2s1 U91 (.Q(N813), .DIN1(N86), .DIN2(N443));
and2s1 U92 (.Q(N816), .DIN1(N86), .DIN2(N460));
and2s1 U93 (.Q(N819), .DIN1(N86), .DIN2(N477));
and2s1 U94 (.Q(N822), .DIN1(N86), .DIN2(N494));
and2s1 U95 (.Q(N825), .DIN1(N86), .DIN2(N511));
and2s1 U96 (.Q(N828), .DIN1(N86), .DIN2(N528));
and2s1 U97 (.Q(N831), .DIN1(N103), .DIN2(N273));
and2s1 U98 (.Q(N834), .DIN1(N103), .DIN2(N290));
and2s1 U99 (.Q(N837), .DIN1(N103), .DIN2(N307));
and2s1 U100 (.Q(N840), .DIN1(N103), .DIN2(N324));
and2s1 U101 (.Q(N843), .DIN1(N103), .DIN2(N341));
and2s1 U102 (.Q(N846), .DIN1(N103), .DIN2(N358));
and2s1 U103 (.Q(N849), .DIN1(N103), .DIN2(N375));
and2s1 U104 (.Q(N852), .DIN1(N103), .DIN2(N392));
and2s1 U105 (.Q(N855), .DIN1(N103), .DIN2(N409));
and2s1 U106 (.Q(N858), .DIN1(N103), .DIN2(N426));
and2s1 U107 (.Q(N861), .DIN1(N103), .DIN2(N443));
and2s1 U108 (.Q(N864), .DIN1(N103), .DIN2(N460));
and2s1 U109 (.Q(N867), .DIN1(N103), .DIN2(N477));
and2s1 U110 (.Q(N870), .DIN1(N103), .DIN2(N494));
and2s1 U111 (.Q(N873), .DIN1(N103), .DIN2(N511));
and2s1 U112 (.Q(N876), .DIN1(N103), .DIN2(N528));
and2s1 U113 (.Q(N879), .DIN1(N120), .DIN2(N273));
and2s1 U114 (.Q(N882), .DIN1(N120), .DIN2(N290));
and2s1 U115 (.Q(N885), .DIN1(N120), .DIN2(N307));
and2s1 U116 (.Q(N888), .DIN1(N120), .DIN2(N324));
and2s1 U117 (.Q(N891), .DIN1(N120), .DIN2(N341));
and2s1 U118 (.Q(N894), .DIN1(N120), .DIN2(N358));
and2s1 U119 (.Q(N897), .DIN1(N120), .DIN2(N375));
and2s1 U120 (.Q(N900), .DIN1(N120), .DIN2(N392));
and2s1 U121 (.Q(N903), .DIN1(N120), .DIN2(N409));
and2s1 U122 (.Q(N906), .DIN1(N120), .DIN2(N426));
and2s1 U123 (.Q(N909), .DIN1(N120), .DIN2(N443));
and2s1 U124 (.Q(N912), .DIN1(N120), .DIN2(N460));
and2s1 U125 (.Q(N915), .DIN1(N120), .DIN2(N477));
and2s1 U126 (.Q(N918), .DIN1(N120), .DIN2(N494));
and2s1 U127 (.Q(N921), .DIN1(N120), .DIN2(N511));
and2s1 U128 (.Q(N924), .DIN1(N120), .DIN2(N528));
and2s1 U129 (.Q(N927), .DIN1(N137), .DIN2(N273));
and2s1 U130 (.Q(N930), .DIN1(N137), .DIN2(N290));
and2s1 U131 (.Q(N933), .DIN1(N137), .DIN2(N307));
and2s1 U132 (.Q(N936), .DIN1(N137), .DIN2(N324));
and2s1 U133 (.Q(N939), .DIN1(N137), .DIN2(N341));
and2s1 U134 (.Q(N942), .DIN1(N137), .DIN2(N358));
and2s1 U135 (.Q(N945), .DIN1(N137), .DIN2(N375));
and2s1 U136 (.Q(N948), .DIN1(N137), .DIN2(N392));
and2s1 U137 (.Q(N951), .DIN1(N137), .DIN2(N409));
and2s1 U138 (.Q(N954), .DIN1(N137), .DIN2(N426));
and2s1 U139 (.Q(N957), .DIN1(N137), .DIN2(N443));
and2s1 U140 (.Q(N960), .DIN1(N137), .DIN2(N460));
and2s1 U141 (.Q(N963), .DIN1(N137), .DIN2(N477));
and2s1 U142 (.Q(N966), .DIN1(N137), .DIN2(N494));
and2s1 U143 (.Q(N969), .DIN1(N137), .DIN2(N511));
and2s1 U144 (.Q(N972), .DIN1(N137), .DIN2(N528));
and2s1 U145 (.Q(N975), .DIN1(N154), .DIN2(N273));
and2s1 U146 (.Q(N978), .DIN1(N154), .DIN2(N290));
and2s1 U147 (.Q(N981), .DIN1(N154), .DIN2(N307));
and2s1 U148 (.Q(N984), .DIN1(N154), .DIN2(N324));
and2s1 U149 (.Q(N987), .DIN1(N154), .DIN2(N341));
and2s1 U150 (.Q(N990), .DIN1(N154), .DIN2(N358));
and2s1 U151 (.Q(N993), .DIN1(N154), .DIN2(N375));
and2s1 U152 (.Q(N996), .DIN1(N154), .DIN2(N392));
and2s1 U153 (.Q(N999), .DIN1(N154), .DIN2(N409));
and2s1 U154 (.Q(N1002), .DIN1(N154), .DIN2(N426));
and2s1 U155 (.Q(N1005), .DIN1(N154), .DIN2(N443));
and2s1 U156 (.Q(N1008), .DIN1(N154), .DIN2(N460));
and2s1 U157 (.Q(N1011), .DIN1(N154), .DIN2(N477));
and2s1 U158 (.Q(N1014), .DIN1(N154), .DIN2(N494));
and2s1 U159 (.Q(N1017), .DIN1(N154), .DIN2(N511));
and2s1 U160 (.Q(N1020), .DIN1(N154), .DIN2(N528));
and2s1 U161 (.Q(N1023), .DIN1(N171), .DIN2(N273));
and2s1 U162 (.Q(N1026), .DIN1(N171), .DIN2(N290));
and2s1 U163 (.Q(N1029), .DIN1(N171), .DIN2(N307));
and2s1 U164 (.Q(N1032), .DIN1(N171), .DIN2(N324));
and2s1 U165 (.Q(N1035), .DIN1(N171), .DIN2(N341));
and2s1 U166 (.Q(N1038), .DIN1(N171), .DIN2(N358));
and2s1 U167 (.Q(N1041), .DIN1(N171), .DIN2(N375));
and2s1 U168 (.Q(N1044), .DIN1(N171), .DIN2(N392));
and2s1 U169 (.Q(N1047), .DIN1(N171), .DIN2(N409));
and2s1 U170 (.Q(N1050), .DIN1(N171), .DIN2(N426));
and2s1 U171 (.Q(N1053), .DIN1(N171), .DIN2(N443));
and2s1 U172 (.Q(N1056), .DIN1(N171), .DIN2(N460));
and2s1 U173 (.Q(N1059), .DIN1(N171), .DIN2(N477));
and2s1 U174 (.Q(N1062), .DIN1(N171), .DIN2(N494));
and2s1 U175 (.Q(N1065), .DIN1(N171), .DIN2(N511));
and2s1 U176 (.Q(N1068), .DIN1(N171), .DIN2(N528));
and2s1 U177 (.Q(N1071), .DIN1(N188), .DIN2(N273));
and2s1 U178 (.Q(N1074), .DIN1(N188), .DIN2(N290));
and2s1 U179 (.Q(N1077), .DIN1(N188), .DIN2(N307));
and2s1 U180 (.Q(N1080), .DIN1(N188), .DIN2(N324));
and2s1 U181 (.Q(N1083), .DIN1(N188), .DIN2(N341));
and2s1 U182 (.Q(N1086), .DIN1(N188), .DIN2(N358));
and2s1 U183 (.Q(N1089), .DIN1(N188), .DIN2(N375));
and2s1 U184 (.Q(N1092), .DIN1(N188), .DIN2(N392));
and2s1 U185 (.Q(N1095), .DIN1(N188), .DIN2(N409));
and2s1 U186 (.Q(N1098), .DIN1(N188), .DIN2(N426));
and2s1 U187 (.Q(N1101), .DIN1(N188), .DIN2(N443));
and2s1 U188 (.Q(N1104), .DIN1(N188), .DIN2(N460));
and2s1 U189 (.Q(N1107), .DIN1(N188), .DIN2(N477));
and2s1 U190 (.Q(N1110), .DIN1(N188), .DIN2(N494));
and2s1 U191 (.Q(N1113), .DIN1(N188), .DIN2(N511));
and2s1 U192 (.Q(N1116), .DIN1(N188), .DIN2(N528));
and2s1 U193 (.Q(N1119), .DIN1(N205), .DIN2(N273));
and2s1 U194 (.Q(N1122), .DIN1(N205), .DIN2(N290));
and2s1 U195 (.Q(N1125), .DIN1(N205), .DIN2(N307));
and2s1 U196 (.Q(N1128), .DIN1(N205), .DIN2(N324));
and2s1 U197 (.Q(N1131), .DIN1(N205), .DIN2(N341));
and2s1 U198 (.Q(N1134), .DIN1(N205), .DIN2(N358));
and2s1 U199 (.Q(N1137), .DIN1(N205), .DIN2(N375));
and2s1 U200 (.Q(N1140), .DIN1(N205), .DIN2(N392));
and2s1 U201 (.Q(N1143), .DIN1(N205), .DIN2(N409));
and2s1 U202 (.Q(N1146), .DIN1(N205), .DIN2(N426));
and2s1 U203 (.Q(N1149), .DIN1(N205), .DIN2(N443));
and2s1 U204 (.Q(N1152), .DIN1(N205), .DIN2(N460));
and2s1 U205 (.Q(N1155), .DIN1(N205), .DIN2(N477));
and2s1 U206 (.Q(N1158), .DIN1(N205), .DIN2(N494));
and2s1 U207 (.Q(N1161), .DIN1(N205), .DIN2(N511));
and2s1 U208 (.Q(N1164), .DIN1(N205), .DIN2(N528));
and2s1 U209 (.Q(N1167), .DIN1(N222), .DIN2(N273));
and2s1 U210 (.Q(N1170), .DIN1(N222), .DIN2(N290));
and2s1 U211 (.Q(N1173), .DIN1(N222), .DIN2(N307));
and2s1 U212 (.Q(N1176), .DIN1(N222), .DIN2(N324));
and2s1 U213 (.Q(N1179), .DIN1(N222), .DIN2(N341));
and2s1 U214 (.Q(N1182), .DIN1(N222), .DIN2(N358));
and2s1 U215 (.Q(N1185), .DIN1(N222), .DIN2(N375));
and2s1 U216 (.Q(N1188), .DIN1(N222), .DIN2(N392));
and2s1 U217 (.Q(N1191), .DIN1(N222), .DIN2(N409));
and2s1 U218 (.Q(N1194), .DIN1(N222), .DIN2(N426));
and2s1 U219 (.Q(N1197), .DIN1(N222), .DIN2(N443));
and2s1 U220 (.Q(N1200), .DIN1(N222), .DIN2(N460));
and2s1 U221 (.Q(N1203), .DIN1(N222), .DIN2(N477));
and2s1 U222 (.Q(N1206), .DIN1(N222), .DIN2(N494));
and2s1 U223 (.Q(N1209), .DIN1(N222), .DIN2(N511));
and2s1 U224 (.Q(N1212), .DIN1(N222), .DIN2(N528));
and2s1 U225 (.Q(N1215), .DIN1(N239), .DIN2(N273));
and2s1 U226 (.Q(N1218), .DIN1(N239), .DIN2(N290));
and2s1 U227 (.Q(N1221), .DIN1(N239), .DIN2(N307));
and2s1 U228 (.Q(N1224), .DIN1(N239), .DIN2(N324));
and2s1 U229 (.Q(N1227), .DIN1(N239), .DIN2(N341));
and2s1 U230 (.Q(N1230), .DIN1(N239), .DIN2(N358));
and2s1 U231 (.Q(N1233), .DIN1(N239), .DIN2(N375));
and2s1 U232 (.Q(N1236), .DIN1(N239), .DIN2(N392));
and2s1 U233 (.Q(N1239), .DIN1(N239), .DIN2(N409));
and2s1 U234 (.Q(N1242), .DIN1(N239), .DIN2(N426));
and2s1 U235 (.Q(N1245), .DIN1(N239), .DIN2(N443));
and2s1 U236 (.Q(N1248), .DIN1(N239), .DIN2(N460));
and2s1 U237 (.Q(N1251), .DIN1(N239), .DIN2(N477));
and2s1 U238 (.Q(N1254), .DIN1(N239), .DIN2(N494));
and2s1 U239 (.Q(N1257), .DIN1(N239), .DIN2(N511));
and2s1 U240 (.Q(N1260), .DIN1(N239), .DIN2(N528));
and2s1 U241 (.Q(N1263), .DIN1(N256), .DIN2(N273));
and2s1 U242 (.Q(N1266), .DIN1(N256), .DIN2(N290));
and2s1 U243 (.Q(N1269), .DIN1(N256), .DIN2(N307));
and2s1 U244 (.Q(N1272), .DIN1(N256), .DIN2(N324));
and2s1 U245 (.Q(N1275), .DIN1(N256), .DIN2(N341));
and2s1 U246 (.Q(N1278), .DIN1(N256), .DIN2(N358));
and2s1 U247 (.Q(N1281), .DIN1(N256), .DIN2(N375));
and2s1 U248 (.Q(N1284), .DIN1(N256), .DIN2(N392));
and2s1 U249 (.Q(N1287), .DIN1(N256), .DIN2(N409));
and2s1 U250 (.Q(N1290), .DIN1(N256), .DIN2(N426));
and2s1 U251 (.Q(N1293), .DIN1(N256), .DIN2(N443));
and2s1 U252 (.Q(N1296), .DIN1(N256), .DIN2(N460));
and2s1 U253 (.Q(N1299), .DIN1(N256), .DIN2(N477));
and2s1 U254 (.Q(N1302), .DIN1(N256), .DIN2(N494));
and2s1 U255 (.Q(N1305), .DIN1(N256), .DIN2(N511));
and2s1 U256 (.Q(N1308), .DIN1(N256), .DIN2(N528));
hi1s1 U257 (.Q(N1311), .DIN(N591));
hi1s1 U258 (.Q(N1315), .DIN(N639));
hi1s1 U259 (.Q(N1319), .DIN(N687));
hi1s1 U260 (.Q(N1323), .DIN(N735));
hi1s1 U261 (.Q(N1327), .DIN(N783));
hi1s1 U262 (.Q(N1331), .DIN(N831));
hi1s1 U263 (.Q(N1335), .DIN(N879));
hi1s1 U264 (.Q(N1339), .DIN(N927));
hi1s1 U265 (.Q(N1343), .DIN(N975));
hi1s1 U266 (.Q(N1347), .DIN(N1023));
hi1s1 U267 (.Q(N1351), .DIN(N1071));
hi1s1 U268 (.Q(N1355), .DIN(N1119));
hi1s1 U269 (.Q(N1359), .DIN(N1167));
hi1s1 U270 (.Q(N1363), .DIN(N1215));
hi1s1 U271 (.Q(N1367), .DIN(N1263));
nor2s1 U272 (.Q(N1371), .DIN1(N591), .DIN2(N1311));
hi1s1 U273 (.Q(N1372), .DIN(N1311));
nor2s1 U274 (.Q(N1373), .DIN1(N639), .DIN2(N1315));
hi1s1 U275 (.Q(N1374), .DIN(N1315));
nor2s1 U276 (.Q(N1375), .DIN1(N687), .DIN2(N1319));
hi1s1 U277 (.Q(N1376), .DIN(N1319));
nor2s1 U278 (.Q(N1377), .DIN1(N735), .DIN2(N1323));
hi1s1 U279 (.Q(N1378), .DIN(N1323));
nor2s1 U280 (.Q(N1379), .DIN1(N783), .DIN2(N1327));
hi1s1 U281 (.Q(N1380), .DIN(N1327));
nor2s1 U282 (.Q(N1381), .DIN1(N831), .DIN2(N1331));
hi1s1 U283 (.Q(N1382), .DIN(N1331));
nor2s1 U284 (.Q(N1383), .DIN1(N879), .DIN2(N1335));
hi1s1 U285 (.Q(N1384), .DIN(N1335));
nor2s1 U286 (.Q(N1385), .DIN1(N927), .DIN2(N1339));
hi1s1 U287 (.Q(N1386), .DIN(N1339));
nor2s1 U288 (.Q(N1387), .DIN1(N975), .DIN2(N1343));
hi1s1 U289 (.Q(N1388), .DIN(N1343));
nor2s1 U290 (.Q(N1389), .DIN1(N1023), .DIN2(N1347));
hi1s1 U291 (.Q(N1390), .DIN(N1347));
nor2s1 U292 (.Q(N1391), .DIN1(N1071), .DIN2(N1351));
hi1s1 U293 (.Q(N1392), .DIN(N1351));
nor2s1 U294 (.Q(N1393), .DIN1(N1119), .DIN2(N1355));
hi1s1 U295 (.Q(N1394), .DIN(N1355));
nor2s1 U296 (.Q(N1395), .DIN1(N1167), .DIN2(N1359));
hi1s1 U297 (.Q(N1396), .DIN(N1359));
nor2s1 U298 (.Q(N1397), .DIN1(N1215), .DIN2(N1363));
hi1s1 U299 (.Q(N1398), .DIN(N1363));
nor2s1 U300 (.Q(N1399), .DIN1(N1263), .DIN2(N1367));
hi1s1 U301 (.Q(N1400), .DIN(N1367));
nor2s1 U302 (.Q(N1401), .DIN1(N1371), .DIN2(N1372));
nor2s1 U303 (.Q(N1404), .DIN1(N1373), .DIN2(N1374));
nor2s1 U304 (.Q(N1407), .DIN1(N1375), .DIN2(N1376));
nor2s1 U305 (.Q(N1410), .DIN1(N1377), .DIN2(N1378));
nor2s1 U306 (.Q(N1413), .DIN1(N1379), .DIN2(N1380));
nor2s1 U307 (.Q(N1416), .DIN1(N1381), .DIN2(N1382));
nor2s1 U308 (.Q(N1419), .DIN1(N1383), .DIN2(N1384));
nor2s1 U309 (.Q(N1422), .DIN1(N1385), .DIN2(N1386));
nor2s1 U310 (.Q(N1425), .DIN1(N1387), .DIN2(N1388));
nor2s1 U311 (.Q(N1428), .DIN1(N1389), .DIN2(N1390));
nor2s1 U312 (.Q(N1431), .DIN1(N1391), .DIN2(N1392));
nor2s1 U313 (.Q(N1434), .DIN1(N1393), .DIN2(N1394));
nor2s1 U314 (.Q(N1437), .DIN1(N1395), .DIN2(N1396));
nor2s1 U315 (.Q(N1440), .DIN1(N1397), .DIN2(N1398));
nor2s1 U316 (.Q(N1443), .DIN1(N1399), .DIN2(N1400));
nor2s1 U317 (.Q(N1446), .DIN1(N1401), .DIN2(N546));
nor2s1 U318 (.Q(N1450), .DIN1(N1404), .DIN2(N594));
nor2s1 U319 (.Q(N1454), .DIN1(N1407), .DIN2(N642));
nor2s1 U320 (.Q(N1458), .DIN1(N1410), .DIN2(N690));
nor2s1 U321 (.Q(N1462), .DIN1(N1413), .DIN2(N738));
nor2s1 U322 (.Q(N1466), .DIN1(N1416), .DIN2(N786));
nor2s1 U323 (.Q(N1470), .DIN1(N1419), .DIN2(N834));
nor2s1 U324 (.Q(N1474), .DIN1(N1422), .DIN2(N882));
nor2s1 U325 (.Q(N1478), .DIN1(N1425), .DIN2(N930));
nor2s1 U326 (.Q(N1482), .DIN1(N1428), .DIN2(N978));
nor2s1 U327 (.Q(N1486), .DIN1(N1431), .DIN2(N1026));
nor2s1 U328 (.Q(N1490), .DIN1(N1434), .DIN2(N1074));
nor2s1 U329 (.Q(N1494), .DIN1(N1437), .DIN2(N1122));
nor2s1 U330 (.Q(N1498), .DIN1(N1440), .DIN2(N1170));
nor2s1 U331 (.Q(N1502), .DIN1(N1443), .DIN2(N1218));
nor2s1 U332 (.Q(N1506), .DIN1(N1401), .DIN2(N1446));
nor2s1 U333 (.Q(N1507), .DIN1(N1446), .DIN2(N546));
nor2s1 U334 (.Q(N1508), .DIN1(N1311), .DIN2(N1446));
nor2s1 U335 (.Q(N1511), .DIN1(N1404), .DIN2(N1450));
nor2s1 U336 (.Q(N1512), .DIN1(N1450), .DIN2(N594));
nor2s1 U337 (.Q(N1513), .DIN1(N1315), .DIN2(N1450));
nor2s1 U338 (.Q(N1516), .DIN1(N1407), .DIN2(N1454));
nor2s1 U339 (.Q(N1517), .DIN1(N1454), .DIN2(N642));
nor2s1 U340 (.Q(N1518), .DIN1(N1319), .DIN2(N1454));
nor2s1 U341 (.Q(N1521), .DIN1(N1410), .DIN2(N1458));
nor2s1 U342 (.Q(N1522), .DIN1(N1458), .DIN2(N690));
nor2s1 U343 (.Q(N1523), .DIN1(N1323), .DIN2(N1458));
nor2s1 U344 (.Q(N1526), .DIN1(N1413), .DIN2(N1462));
nor2s1 U345 (.Q(N1527), .DIN1(N1462), .DIN2(N738));
nor2s1 U346 (.Q(N1528), .DIN1(N1327), .DIN2(N1462));
nor2s1 U347 (.Q(N1531), .DIN1(N1416), .DIN2(N1466));
nor2s1 U348 (.Q(N1532), .DIN1(N1466), .DIN2(N786));
nor2s1 U349 (.Q(N1533), .DIN1(N1331), .DIN2(N1466));
nor2s1 U350 (.Q(N1536), .DIN1(N1419), .DIN2(N1470));
nor2s1 U351 (.Q(N1537), .DIN1(N1470), .DIN2(N834));
nor2s1 U352 (.Q(N1538), .DIN1(N1335), .DIN2(N1470));
nor2s1 U353 (.Q(N1541), .DIN1(N1422), .DIN2(N1474));
nor2s1 U354 (.Q(N1542), .DIN1(N1474), .DIN2(N882));
nor2s1 U355 (.Q(N1543), .DIN1(N1339), .DIN2(N1474));
nor2s1 U356 (.Q(N1546), .DIN1(N1425), .DIN2(N1478));
nor2s1 U357 (.Q(N1547), .DIN1(N1478), .DIN2(N930));
nor2s1 U358 (.Q(N1548), .DIN1(N1343), .DIN2(N1478));
nor2s1 U359 (.Q(N1551), .DIN1(N1428), .DIN2(N1482));
nor2s1 U360 (.Q(N1552), .DIN1(N1482), .DIN2(N978));
nor2s1 U361 (.Q(N1553), .DIN1(N1347), .DIN2(N1482));
nor2s1 U362 (.Q(N1556), .DIN1(N1431), .DIN2(N1486));
nor2s1 U363 (.Q(N1557), .DIN1(N1486), .DIN2(N1026));
nor2s1 U364 (.Q(N1558), .DIN1(N1351), .DIN2(N1486));
nor2s1 U365 (.Q(N1561), .DIN1(N1434), .DIN2(N1490));
nor2s1 U366 (.Q(N1562), .DIN1(N1490), .DIN2(N1074));
nor2s1 U367 (.Q(N1563), .DIN1(N1355), .DIN2(N1490));
nor2s1 U368 (.Q(N1566), .DIN1(N1437), .DIN2(N1494));
nor2s1 U369 (.Q(N1567), .DIN1(N1494), .DIN2(N1122));
nor2s1 U370 (.Q(N1568), .DIN1(N1359), .DIN2(N1494));
nor2s1 U371 (.Q(N1571), .DIN1(N1440), .DIN2(N1498));
nor2s1 U372 (.Q(N1572), .DIN1(N1498), .DIN2(N1170));
nor2s1 U373 (.Q(N1573), .DIN1(N1363), .DIN2(N1498));
nor2s1 U374 (.Q(N1576), .DIN1(N1443), .DIN2(N1502));
nor2s1 U375 (.Q(N1577), .DIN1(N1502), .DIN2(N1218));
nor2s1 U376 (.Q(N1578), .DIN1(N1367), .DIN2(N1502));
nor2s1 U377 (.Q(N1581), .DIN1(N1506), .DIN2(N1507));
nor2s1 U378 (.Q(N1582), .DIN1(N1511), .DIN2(N1512));
nor2s1 U379 (.Q(N1585), .DIN1(N1516), .DIN2(N1517));
nor2s1 U380 (.Q(N1588), .DIN1(N1521), .DIN2(N1522));
nor2s1 U381 (.Q(N1591), .DIN1(N1526), .DIN2(N1527));
nor2s1 U382 (.Q(N1594), .DIN1(N1531), .DIN2(N1532));
nor2s1 U383 (.Q(N1597), .DIN1(N1536), .DIN2(N1537));
nor2s1 U384 (.Q(N1600), .DIN1(N1541), .DIN2(N1542));
nor2s1 U385 (.Q(N1603), .DIN1(N1546), .DIN2(N1547));
nor2s1 U386 (.Q(N1606), .DIN1(N1551), .DIN2(N1552));
nor2s1 U387 (.Q(N1609), .DIN1(N1556), .DIN2(N1557));
nor2s1 U388 (.Q(N1612), .DIN1(N1561), .DIN2(N1562));
nor2s1 U389 (.Q(N1615), .DIN1(N1566), .DIN2(N1567));
nor2s1 U390 (.Q(N1618), .DIN1(N1571), .DIN2(N1572));
nor2s1 U391 (.Q(N1621), .DIN1(N1576), .DIN2(N1577));
nor2s1 U392 (.Q(N1624), .DIN1(N1266), .DIN2(N1578));
nor2s1 U393 (.Q(N1628), .DIN1(N1582), .DIN2(N1508));
nor2s1 U394 (.Q(N1632), .DIN1(N1585), .DIN2(N1513));
nor2s1 U395 (.Q(N1636), .DIN1(N1588), .DIN2(N1518));
nor2s1 U396 (.Q(N1640), .DIN1(N1591), .DIN2(N1523));
nor2s1 U397 (.Q(N1644), .DIN1(N1594), .DIN2(N1528));
nor2s1 U398 (.Q(N1648), .DIN1(N1597), .DIN2(N1533));
nor2s1 U399 (.Q(N1652), .DIN1(N1600), .DIN2(N1538));
nor2s1 U400 (.Q(N1656), .DIN1(N1603), .DIN2(N1543));
nor2s1 U401 (.Q(N1660), .DIN1(N1606), .DIN2(N1548));
nor2s1 U402 (.Q(N1664), .DIN1(N1609), .DIN2(N1553));
nor2s1 U403 (.Q(N1668), .DIN1(N1612), .DIN2(N1558));
nor2s1 U404 (.Q(N1672), .DIN1(N1615), .DIN2(N1563));
nor2s1 U405 (.Q(N1676), .DIN1(N1618), .DIN2(N1568));
nor2s1 U406 (.Q(N1680), .DIN1(N1621), .DIN2(N1573));
nor2s1 U407 (.Q(N1684), .DIN1(N1266), .DIN2(N1624));
nor2s1 U408 (.Q(N1685), .DIN1(N1624), .DIN2(N1578));
nor2s1 U409 (.Q(N1686), .DIN1(N1582), .DIN2(N1628));
nor2s1 U410 (.Q(N1687), .DIN1(N1628), .DIN2(N1508));
nor2s1 U411 (.Q(N1688), .DIN1(N1585), .DIN2(N1632));
nor2s1 U412 (.Q(N1689), .DIN1(N1632), .DIN2(N1513));
nor2s1 U413 (.Q(N1690), .DIN1(N1588), .DIN2(N1636));
nor2s1 U414 (.Q(N1691), .DIN1(N1636), .DIN2(N1518));
nor2s1 U415 (.Q(N1692), .DIN1(N1591), .DIN2(N1640));
nor2s1 U416 (.Q(N1693), .DIN1(N1640), .DIN2(N1523));
nor2s1 U417 (.Q(N1694), .DIN1(N1594), .DIN2(N1644));
nor2s1 U418 (.Q(N1695), .DIN1(N1644), .DIN2(N1528));
nor2s1 U419 (.Q(N1696), .DIN1(N1597), .DIN2(N1648));
nor2s1 U420 (.Q(N1697), .DIN1(N1648), .DIN2(N1533));
nor2s1 U421 (.Q(N1698), .DIN1(N1600), .DIN2(N1652));
nor2s1 U422 (.Q(N1699), .DIN1(N1652), .DIN2(N1538));
nor2s1 U423 (.Q(N1700), .DIN1(N1603), .DIN2(N1656));
nor2s1 U424 (.Q(N1701), .DIN1(N1656), .DIN2(N1543));
nor2s1 U425 (.Q(N1702), .DIN1(N1606), .DIN2(N1660));
nor2s1 U426 (.Q(N1703), .DIN1(N1660), .DIN2(N1548));
nor2s1 U427 (.Q(N1704), .DIN1(N1609), .DIN2(N1664));
nor2s1 U428 (.Q(N1705), .DIN1(N1664), .DIN2(N1553));
nor2s1 U429 (.Q(N1706), .DIN1(N1612), .DIN2(N1668));
nor2s1 U430 (.Q(N1707), .DIN1(N1668), .DIN2(N1558));
nor2s1 U431 (.Q(N1708), .DIN1(N1615), .DIN2(N1672));
nor2s1 U432 (.Q(N1709), .DIN1(N1672), .DIN2(N1563));
nor2s1 U433 (.Q(N1710), .DIN1(N1618), .DIN2(N1676));
nor2s1 U434 (.Q(N1711), .DIN1(N1676), .DIN2(N1568));
nor2s1 U435 (.Q(N1712), .DIN1(N1621), .DIN2(N1680));
nor2s1 U436 (.Q(N1713), .DIN1(N1680), .DIN2(N1573));
nor2s1 U437 (.Q(N1714), .DIN1(N1684), .DIN2(N1685));
nor2s1 U438 (.Q(N1717), .DIN1(N1686), .DIN2(N1687));
nor2s1 U439 (.Q(N1720), .DIN1(N1688), .DIN2(N1689));
nor2s1 U440 (.Q(N1723), .DIN1(N1690), .DIN2(N1691));
nor2s1 U441 (.Q(N1726), .DIN1(N1692), .DIN2(N1693));
nor2s1 U442 (.Q(N1729), .DIN1(N1694), .DIN2(N1695));
nor2s1 U443 (.Q(N1732), .DIN1(N1696), .DIN2(N1697));
nor2s1 U444 (.Q(N1735), .DIN1(N1698), .DIN2(N1699));
nor2s1 U445 (.Q(N1738), .DIN1(N1700), .DIN2(N1701));
nor2s1 U446 (.Q(N1741), .DIN1(N1702), .DIN2(N1703));
nor2s1 U447 (.Q(N1744), .DIN1(N1704), .DIN2(N1705));
nor2s1 U448 (.Q(N1747), .DIN1(N1706), .DIN2(N1707));
nor2s1 U449 (.Q(N1750), .DIN1(N1708), .DIN2(N1709));
nor2s1 U450 (.Q(N1753), .DIN1(N1710), .DIN2(N1711));
nor2s1 U451 (.Q(N1756), .DIN1(N1712), .DIN2(N1713));
nor2s1 U452 (.Q(N1759), .DIN1(N1714), .DIN2(N1221));
nor2s1 U453 (.Q(N1763), .DIN1(N1717), .DIN2(N549));
nor2s1 U454 (.Q(N1767), .DIN1(N1720), .DIN2(N597));
nor2s1 U455 (.Q(N1771), .DIN1(N1723), .DIN2(N645));
nor2s1 U456 (.Q(N1775), .DIN1(N1726), .DIN2(N693));
nor2s1 U457 (.Q(N1779), .DIN1(N1729), .DIN2(N741));
nor2s1 U458 (.Q(N1783), .DIN1(N1732), .DIN2(N789));
nor2s1 U459 (.Q(N1787), .DIN1(N1735), .DIN2(N837));
nor2s1 U460 (.Q(N1791), .DIN1(N1738), .DIN2(N885));
nor2s1 U461 (.Q(N1795), .DIN1(N1741), .DIN2(N933));
nor2s1 U462 (.Q(N1799), .DIN1(N1744), .DIN2(N981));
nor2s1 U463 (.Q(N1803), .DIN1(N1747), .DIN2(N1029));
nor2s1 U464 (.Q(N1807), .DIN1(N1750), .DIN2(N1077));
nor2s1 U465 (.Q(N1811), .DIN1(N1753), .DIN2(N1125));
nor2s1 U466 (.Q(N1815), .DIN1(N1756), .DIN2(N1173));
nor2s1 U467 (.Q(N1819), .DIN1(N1714), .DIN2(N1759));
nor2s1 U468 (.Q(N1820), .DIN1(N1759), .DIN2(N1221));
nor2s1 U469 (.Q(N1821), .DIN1(N1624), .DIN2(N1759));
nor2s1 U470 (.Q(N1824), .DIN1(N1717), .DIN2(N1763));
nor2s1 U471 (.Q(N1825), .DIN1(N1763), .DIN2(N549));
nor2s1 U472 (.Q(N1826), .DIN1(N1628), .DIN2(N1763));
nor2s1 U473 (.Q(N1829), .DIN1(N1720), .DIN2(N1767));
nor2s1 U474 (.Q(N1830), .DIN1(N1767), .DIN2(N597));
nor2s1 U475 (.Q(N1831), .DIN1(N1632), .DIN2(N1767));
nor2s1 U476 (.Q(N1834), .DIN1(N1723), .DIN2(N1771));
nor2s1 U477 (.Q(N1835), .DIN1(N1771), .DIN2(N645));
nor2s1 U478 (.Q(N1836), .DIN1(N1636), .DIN2(N1771));
nor2s1 U479 (.Q(N1839), .DIN1(N1726), .DIN2(N1775));
nor2s1 U480 (.Q(N1840), .DIN1(N1775), .DIN2(N693));
nor2s1 U481 (.Q(N1841), .DIN1(N1640), .DIN2(N1775));
nor2s1 U482 (.Q(N1844), .DIN1(N1729), .DIN2(N1779));
nor2s1 U483 (.Q(N1845), .DIN1(N1779), .DIN2(N741));
nor2s1 U484 (.Q(N1846), .DIN1(N1644), .DIN2(N1779));
nor2s1 U485 (.Q(N1849), .DIN1(N1732), .DIN2(N1783));
nor2s1 U486 (.Q(N1850), .DIN1(N1783), .DIN2(N789));
nor2s1 U487 (.Q(N1851), .DIN1(N1648), .DIN2(N1783));
nor2s1 U488 (.Q(N1854), .DIN1(N1735), .DIN2(N1787));
nor2s1 U489 (.Q(N1855), .DIN1(N1787), .DIN2(N837));
nor2s1 U490 (.Q(N1856), .DIN1(N1652), .DIN2(N1787));
nor2s1 U491 (.Q(N1859), .DIN1(N1738), .DIN2(N1791));
nor2s1 U492 (.Q(N1860), .DIN1(N1791), .DIN2(N885));
nor2s1 U493 (.Q(N1861), .DIN1(N1656), .DIN2(N1791));
nor2s1 U494 (.Q(N1864), .DIN1(N1741), .DIN2(N1795));
nor2s1 U495 (.Q(N1865), .DIN1(N1795), .DIN2(N933));
nor2s1 U496 (.Q(N1866), .DIN1(N1660), .DIN2(N1795));
nor2s1 U497 (.Q(N1869), .DIN1(N1744), .DIN2(N1799));
nor2s1 U498 (.Q(N1870), .DIN1(N1799), .DIN2(N981));
nor2s1 U499 (.Q(N1871), .DIN1(N1664), .DIN2(N1799));
nor2s1 U500 (.Q(N1874), .DIN1(N1747), .DIN2(N1803));
nor2s1 U501 (.Q(N1875), .DIN1(N1803), .DIN2(N1029));
nor2s1 U502 (.Q(N1876), .DIN1(N1668), .DIN2(N1803));
nor2s1 U503 (.Q(N1879), .DIN1(N1750), .DIN2(N1807));
nor2s1 U504 (.Q(N1880), .DIN1(N1807), .DIN2(N1077));
nor2s1 U505 (.Q(N1881), .DIN1(N1672), .DIN2(N1807));
nor2s1 U506 (.Q(N1884), .DIN1(N1753), .DIN2(N1811));
nor2s1 U507 (.Q(N1885), .DIN1(N1811), .DIN2(N1125));
nor2s1 U508 (.Q(N1886), .DIN1(N1676), .DIN2(N1811));
nor2s1 U509 (.Q(N1889), .DIN1(N1756), .DIN2(N1815));
nor2s1 U510 (.Q(N1890), .DIN1(N1815), .DIN2(N1173));
nor2s1 U511 (.Q(N1891), .DIN1(N1680), .DIN2(N1815));
nor2s1 U512 (.Q(N1894), .DIN1(N1819), .DIN2(N1820));
nor2s1 U513 (.Q(N1897), .DIN1(N1269), .DIN2(N1821));
nor2s1 U514 (.Q(N1901), .DIN1(N1824), .DIN2(N1825));
nor2s1 U515 (.Q(N1902), .DIN1(N1829), .DIN2(N1830));
nor2s1 U516 (.Q(N1905), .DIN1(N1834), .DIN2(N1835));
nor2s1 U517 (.Q(N1908), .DIN1(N1839), .DIN2(N1840));
nor2s1 U518 (.Q(N1911), .DIN1(N1844), .DIN2(N1845));
nor2s1 U519 (.Q(N1914), .DIN1(N1849), .DIN2(N1850));
nor2s1 U520 (.Q(N1917), .DIN1(N1854), .DIN2(N1855));
nor2s1 U521 (.Q(N1920), .DIN1(N1859), .DIN2(N1860));
nor2s1 U522 (.Q(N1923), .DIN1(N1864), .DIN2(N1865));
nor2s1 U523 (.Q(N1926), .DIN1(N1869), .DIN2(N1870));
nor2s1 U524 (.Q(N1929), .DIN1(N1874), .DIN2(N1875));
nor2s1 U525 (.Q(N1932), .DIN1(N1879), .DIN2(N1880));
nor2s1 U526 (.Q(N1935), .DIN1(N1884), .DIN2(N1885));
nor2s1 U527 (.Q(N1938), .DIN1(N1889), .DIN2(N1890));
nor2s1 U528 (.Q(N1941), .DIN1(N1894), .DIN2(N1891));
nor2s1 U529 (.Q(N1945), .DIN1(N1269), .DIN2(N1897));
nor2s1 U530 (.Q(N1946), .DIN1(N1897), .DIN2(N1821));
nor2s1 U531 (.Q(N1947), .DIN1(N1902), .DIN2(N1826));
nor2s1 U532 (.Q(N1951), .DIN1(N1905), .DIN2(N1831));
nor2s1 U533 (.Q(N1955), .DIN1(N1908), .DIN2(N1836));
nor2s1 U534 (.Q(N1959), .DIN1(N1911), .DIN2(N1841));
nor2s1 U535 (.Q(N1963), .DIN1(N1914), .DIN2(N1846));
nor2s1 U536 (.Q(N1967), .DIN1(N1917), .DIN2(N1851));
nor2s1 U537 (.Q(N1971), .DIN1(N1920), .DIN2(N1856));
nor2s1 U538 (.Q(N1975), .DIN1(N1923), .DIN2(N1861));
nor2s1 U539 (.Q(N1979), .DIN1(N1926), .DIN2(N1866));
nor2s1 U540 (.Q(N1983), .DIN1(N1929), .DIN2(N1871));
nor2s1 U541 (.Q(N1987), .DIN1(N1932), .DIN2(N1876));
nor2s1 U542 (.Q(N1991), .DIN1(N1935), .DIN2(N1881));
nor2s1 U543 (.Q(N1995), .DIN1(N1938), .DIN2(N1886));
nor2s1 U544 (.Q(N1999), .DIN1(N1894), .DIN2(N1941));
nor2s1 U545 (.Q(N2000), .DIN1(N1941), .DIN2(N1891));
nor2s1 U546 (.Q(N2001), .DIN1(N1945), .DIN2(N1946));
nor2s1 U547 (.Q(N2004), .DIN1(N1902), .DIN2(N1947));
nor2s1 U548 (.Q(N2005), .DIN1(N1947), .DIN2(N1826));
nor2s1 U549 (.Q(N2006), .DIN1(N1905), .DIN2(N1951));
nor2s1 U550 (.Q(N2007), .DIN1(N1951), .DIN2(N1831));
nor2s1 U551 (.Q(N2008), .DIN1(N1908), .DIN2(N1955));
nor2s1 U552 (.Q(N2009), .DIN1(N1955), .DIN2(N1836));
nor2s1 U553 (.Q(N2010), .DIN1(N1911), .DIN2(N1959));
nor2s1 U554 (.Q(N2011), .DIN1(N1959), .DIN2(N1841));
nor2s1 U555 (.Q(N2012), .DIN1(N1914), .DIN2(N1963));
nor2s1 U556 (.Q(N2013), .DIN1(N1963), .DIN2(N1846));
nor2s1 U557 (.Q(N2014), .DIN1(N1917), .DIN2(N1967));
nor2s1 U558 (.Q(N2015), .DIN1(N1967), .DIN2(N1851));
nor2s1 U559 (.Q(N2016), .DIN1(N1920), .DIN2(N1971));
nor2s1 U560 (.Q(N2017), .DIN1(N1971), .DIN2(N1856));
nor2s1 U561 (.Q(N2018), .DIN1(N1923), .DIN2(N1975));
nor2s1 U562 (.Q(N2019), .DIN1(N1975), .DIN2(N1861));
nor2s1 U563 (.Q(N2020), .DIN1(N1926), .DIN2(N1979));
nor2s1 U564 (.Q(N2021), .DIN1(N1979), .DIN2(N1866));
nor2s1 U565 (.Q(N2022), .DIN1(N1929), .DIN2(N1983));
nor2s1 U566 (.Q(N2023), .DIN1(N1983), .DIN2(N1871));
nor2s1 U567 (.Q(N2024), .DIN1(N1932), .DIN2(N1987));
nor2s1 U568 (.Q(N2025), .DIN1(N1987), .DIN2(N1876));
nor2s1 U569 (.Q(N2026), .DIN1(N1935), .DIN2(N1991));
nor2s1 U570 (.Q(N2027), .DIN1(N1991), .DIN2(N1881));
nor2s1 U571 (.Q(N2028), .DIN1(N1938), .DIN2(N1995));
nor2s1 U572 (.Q(N2029), .DIN1(N1995), .DIN2(N1886));
nor2s1 U573 (.Q(N2030), .DIN1(N1999), .DIN2(N2000));
nor2s1 U574 (.Q(N2033), .DIN1(N2001), .DIN2(N1224));
nor2s1 U575 (.Q(N2037), .DIN1(N2004), .DIN2(N2005));
nor2s1 U576 (.Q(N2040), .DIN1(N2006), .DIN2(N2007));
nor2s1 U577 (.Q(N2043), .DIN1(N2008), .DIN2(N2009));
nor2s1 U578 (.Q(N2046), .DIN1(N2010), .DIN2(N2011));
nor2s1 U579 (.Q(N2049), .DIN1(N2012), .DIN2(N2013));
nor2s1 U580 (.Q(N2052), .DIN1(N2014), .DIN2(N2015));
nor2s1 U581 (.Q(N2055), .DIN1(N2016), .DIN2(N2017));
nor2s1 U582 (.Q(N2058), .DIN1(N2018), .DIN2(N2019));
nor2s1 U583 (.Q(N2061), .DIN1(N2020), .DIN2(N2021));
nor2s1 U584 (.Q(N2064), .DIN1(N2022), .DIN2(N2023));
nor2s1 U585 (.Q(N2067), .DIN1(N2024), .DIN2(N2025));
nor2s1 U586 (.Q(N2070), .DIN1(N2026), .DIN2(N2027));
nor2s1 U587 (.Q(N2073), .DIN1(N2028), .DIN2(N2029));
nor2s1 U588 (.Q(N2076), .DIN1(N2030), .DIN2(N1176));
nor2s1 U589 (.Q(N2080), .DIN1(N2001), .DIN2(N2033));
nor2s1 U590 (.Q(N2081), .DIN1(N2033), .DIN2(N1224));
nor2s1 U591 (.Q(N2082), .DIN1(N1897), .DIN2(N2033));
nor2s1 U592 (.Q(N2085), .DIN1(N2037), .DIN2(N552));
nor2s1 U593 (.Q(N2089), .DIN1(N2040), .DIN2(N600));
nor2s1 U594 (.Q(N2093), .DIN1(N2043), .DIN2(N648));
nor2s1 U595 (.Q(N2097), .DIN1(N2046), .DIN2(N696));
nor2s1 U596 (.Q(N2101), .DIN1(N2049), .DIN2(N744));
nor2s1 U597 (.Q(N2105), .DIN1(N2052), .DIN2(N792));
nor2s1 U598 (.Q(N2109), .DIN1(N2055), .DIN2(N840));
nor2s1 U599 (.Q(N2113), .DIN1(N2058), .DIN2(N888));
nor2s1 U600 (.Q(N2117), .DIN1(N2061), .DIN2(N936));
nor2s1 U601 (.Q(N2121), .DIN1(N2064), .DIN2(N984));
nor2s1 U602 (.Q(N2125), .DIN1(N2067), .DIN2(N1032));
nor2s1 U603 (.Q(N2129), .DIN1(N2070), .DIN2(N1080));
nor2s1 U604 (.Q(N2133), .DIN1(N2073), .DIN2(N1128));
nor2s1 U605 (.Q(N2137), .DIN1(N2030), .DIN2(N2076));
nor2s1 U606 (.Q(N2138), .DIN1(N2076), .DIN2(N1176));
nor2s1 U607 (.Q(N2139), .DIN1(N1941), .DIN2(N2076));
nor2s1 U608 (.Q(N2142), .DIN1(N2080), .DIN2(N2081));
nor2s1 U609 (.Q(N2145), .DIN1(N1272), .DIN2(N2082));
nor2s1 U610 (.Q(N2149), .DIN1(N2037), .DIN2(N2085));
nor2s1 U611 (.Q(N2150), .DIN1(N2085), .DIN2(N552));
nor2s1 U612 (.Q(N2151), .DIN1(N1947), .DIN2(N2085));
nor2s1 U613 (.Q(N2154), .DIN1(N2040), .DIN2(N2089));
nor2s1 U614 (.Q(N2155), .DIN1(N2089), .DIN2(N600));
nor2s1 U615 (.Q(N2156), .DIN1(N1951), .DIN2(N2089));
nor2s1 U616 (.Q(N2159), .DIN1(N2043), .DIN2(N2093));
nor2s1 U617 (.Q(N2160), .DIN1(N2093), .DIN2(N648));
nor2s1 U618 (.Q(N2161), .DIN1(N1955), .DIN2(N2093));
nor2s1 U619 (.Q(N2164), .DIN1(N2046), .DIN2(N2097));
nor2s1 U620 (.Q(N2165), .DIN1(N2097), .DIN2(N696));
nor2s1 U621 (.Q(N2166), .DIN1(N1959), .DIN2(N2097));
nor2s1 U622 (.Q(N2169), .DIN1(N2049), .DIN2(N2101));
nor2s1 U623 (.Q(N2170), .DIN1(N2101), .DIN2(N744));
nor2s1 U624 (.Q(N2171), .DIN1(N1963), .DIN2(N2101));
nor2s1 U625 (.Q(N2174), .DIN1(N2052), .DIN2(N2105));
nor2s1 U626 (.Q(N2175), .DIN1(N2105), .DIN2(N792));
nor2s1 U627 (.Q(N2176), .DIN1(N1967), .DIN2(N2105));
nor2s1 U628 (.Q(N2179), .DIN1(N2055), .DIN2(N2109));
nor2s1 U629 (.Q(N2180), .DIN1(N2109), .DIN2(N840));
nor2s1 U630 (.Q(N2181), .DIN1(N1971), .DIN2(N2109));
nor2s1 U631 (.Q(N2184), .DIN1(N2058), .DIN2(N2113));
nor2s1 U632 (.Q(N2185), .DIN1(N2113), .DIN2(N888));
nor2s1 U633 (.Q(N2186), .DIN1(N1975), .DIN2(N2113));
nor2s1 U634 (.Q(N2189), .DIN1(N2061), .DIN2(N2117));
nor2s1 U635 (.Q(N2190), .DIN1(N2117), .DIN2(N936));
nor2s1 U636 (.Q(N2191), .DIN1(N1979), .DIN2(N2117));
nor2s1 U637 (.Q(N2194), .DIN1(N2064), .DIN2(N2121));
nor2s1 U638 (.Q(N2195), .DIN1(N2121), .DIN2(N984));
nor2s1 U639 (.Q(N2196), .DIN1(N1983), .DIN2(N2121));
nor2s1 U640 (.Q(N2199), .DIN1(N2067), .DIN2(N2125));
nor2s1 U641 (.Q(N2200), .DIN1(N2125), .DIN2(N1032));
nor2s1 U642 (.Q(N2201), .DIN1(N1987), .DIN2(N2125));
nor2s1 U643 (.Q(N2204), .DIN1(N2070), .DIN2(N2129));
nor2s1 U644 (.Q(N2205), .DIN1(N2129), .DIN2(N1080));
nor2s1 U645 (.Q(N2206), .DIN1(N1991), .DIN2(N2129));
nor2s1 U646 (.Q(N2209), .DIN1(N2073), .DIN2(N2133));
nor2s1 U647 (.Q(N2210), .DIN1(N2133), .DIN2(N1128));
nor2s1 U648 (.Q(N2211), .DIN1(N1995), .DIN2(N2133));
nor2s1 U649 (.Q(N2214), .DIN1(N2137), .DIN2(N2138));
nor2s1 U650 (.Q(N2217), .DIN1(N2142), .DIN2(N2139));
nor2s1 U651 (.Q(N2221), .DIN1(N1272), .DIN2(N2145));
nor2s1 U652 (.Q(N2222), .DIN1(N2145), .DIN2(N2082));
nor2s1 U653 (.Q(N2223), .DIN1(N2149), .DIN2(N2150));
nor2s1 U654 (.Q(N2224), .DIN1(N2154), .DIN2(N2155));
nor2s1 U655 (.Q(N2227), .DIN1(N2159), .DIN2(N2160));
nor2s1 U656 (.Q(N2230), .DIN1(N2164), .DIN2(N2165));
nor2s1 U657 (.Q(N2233), .DIN1(N2169), .DIN2(N2170));
nor2s1 U658 (.Q(N2236), .DIN1(N2174), .DIN2(N2175));
nor2s1 U659 (.Q(N2239), .DIN1(N2179), .DIN2(N2180));
nor2s1 U660 (.Q(N2242), .DIN1(N2184), .DIN2(N2185));
nor2s1 U661 (.Q(N2245), .DIN1(N2189), .DIN2(N2190));
nor2s1 U662 (.Q(N2248), .DIN1(N2194), .DIN2(N2195));
nor2s1 U663 (.Q(N2251), .DIN1(N2199), .DIN2(N2200));
nor2s1 U664 (.Q(N2254), .DIN1(N2204), .DIN2(N2205));
nor2s1 U665 (.Q(N2257), .DIN1(N2209), .DIN2(N2210));
nor2s1 U666 (.Q(N2260), .DIN1(N2214), .DIN2(N2211));
nor2s1 U667 (.Q(N2264), .DIN1(N2142), .DIN2(N2217));
nor2s1 U668 (.Q(N2265), .DIN1(N2217), .DIN2(N2139));
nor2s1 U669 (.Q(N2266), .DIN1(N2221), .DIN2(N2222));
nor2s1 U670 (.Q(N2269), .DIN1(N2224), .DIN2(N2151));
nor2s1 U671 (.Q(N2273), .DIN1(N2227), .DIN2(N2156));
nor2s1 U672 (.Q(N2277), .DIN1(N2230), .DIN2(N2161));
nor2s1 U673 (.Q(N2281), .DIN1(N2233), .DIN2(N2166));
nor2s1 U674 (.Q(N2285), .DIN1(N2236), .DIN2(N2171));
nor2s1 U675 (.Q(N2289), .DIN1(N2239), .DIN2(N2176));
nor2s1 U676 (.Q(N2293), .DIN1(N2242), .DIN2(N2181));
nor2s1 U677 (.Q(N2297), .DIN1(N2245), .DIN2(N2186));
nor2s1 U678 (.Q(N2301), .DIN1(N2248), .DIN2(N2191));
nor2s1 U679 (.Q(N2305), .DIN1(N2251), .DIN2(N2196));
nor2s1 U680 (.Q(N2309), .DIN1(N2254), .DIN2(N2201));
nor2s1 U681 (.Q(N2313), .DIN1(N2257), .DIN2(N2206));
nor2s1 U682 (.Q(N2317), .DIN1(N2214), .DIN2(N2260));
nor2s1 U683 (.Q(N2318), .DIN1(N2260), .DIN2(N2211));
nor2s1 U684 (.Q(N2319), .DIN1(N2264), .DIN2(N2265));
nor2s1 U685 (.Q(N2322), .DIN1(N2266), .DIN2(N1227));
nor2s1 U686 (.Q(N2326), .DIN1(N2224), .DIN2(N2269));
nor2s1 U687 (.Q(N2327), .DIN1(N2269), .DIN2(N2151));
nor2s1 U688 (.Q(N2328), .DIN1(N2227), .DIN2(N2273));
nor2s1 U689 (.Q(N2329), .DIN1(N2273), .DIN2(N2156));
nor2s1 U690 (.Q(N2330), .DIN1(N2230), .DIN2(N2277));
nor2s1 U691 (.Q(N2331), .DIN1(N2277), .DIN2(N2161));
nor2s1 U692 (.Q(N2332), .DIN1(N2233), .DIN2(N2281));
nor2s1 U693 (.Q(N2333), .DIN1(N2281), .DIN2(N2166));
nor2s1 U694 (.Q(N2334), .DIN1(N2236), .DIN2(N2285));
nor2s1 U695 (.Q(N2335), .DIN1(N2285), .DIN2(N2171));
nor2s1 U696 (.Q(N2336), .DIN1(N2239), .DIN2(N2289));
nor2s1 U697 (.Q(N2337), .DIN1(N2289), .DIN2(N2176));
nor2s1 U698 (.Q(N2338), .DIN1(N2242), .DIN2(N2293));
nor2s1 U699 (.Q(N2339), .DIN1(N2293), .DIN2(N2181));
nor2s1 U700 (.Q(N2340), .DIN1(N2245), .DIN2(N2297));
nor2s1 U701 (.Q(N2341), .DIN1(N2297), .DIN2(N2186));
nor2s1 U702 (.Q(N2342), .DIN1(N2248), .DIN2(N2301));
nor2s1 U703 (.Q(N2343), .DIN1(N2301), .DIN2(N2191));
nor2s1 U704 (.Q(N2344), .DIN1(N2251), .DIN2(N2305));
nor2s1 U705 (.Q(N2345), .DIN1(N2305), .DIN2(N2196));
nor2s1 U706 (.Q(N2346), .DIN1(N2254), .DIN2(N2309));
nor2s1 U707 (.Q(N2347), .DIN1(N2309), .DIN2(N2201));
nor2s1 U708 (.Q(N2348), .DIN1(N2257), .DIN2(N2313));
nor2s1 U709 (.Q(N2349), .DIN1(N2313), .DIN2(N2206));
nor2s1 U710 (.Q(N2350), .DIN1(N2317), .DIN2(N2318));
nor2s1 U711 (.Q(N2353), .DIN1(N2319), .DIN2(N1179));
nor2s1 U712 (.Q(N2357), .DIN1(N2266), .DIN2(N2322));
nor2s1 U713 (.Q(N2358), .DIN1(N2322), .DIN2(N1227));
nor2s1 U714 (.Q(N2359), .DIN1(N2145), .DIN2(N2322));
nor2s1 U715 (.Q(N2362), .DIN1(N2326), .DIN2(N2327));
nor2s1 U716 (.Q(N2365), .DIN1(N2328), .DIN2(N2329));
nor2s1 U717 (.Q(N2368), .DIN1(N2330), .DIN2(N2331));
nor2s1 U718 (.Q(N2371), .DIN1(N2332), .DIN2(N2333));
nor2s1 U719 (.Q(N2374), .DIN1(N2334), .DIN2(N2335));
nor2s1 U720 (.Q(N2377), .DIN1(N2336), .DIN2(N2337));
nor2s1 U721 (.Q(N2380), .DIN1(N2338), .DIN2(N2339));
nor2s1 U722 (.Q(N2383), .DIN1(N2340), .DIN2(N2341));
nor2s1 U723 (.Q(N2386), .DIN1(N2342), .DIN2(N2343));
nor2s1 U724 (.Q(N2389), .DIN1(N2344), .DIN2(N2345));
nor2s1 U725 (.Q(N2392), .DIN1(N2346), .DIN2(N2347));
nor2s1 U726 (.Q(N2395), .DIN1(N2348), .DIN2(N2349));
nor2s1 U727 (.Q(N2398), .DIN1(N2350), .DIN2(N1131));
nor2s1 U728 (.Q(N2402), .DIN1(N2319), .DIN2(N2353));
nor2s1 U729 (.Q(N2403), .DIN1(N2353), .DIN2(N1179));
nor2s1 U730 (.Q(N2404), .DIN1(N2217), .DIN2(N2353));
nor2s1 U731 (.Q(N2407), .DIN1(N2357), .DIN2(N2358));
nor2s1 U732 (.Q(N2410), .DIN1(N1275), .DIN2(N2359));
nor2s1 U733 (.Q(N2414), .DIN1(N2362), .DIN2(N555));
nor2s1 U734 (.Q(N2418), .DIN1(N2365), .DIN2(N603));
nor2s1 U735 (.Q(N2422), .DIN1(N2368), .DIN2(N651));
nor2s1 U736 (.Q(N2426), .DIN1(N2371), .DIN2(N699));
nor2s1 U737 (.Q(N2430), .DIN1(N2374), .DIN2(N747));
nor2s1 U738 (.Q(N2434), .DIN1(N2377), .DIN2(N795));
nor2s1 U739 (.Q(N2438), .DIN1(N2380), .DIN2(N843));
nor2s1 U740 (.Q(N2442), .DIN1(N2383), .DIN2(N891));
nor2s1 U741 (.Q(N2446), .DIN1(N2386), .DIN2(N939));
nor2s1 U742 (.Q(N2450), .DIN1(N2389), .DIN2(N987));
nor2s1 U743 (.Q(N2454), .DIN1(N2392), .DIN2(N1035));
nor2s1 U744 (.Q(N2458), .DIN1(N2395), .DIN2(N1083));
nor2s1 U745 (.Q(N2462), .DIN1(N2350), .DIN2(N2398));
nor2s1 U746 (.Q(N2463), .DIN1(N2398), .DIN2(N1131));
nor2s1 U747 (.Q(N2464), .DIN1(N2260), .DIN2(N2398));
nor2s1 U748 (.Q(N2467), .DIN1(N2402), .DIN2(N2403));
nor2s1 U749 (.Q(N2470), .DIN1(N2407), .DIN2(N2404));
nor2s1 U750 (.Q(N2474), .DIN1(N1275), .DIN2(N2410));
nor2s1 U751 (.Q(N2475), .DIN1(N2410), .DIN2(N2359));
nor2s1 U752 (.Q(N2476), .DIN1(N2362), .DIN2(N2414));
nor2s1 U753 (.Q(N2477), .DIN1(N2414), .DIN2(N555));
nor2s1 U754 (.Q(N2478), .DIN1(N2269), .DIN2(N2414));
nor2s1 U755 (.Q(N2481), .DIN1(N2365), .DIN2(N2418));
nor2s1 U756 (.Q(N2482), .DIN1(N2418), .DIN2(N603));
nor2s1 U757 (.Q(N2483), .DIN1(N2273), .DIN2(N2418));
nor2s1 U758 (.Q(N2486), .DIN1(N2368), .DIN2(N2422));
nor2s1 U759 (.Q(N2487), .DIN1(N2422), .DIN2(N651));
nor2s1 U760 (.Q(N2488), .DIN1(N2277), .DIN2(N2422));
nor2s1 U761 (.Q(N2491), .DIN1(N2371), .DIN2(N2426));
nor2s1 U762 (.Q(N2492), .DIN1(N2426), .DIN2(N699));
nor2s1 U763 (.Q(N2493), .DIN1(N2281), .DIN2(N2426));
nor2s1 U764 (.Q(N2496), .DIN1(N2374), .DIN2(N2430));
nor2s1 U765 (.Q(N2497), .DIN1(N2430), .DIN2(N747));
nor2s1 U766 (.Q(N2498), .DIN1(N2285), .DIN2(N2430));
nor2s1 U767 (.Q(N2501), .DIN1(N2377), .DIN2(N2434));
nor2s1 U768 (.Q(N2502), .DIN1(N2434), .DIN2(N795));
nor2s1 U769 (.Q(N2503), .DIN1(N2289), .DIN2(N2434));
nor2s1 U770 (.Q(N2506), .DIN1(N2380), .DIN2(N2438));
nor2s1 U771 (.Q(N2507), .DIN1(N2438), .DIN2(N843));
nor2s1 U772 (.Q(N2508), .DIN1(N2293), .DIN2(N2438));
nor2s1 U773 (.Q(N2511), .DIN1(N2383), .DIN2(N2442));
nor2s1 U774 (.Q(N2512), .DIN1(N2442), .DIN2(N891));
nor2s1 U775 (.Q(N2513), .DIN1(N2297), .DIN2(N2442));
nor2s1 U776 (.Q(N2516), .DIN1(N2386), .DIN2(N2446));
nor2s1 U777 (.Q(N2517), .DIN1(N2446), .DIN2(N939));
nor2s1 U778 (.Q(N2518), .DIN1(N2301), .DIN2(N2446));
nor2s1 U779 (.Q(N2521), .DIN1(N2389), .DIN2(N2450));
nor2s1 U780 (.Q(N2522), .DIN1(N2450), .DIN2(N987));
nor2s1 U781 (.Q(N2523), .DIN1(N2305), .DIN2(N2450));
nor2s1 U782 (.Q(N2526), .DIN1(N2392), .DIN2(N2454));
nor2s1 U783 (.Q(N2527), .DIN1(N2454), .DIN2(N1035));
nor2s1 U784 (.Q(N2528), .DIN1(N2309), .DIN2(N2454));
nor2s1 U785 (.Q(N2531), .DIN1(N2395), .DIN2(N2458));
nor2s1 U786 (.Q(N2532), .DIN1(N2458), .DIN2(N1083));
nor2s1 U787 (.Q(N2533), .DIN1(N2313), .DIN2(N2458));
nor2s1 U788 (.Q(N2536), .DIN1(N2462), .DIN2(N2463));
nor2s1 U789 (.Q(N2539), .DIN1(N2467), .DIN2(N2464));
nor2s1 U790 (.Q(N2543), .DIN1(N2407), .DIN2(N2470));
nor2s1 U791 (.Q(N2544), .DIN1(N2470), .DIN2(N2404));
nor2s1 U792 (.Q(N2545), .DIN1(N2474), .DIN2(N2475));
nor2s1 U793 (.Q(N2548), .DIN1(N2476), .DIN2(N2477));
nor2s1 U794 (.Q(N2549), .DIN1(N2481), .DIN2(N2482));
nor2s1 U795 (.Q(N2552), .DIN1(N2486), .DIN2(N2487));
nor2s1 U796 (.Q(N2555), .DIN1(N2491), .DIN2(N2492));
nor2s1 U797 (.Q(N2558), .DIN1(N2496), .DIN2(N2497));
nor2s1 U798 (.Q(N2561), .DIN1(N2501), .DIN2(N2502));
nor2s1 U799 (.Q(N2564), .DIN1(N2506), .DIN2(N2507));
nor2s1 U800 (.Q(N2567), .DIN1(N2511), .DIN2(N2512));
nor2s1 U801 (.Q(N2570), .DIN1(N2516), .DIN2(N2517));
nor2s1 U802 (.Q(N2573), .DIN1(N2521), .DIN2(N2522));
nor2s1 U803 (.Q(N2576), .DIN1(N2526), .DIN2(N2527));
nor2s1 U804 (.Q(N2579), .DIN1(N2531), .DIN2(N2532));
nor2s1 U805 (.Q(N2582), .DIN1(N2536), .DIN2(N2533));
nor2s1 U806 (.Q(N2586), .DIN1(N2467), .DIN2(N2539));
nor2s1 U807 (.Q(N2587), .DIN1(N2539), .DIN2(N2464));
nor2s1 U808 (.Q(N2588), .DIN1(N2543), .DIN2(N2544));
nor2s1 U809 (.Q(N2591), .DIN1(N2545), .DIN2(N1230));
nor2s1 U810 (.Q(N2595), .DIN1(N2549), .DIN2(N2478));
nor2s1 U811 (.Q(N2599), .DIN1(N2552), .DIN2(N2483));
nor2s1 U812 (.Q(N2603), .DIN1(N2555), .DIN2(N2488));
nor2s1 U813 (.Q(N2607), .DIN1(N2558), .DIN2(N2493));
nor2s1 U814 (.Q(N2611), .DIN1(N2561), .DIN2(N2498));
nor2s1 U815 (.Q(N2615), .DIN1(N2564), .DIN2(N2503));
nor2s1 U816 (.Q(N2619), .DIN1(N2567), .DIN2(N2508));
nor2s1 U817 (.Q(N2623), .DIN1(N2570), .DIN2(N2513));
nor2s1 U818 (.Q(N2627), .DIN1(N2573), .DIN2(N2518));
nor2s1 U819 (.Q(N2631), .DIN1(N2576), .DIN2(N2523));
nor2s1 U820 (.Q(N2635), .DIN1(N2579), .DIN2(N2528));
nor2s1 U821 (.Q(N2639), .DIN1(N2536), .DIN2(N2582));
nor2s1 U822 (.Q(N2640), .DIN1(N2582), .DIN2(N2533));
nor2s1 U823 (.Q(N2641), .DIN1(N2586), .DIN2(N2587));
nor2s1 U824 (.Q(N2644), .DIN1(N2588), .DIN2(N1182));
nor2s1 U825 (.Q(N2648), .DIN1(N2545), .DIN2(N2591));
nor2s1 U826 (.Q(N2649), .DIN1(N2591), .DIN2(N1230));
nor2s1 U827 (.Q(N2650), .DIN1(N2410), .DIN2(N2591));
nor2s1 U828 (.Q(N2653), .DIN1(N2549), .DIN2(N2595));
nor2s1 U829 (.Q(N2654), .DIN1(N2595), .DIN2(N2478));
nor2s1 U830 (.Q(N2655), .DIN1(N2552), .DIN2(N2599));
nor2s1 U831 (.Q(N2656), .DIN1(N2599), .DIN2(N2483));
nor2s1 U832 (.Q(N2657), .DIN1(N2555), .DIN2(N2603));
nor2s1 U833 (.Q(N2658), .DIN1(N2603), .DIN2(N2488));
nor2s1 U834 (.Q(N2659), .DIN1(N2558), .DIN2(N2607));
nor2s1 U835 (.Q(N2660), .DIN1(N2607), .DIN2(N2493));
nor2s1 U836 (.Q(N2661), .DIN1(N2561), .DIN2(N2611));
nor2s1 U837 (.Q(N2662), .DIN1(N2611), .DIN2(N2498));
nor2s1 U838 (.Q(N2663), .DIN1(N2564), .DIN2(N2615));
nor2s1 U839 (.Q(N2664), .DIN1(N2615), .DIN2(N2503));
nor2s1 U840 (.Q(N2665), .DIN1(N2567), .DIN2(N2619));
nor2s1 U841 (.Q(N2666), .DIN1(N2619), .DIN2(N2508));
nor2s1 U842 (.Q(N2667), .DIN1(N2570), .DIN2(N2623));
nor2s1 U843 (.Q(N2668), .DIN1(N2623), .DIN2(N2513));
nor2s1 U844 (.Q(N2669), .DIN1(N2573), .DIN2(N2627));
nor2s1 U845 (.Q(N2670), .DIN1(N2627), .DIN2(N2518));
nor2s1 U846 (.Q(N2671), .DIN1(N2576), .DIN2(N2631));
nor2s1 U847 (.Q(N2672), .DIN1(N2631), .DIN2(N2523));
nor2s1 U848 (.Q(N2673), .DIN1(N2579), .DIN2(N2635));
nor2s1 U849 (.Q(N2674), .DIN1(N2635), .DIN2(N2528));
nor2s1 U850 (.Q(N2675), .DIN1(N2639), .DIN2(N2640));
nor2s1 U851 (.Q(N2678), .DIN1(N2641), .DIN2(N1134));
nor2s1 U852 (.Q(N2682), .DIN1(N2588), .DIN2(N2644));
nor2s1 U853 (.Q(N2683), .DIN1(N2644), .DIN2(N1182));
nor2s1 U854 (.Q(N2684), .DIN1(N2470), .DIN2(N2644));
nor2s1 U855 (.Q(N2687), .DIN1(N2648), .DIN2(N2649));
nor2s1 U856 (.Q(N2690), .DIN1(N1278), .DIN2(N2650));
nor2s1 U857 (.Q(N2694), .DIN1(N2653), .DIN2(N2654));
nor2s1 U858 (.Q(N2697), .DIN1(N2655), .DIN2(N2656));
nor2s1 U859 (.Q(N2700), .DIN1(N2657), .DIN2(N2658));
nor2s1 U860 (.Q(N2703), .DIN1(N2659), .DIN2(N2660));
nor2s1 U861 (.Q(N2706), .DIN1(N2661), .DIN2(N2662));
nor2s1 U862 (.Q(N2709), .DIN1(N2663), .DIN2(N2664));
nor2s1 U863 (.Q(N2712), .DIN1(N2665), .DIN2(N2666));
nor2s1 U864 (.Q(N2715), .DIN1(N2667), .DIN2(N2668));
nor2s1 U865 (.Q(N2718), .DIN1(N2669), .DIN2(N2670));
nor2s1 U866 (.Q(N2721), .DIN1(N2671), .DIN2(N2672));
nor2s1 U867 (.Q(N2724), .DIN1(N2673), .DIN2(N2674));
nor2s1 U868 (.Q(N2727), .DIN1(N2675), .DIN2(N1086));
nor2s1 U869 (.Q(N2731), .DIN1(N2641), .DIN2(N2678));
nor2s1 U870 (.Q(N2732), .DIN1(N2678), .DIN2(N1134));
nor2s1 U871 (.Q(N2733), .DIN1(N2539), .DIN2(N2678));
nor2s1 U872 (.Q(N2736), .DIN1(N2682), .DIN2(N2683));
nor2s1 U873 (.Q(N2739), .DIN1(N2687), .DIN2(N2684));
nor2s1 U874 (.Q(N2743), .DIN1(N1278), .DIN2(N2690));
nor2s1 U875 (.Q(N2744), .DIN1(N2690), .DIN2(N2650));
nor2s1 U876 (.Q(N2745), .DIN1(N2694), .DIN2(N558));
nor2s1 U877 (.Q(N2749), .DIN1(N2697), .DIN2(N606));
nor2s1 U878 (.Q(N2753), .DIN1(N2700), .DIN2(N654));
nor2s1 U879 (.Q(N2757), .DIN1(N2703), .DIN2(N702));
nor2s1 U880 (.Q(N2761), .DIN1(N2706), .DIN2(N750));
nor2s1 U881 (.Q(N2765), .DIN1(N2709), .DIN2(N798));
nor2s1 U882 (.Q(N2769), .DIN1(N2712), .DIN2(N846));
nor2s1 U883 (.Q(N2773), .DIN1(N2715), .DIN2(N894));
nor2s1 U884 (.Q(N2777), .DIN1(N2718), .DIN2(N942));
nor2s1 U885 (.Q(N2781), .DIN1(N2721), .DIN2(N990));
nor2s1 U886 (.Q(N2785), .DIN1(N2724), .DIN2(N1038));
nor2s1 U887 (.Q(N2789), .DIN1(N2675), .DIN2(N2727));
nor2s1 U888 (.Q(N2790), .DIN1(N2727), .DIN2(N1086));
nor2s1 U889 (.Q(N2791), .DIN1(N2582), .DIN2(N2727));
nor2s1 U890 (.Q(N2794), .DIN1(N2731), .DIN2(N2732));
nor2s1 U891 (.Q(N2797), .DIN1(N2736), .DIN2(N2733));
nor2s1 U892 (.Q(N2801), .DIN1(N2687), .DIN2(N2739));
nor2s1 U893 (.Q(N2802), .DIN1(N2739), .DIN2(N2684));
nor2s1 U894 (.Q(N2803), .DIN1(N2743), .DIN2(N2744));
nor2s1 U895 (.Q(N2806), .DIN1(N2694), .DIN2(N2745));
nor2s1 U896 (.Q(N2807), .DIN1(N2745), .DIN2(N558));
nor2s1 U897 (.Q(N2808), .DIN1(N2595), .DIN2(N2745));
nor2s1 U898 (.Q(N2811), .DIN1(N2697), .DIN2(N2749));
nor2s1 U899 (.Q(N2812), .DIN1(N2749), .DIN2(N606));
nor2s1 U900 (.Q(N2813), .DIN1(N2599), .DIN2(N2749));
nor2s1 U901 (.Q(N2816), .DIN1(N2700), .DIN2(N2753));
nor2s1 U902 (.Q(N2817), .DIN1(N2753), .DIN2(N654));
nor2s1 U903 (.Q(N2818), .DIN1(N2603), .DIN2(N2753));
nor2s1 U904 (.Q(N2821), .DIN1(N2703), .DIN2(N2757));
nor2s1 U905 (.Q(N2822), .DIN1(N2757), .DIN2(N702));
nor2s1 U906 (.Q(N2823), .DIN1(N2607), .DIN2(N2757));
nor2s1 U907 (.Q(N2826), .DIN1(N2706), .DIN2(N2761));
nor2s1 U908 (.Q(N2827), .DIN1(N2761), .DIN2(N750));
nor2s1 U909 (.Q(N2828), .DIN1(N2611), .DIN2(N2761));
nor2s1 U910 (.Q(N2831), .DIN1(N2709), .DIN2(N2765));
nor2s1 U911 (.Q(N2832), .DIN1(N2765), .DIN2(N798));
nor2s1 U912 (.Q(N2833), .DIN1(N2615), .DIN2(N2765));
nor2s1 U913 (.Q(N2836), .DIN1(N2712), .DIN2(N2769));
nor2s1 U914 (.Q(N2837), .DIN1(N2769), .DIN2(N846));
nor2s1 U915 (.Q(N2838), .DIN1(N2619), .DIN2(N2769));
nor2s1 U916 (.Q(N2841), .DIN1(N2715), .DIN2(N2773));
nor2s1 U917 (.Q(N2842), .DIN1(N2773), .DIN2(N894));
nor2s1 U918 (.Q(N2843), .DIN1(N2623), .DIN2(N2773));
nor2s1 U919 (.Q(N2846), .DIN1(N2718), .DIN2(N2777));
nor2s1 U920 (.Q(N2847), .DIN1(N2777), .DIN2(N942));
nor2s1 U921 (.Q(N2848), .DIN1(N2627), .DIN2(N2777));
nor2s1 U922 (.Q(N2851), .DIN1(N2721), .DIN2(N2781));
nor2s1 U923 (.Q(N2852), .DIN1(N2781), .DIN2(N990));
nor2s1 U924 (.Q(N2853), .DIN1(N2631), .DIN2(N2781));
nor2s1 U925 (.Q(N2856), .DIN1(N2724), .DIN2(N2785));
nor2s1 U926 (.Q(N2857), .DIN1(N2785), .DIN2(N1038));
nor2s1 U927 (.Q(N2858), .DIN1(N2635), .DIN2(N2785));
nor2s1 U928 (.Q(N2861), .DIN1(N2789), .DIN2(N2790));
nor2s1 U929 (.Q(N2864), .DIN1(N2794), .DIN2(N2791));
nor2s1 U930 (.Q(N2868), .DIN1(N2736), .DIN2(N2797));
nor2s1 U931 (.Q(N2869), .DIN1(N2797), .DIN2(N2733));
nor2s1 U932 (.Q(N2870), .DIN1(N2801), .DIN2(N2802));
nor2s1 U933 (.Q(N2873), .DIN1(N2803), .DIN2(N1233));
nor2s1 U934 (.Q(N2877), .DIN1(N2806), .DIN2(N2807));
nor2s1 U935 (.Q(N2878), .DIN1(N2811), .DIN2(N2812));
nor2s1 U936 (.Q(N2881), .DIN1(N2816), .DIN2(N2817));
nor2s1 U937 (.Q(N2884), .DIN1(N2821), .DIN2(N2822));
nor2s1 U938 (.Q(N2887), .DIN1(N2826), .DIN2(N2827));
nor2s1 U939 (.Q(N2890), .DIN1(N2831), .DIN2(N2832));
nor2s1 U940 (.Q(N2893), .DIN1(N2836), .DIN2(N2837));
nor2s1 U941 (.Q(N2896), .DIN1(N2841), .DIN2(N2842));
nor2s1 U942 (.Q(N2899), .DIN1(N2846), .DIN2(N2847));
nor2s1 U943 (.Q(N2902), .DIN1(N2851), .DIN2(N2852));
nor2s1 U944 (.Q(N2905), .DIN1(N2856), .DIN2(N2857));
nor2s1 U945 (.Q(N2908), .DIN1(N2861), .DIN2(N2858));
nor2s1 U946 (.Q(N2912), .DIN1(N2794), .DIN2(N2864));
nor2s1 U947 (.Q(N2913), .DIN1(N2864), .DIN2(N2791));
nor2s1 U948 (.Q(N2914), .DIN1(N2868), .DIN2(N2869));
nor2s1 U949 (.Q(N2917), .DIN1(N2870), .DIN2(N1185));
nor2s1 U950 (.Q(N2921), .DIN1(N2803), .DIN2(N2873));
nor2s1 U951 (.Q(N2922), .DIN1(N2873), .DIN2(N1233));
nor2s1 U952 (.Q(N2923), .DIN1(N2690), .DIN2(N2873));
nor2s1 U953 (.Q(N2926), .DIN1(N2878), .DIN2(N2808));
nor2s1 U954 (.Q(N2930), .DIN1(N2881), .DIN2(N2813));
nor2s1 U955 (.Q(N2934), .DIN1(N2884), .DIN2(N2818));
nor2s1 U956 (.Q(N2938), .DIN1(N2887), .DIN2(N2823));
nor2s1 U957 (.Q(N2942), .DIN1(N2890), .DIN2(N2828));
nor2s1 U958 (.Q(N2946), .DIN1(N2893), .DIN2(N2833));
nor2s1 U959 (.Q(N2950), .DIN1(N2896), .DIN2(N2838));
nor2s1 U960 (.Q(N2954), .DIN1(N2899), .DIN2(N2843));
nor2s1 U961 (.Q(N2958), .DIN1(N2902), .DIN2(N2848));
nor2s1 U962 (.Q(N2962), .DIN1(N2905), .DIN2(N2853));
nor2s1 U963 (.Q(N2966), .DIN1(N2861), .DIN2(N2908));
nor2s1 U964 (.Q(N2967), .DIN1(N2908), .DIN2(N2858));
nor2s1 U965 (.Q(N2968), .DIN1(N2912), .DIN2(N2913));
nor2s1 U966 (.Q(N2971), .DIN1(N2914), .DIN2(N1137));
nor2s1 U967 (.Q(N2975), .DIN1(N2870), .DIN2(N2917));
nor2s1 U968 (.Q(N2976), .DIN1(N2917), .DIN2(N1185));
nor2s1 U969 (.Q(N2977), .DIN1(N2739), .DIN2(N2917));
nor2s1 U970 (.Q(N2980), .DIN1(N2921), .DIN2(N2922));
nor2s1 U971 (.Q(N2983), .DIN1(N1281), .DIN2(N2923));
nor2s1 U972 (.Q(N2987), .DIN1(N2878), .DIN2(N2926));
nor2s1 U973 (.Q(N2988), .DIN1(N2926), .DIN2(N2808));
nor2s1 U974 (.Q(N2989), .DIN1(N2881), .DIN2(N2930));
nor2s1 U975 (.Q(N2990), .DIN1(N2930), .DIN2(N2813));
nor2s1 U976 (.Q(N2991), .DIN1(N2884), .DIN2(N2934));
nor2s1 U977 (.Q(N2992), .DIN1(N2934), .DIN2(N2818));
nor2s1 U978 (.Q(N2993), .DIN1(N2887), .DIN2(N2938));
nor2s1 U979 (.Q(N2994), .DIN1(N2938), .DIN2(N2823));
nor2s1 U980 (.Q(N2995), .DIN1(N2890), .DIN2(N2942));
nor2s1 U981 (.Q(N2996), .DIN1(N2942), .DIN2(N2828));
nor2s1 U982 (.Q(N2997), .DIN1(N2893), .DIN2(N2946));
nor2s1 U983 (.Q(N2998), .DIN1(N2946), .DIN2(N2833));
nor2s1 U984 (.Q(N2999), .DIN1(N2896), .DIN2(N2950));
nor2s1 U985 (.Q(N3000), .DIN1(N2950), .DIN2(N2838));
nor2s1 U986 (.Q(N3001), .DIN1(N2899), .DIN2(N2954));
nor2s1 U987 (.Q(N3002), .DIN1(N2954), .DIN2(N2843));
nor2s1 U988 (.Q(N3003), .DIN1(N2902), .DIN2(N2958));
nor2s1 U989 (.Q(N3004), .DIN1(N2958), .DIN2(N2848));
nor2s1 U990 (.Q(N3005), .DIN1(N2905), .DIN2(N2962));
nor2s1 U991 (.Q(N3006), .DIN1(N2962), .DIN2(N2853));
nor2s1 U992 (.Q(N3007), .DIN1(N2966), .DIN2(N2967));
nor2s1 U993 (.Q(N3010), .DIN1(N2968), .DIN2(N1089));
nor2s1 U994 (.Q(N3014), .DIN1(N2914), .DIN2(N2971));
nor2s1 U995 (.Q(N3015), .DIN1(N2971), .DIN2(N1137));
nor2s1 U996 (.Q(N3016), .DIN1(N2797), .DIN2(N2971));
nor2s1 U997 (.Q(N3019), .DIN1(N2975), .DIN2(N2976));
nor2s1 U998 (.Q(N3022), .DIN1(N2980), .DIN2(N2977));
nor2s1 U999 (.Q(N3026), .DIN1(N1281), .DIN2(N2983));
nor2s1 U1000 (.Q(N3027), .DIN1(N2983), .DIN2(N2923));
nor2s1 U1001 (.Q(N3028), .DIN1(N2987), .DIN2(N2988));
nor2s1 U1002 (.Q(N3031), .DIN1(N2989), .DIN2(N2990));
nor2s1 U1003 (.Q(N3034), .DIN1(N2991), .DIN2(N2992));
nor2s1 U1004 (.Q(N3037), .DIN1(N2993), .DIN2(N2994));
nor2s1 U1005 (.Q(N3040), .DIN1(N2995), .DIN2(N2996));
nor2s1 U1006 (.Q(N3043), .DIN1(N2997), .DIN2(N2998));
nor2s1 U1007 (.Q(N3046), .DIN1(N2999), .DIN2(N3000));
nor2s1 U1008 (.Q(N3049), .DIN1(N3001), .DIN2(N3002));
nor2s1 U1009 (.Q(N3052), .DIN1(N3003), .DIN2(N3004));
nor2s1 U1010 (.Q(N3055), .DIN1(N3005), .DIN2(N3006));
nor2s1 U1011 (.Q(N3058), .DIN1(N3007), .DIN2(N1041));
nor2s1 U1012 (.Q(N3062), .DIN1(N2968), .DIN2(N3010));
nor2s1 U1013 (.Q(N3063), .DIN1(N3010), .DIN2(N1089));
nor2s1 U1014 (.Q(N3064), .DIN1(N2864), .DIN2(N3010));
nor2s1 U1015 (.Q(N3067), .DIN1(N3014), .DIN2(N3015));
nor2s1 U1016 (.Q(N3070), .DIN1(N3019), .DIN2(N3016));
nor2s1 U1017 (.Q(N3074), .DIN1(N2980), .DIN2(N3022));
nor2s1 U1018 (.Q(N3075), .DIN1(N3022), .DIN2(N2977));
nor2s1 U1019 (.Q(N3076), .DIN1(N3026), .DIN2(N3027));
nor2s1 U1020 (.Q(N3079), .DIN1(N3028), .DIN2(N561));
nor2s1 U1021 (.Q(N3083), .DIN1(N3031), .DIN2(N609));
nor2s1 U1022 (.Q(N3087), .DIN1(N3034), .DIN2(N657));
nor2s1 U1023 (.Q(N3091), .DIN1(N3037), .DIN2(N705));
nor2s1 U1024 (.Q(N3095), .DIN1(N3040), .DIN2(N753));
nor2s1 U1025 (.Q(N3099), .DIN1(N3043), .DIN2(N801));
nor2s1 U1026 (.Q(N3103), .DIN1(N3046), .DIN2(N849));
nor2s1 U1027 (.Q(N3107), .DIN1(N3049), .DIN2(N897));
nor2s1 U1028 (.Q(N3111), .DIN1(N3052), .DIN2(N945));
nor2s1 U1029 (.Q(N3115), .DIN1(N3055), .DIN2(N993));
nor2s1 U1030 (.Q(N3119), .DIN1(N3007), .DIN2(N3058));
nor2s1 U1031 (.Q(N3120), .DIN1(N3058), .DIN2(N1041));
nor2s1 U1032 (.Q(N3121), .DIN1(N2908), .DIN2(N3058));
nor2s1 U1033 (.Q(N3124), .DIN1(N3062), .DIN2(N3063));
nor2s1 U1034 (.Q(N3127), .DIN1(N3067), .DIN2(N3064));
nor2s1 U1035 (.Q(N3131), .DIN1(N3019), .DIN2(N3070));
nor2s1 U1036 (.Q(N3132), .DIN1(N3070), .DIN2(N3016));
nor2s1 U1037 (.Q(N3133), .DIN1(N3074), .DIN2(N3075));
nor2s1 U1038 (.Q(N3136), .DIN1(N3076), .DIN2(N1236));
nor2s1 U1039 (.Q(N3140), .DIN1(N3028), .DIN2(N3079));
nor2s1 U1040 (.Q(N3141), .DIN1(N3079), .DIN2(N561));
nor2s1 U1041 (.Q(N3142), .DIN1(N2926), .DIN2(N3079));
nor2s1 U1042 (.Q(N3145), .DIN1(N3031), .DIN2(N3083));
nor2s1 U1043 (.Q(N3146), .DIN1(N3083), .DIN2(N609));
nor2s1 U1044 (.Q(N3147), .DIN1(N2930), .DIN2(N3083));
nor2s1 U1045 (.Q(N3150), .DIN1(N3034), .DIN2(N3087));
nor2s1 U1046 (.Q(N3151), .DIN1(N3087), .DIN2(N657));
nor2s1 U1047 (.Q(N3152), .DIN1(N2934), .DIN2(N3087));
nor2s1 U1048 (.Q(N3155), .DIN1(N3037), .DIN2(N3091));
nor2s1 U1049 (.Q(N3156), .DIN1(N3091), .DIN2(N705));
nor2s1 U1050 (.Q(N3157), .DIN1(N2938), .DIN2(N3091));
nor2s1 U1051 (.Q(N3160), .DIN1(N3040), .DIN2(N3095));
nor2s1 U1052 (.Q(N3161), .DIN1(N3095), .DIN2(N753));
nor2s1 U1053 (.Q(N3162), .DIN1(N2942), .DIN2(N3095));
nor2s1 U1054 (.Q(N3165), .DIN1(N3043), .DIN2(N3099));
nor2s1 U1055 (.Q(N3166), .DIN1(N3099), .DIN2(N801));
nor2s1 U1056 (.Q(N3167), .DIN1(N2946), .DIN2(N3099));
nor2s1 U1057 (.Q(N3170), .DIN1(N3046), .DIN2(N3103));
nor2s1 U1058 (.Q(N3171), .DIN1(N3103), .DIN2(N849));
nor2s1 U1059 (.Q(N3172), .DIN1(N2950), .DIN2(N3103));
nor2s1 U1060 (.Q(N3175), .DIN1(N3049), .DIN2(N3107));
nor2s1 U1061 (.Q(N3176), .DIN1(N3107), .DIN2(N897));
nor2s1 U1062 (.Q(N3177), .DIN1(N2954), .DIN2(N3107));
nor2s1 U1063 (.Q(N3180), .DIN1(N3052), .DIN2(N3111));
nor2s1 U1064 (.Q(N3181), .DIN1(N3111), .DIN2(N945));
nor2s1 U1065 (.Q(N3182), .DIN1(N2958), .DIN2(N3111));
nor2s1 U1066 (.Q(N3185), .DIN1(N3055), .DIN2(N3115));
nor2s1 U1067 (.Q(N3186), .DIN1(N3115), .DIN2(N993));
nor2s1 U1068 (.Q(N3187), .DIN1(N2962), .DIN2(N3115));
nor2s1 U1069 (.Q(N3190), .DIN1(N3119), .DIN2(N3120));
nor2s1 U1070 (.Q(N3193), .DIN1(N3124), .DIN2(N3121));
nor2s1 U1071 (.Q(N3197), .DIN1(N3067), .DIN2(N3127));
nor2s1 U1072 (.Q(N3198), .DIN1(N3127), .DIN2(N3064));
nor2s1 U1073 (.Q(N3199), .DIN1(N3131), .DIN2(N3132));
nor2s1 U1074 (.Q(N3202), .DIN1(N3133), .DIN2(N1188));
nor2s1 U1075 (.Q(N3206), .DIN1(N3076), .DIN2(N3136));
nor2s1 U1076 (.Q(N3207), .DIN1(N3136), .DIN2(N1236));
nor2s1 U1077 (.Q(N3208), .DIN1(N2983), .DIN2(N3136));
nor2s1 U1078 (.Q(N3211), .DIN1(N3140), .DIN2(N3141));
nor2s1 U1079 (.Q(N3212), .DIN1(N3145), .DIN2(N3146));
nor2s1 U1080 (.Q(N3215), .DIN1(N3150), .DIN2(N3151));
nor2s1 U1081 (.Q(N3218), .DIN1(N3155), .DIN2(N3156));
nor2s1 U1082 (.Q(N3221), .DIN1(N3160), .DIN2(N3161));
nor2s1 U1083 (.Q(N3224), .DIN1(N3165), .DIN2(N3166));
nor2s1 U1084 (.Q(N3227), .DIN1(N3170), .DIN2(N3171));
nor2s1 U1085 (.Q(N3230), .DIN1(N3175), .DIN2(N3176));
nor2s1 U1086 (.Q(N3233), .DIN1(N3180), .DIN2(N3181));
nor2s1 U1087 (.Q(N3236), .DIN1(N3185), .DIN2(N3186));
nor2s1 U1088 (.Q(N3239), .DIN1(N3190), .DIN2(N3187));
nor2s1 U1089 (.Q(N3243), .DIN1(N3124), .DIN2(N3193));
nor2s1 U1090 (.Q(N3244), .DIN1(N3193), .DIN2(N3121));
nor2s1 U1091 (.Q(N3245), .DIN1(N3197), .DIN2(N3198));
nor2s1 U1092 (.Q(N3248), .DIN1(N3199), .DIN2(N1140));
nor2s1 U1093 (.Q(N3252), .DIN1(N3133), .DIN2(N3202));
nor2s1 U1094 (.Q(N3253), .DIN1(N3202), .DIN2(N1188));
nor2s1 U1095 (.Q(N3254), .DIN1(N3022), .DIN2(N3202));
nor2s1 U1096 (.Q(N3257), .DIN1(N3206), .DIN2(N3207));
nor2s1 U1097 (.Q(N3260), .DIN1(N1284), .DIN2(N3208));
nor2s1 U1098 (.Q(N3264), .DIN1(N3212), .DIN2(N3142));
nor2s1 U1099 (.Q(N3268), .DIN1(N3215), .DIN2(N3147));
nor2s1 U1100 (.Q(N3272), .DIN1(N3218), .DIN2(N3152));
nor2s1 U1101 (.Q(N3276), .DIN1(N3221), .DIN2(N3157));
nor2s1 U1102 (.Q(N3280), .DIN1(N3224), .DIN2(N3162));
nor2s1 U1103 (.Q(N3284), .DIN1(N3227), .DIN2(N3167));
nor2s1 U1104 (.Q(N3288), .DIN1(N3230), .DIN2(N3172));
nor2s1 U1105 (.Q(N3292), .DIN1(N3233), .DIN2(N3177));
nor2s1 U1106 (.Q(N3296), .DIN1(N3236), .DIN2(N3182));
nor2s1 U1107 (.Q(N3300), .DIN1(N3190), .DIN2(N3239));
nor2s1 U1108 (.Q(N3301), .DIN1(N3239), .DIN2(N3187));
nor2s1 U1109 (.Q(N3302), .DIN1(N3243), .DIN2(N3244));
nor2s1 U1110 (.Q(N3305), .DIN1(N3245), .DIN2(N1092));
nor2s1 U1111 (.Q(N3309), .DIN1(N3199), .DIN2(N3248));
nor2s1 U1112 (.Q(N3310), .DIN1(N3248), .DIN2(N1140));
nor2s1 U1113 (.Q(N3311), .DIN1(N3070), .DIN2(N3248));
nor2s1 U1114 (.Q(N3314), .DIN1(N3252), .DIN2(N3253));
nor2s1 U1115 (.Q(N3317), .DIN1(N3257), .DIN2(N3254));
nor2s1 U1116 (.Q(N3321), .DIN1(N1284), .DIN2(N3260));
nor2s1 U1117 (.Q(N3322), .DIN1(N3260), .DIN2(N3208));
nor2s1 U1118 (.Q(N3323), .DIN1(N3212), .DIN2(N3264));
nor2s1 U1119 (.Q(N3324), .DIN1(N3264), .DIN2(N3142));
nor2s1 U1120 (.Q(N3325), .DIN1(N3215), .DIN2(N3268));
nor2s1 U1121 (.Q(N3326), .DIN1(N3268), .DIN2(N3147));
nor2s1 U1122 (.Q(N3327), .DIN1(N3218), .DIN2(N3272));
nor2s1 U1123 (.Q(N3328), .DIN1(N3272), .DIN2(N3152));
nor2s1 U1124 (.Q(N3329), .DIN1(N3221), .DIN2(N3276));
nor2s1 U1125 (.Q(N3330), .DIN1(N3276), .DIN2(N3157));
nor2s1 U1126 (.Q(N3331), .DIN1(N3224), .DIN2(N3280));
nor2s1 U1127 (.Q(N3332), .DIN1(N3280), .DIN2(N3162));
nor2s1 U1128 (.Q(N3333), .DIN1(N3227), .DIN2(N3284));
nor2s1 U1129 (.Q(N3334), .DIN1(N3284), .DIN2(N3167));
nor2s1 U1130 (.Q(N3335), .DIN1(N3230), .DIN2(N3288));
nor2s1 U1131 (.Q(N3336), .DIN1(N3288), .DIN2(N3172));
nor2s1 U1132 (.Q(N3337), .DIN1(N3233), .DIN2(N3292));
nor2s1 U1133 (.Q(N3338), .DIN1(N3292), .DIN2(N3177));
nor2s1 U1134 (.Q(N3339), .DIN1(N3236), .DIN2(N3296));
nor2s1 U1135 (.Q(N3340), .DIN1(N3296), .DIN2(N3182));
nor2s1 U1136 (.Q(N3341), .DIN1(N3300), .DIN2(N3301));
nor2s1 U1137 (.Q(N3344), .DIN1(N3302), .DIN2(N1044));
nor2s1 U1138 (.Q(N3348), .DIN1(N3245), .DIN2(N3305));
nor2s1 U1139 (.Q(N3349), .DIN1(N3305), .DIN2(N1092));
nor2s1 U1140 (.Q(N3350), .DIN1(N3127), .DIN2(N3305));
nor2s1 U1141 (.Q(N3353), .DIN1(N3309), .DIN2(N3310));
nor2s1 U1142 (.Q(N3356), .DIN1(N3314), .DIN2(N3311));
nor2s1 U1143 (.Q(N3360), .DIN1(N3257), .DIN2(N3317));
nor2s1 U1144 (.Q(N3361), .DIN1(N3317), .DIN2(N3254));
nor2s1 U1145 (.Q(N3362), .DIN1(N3321), .DIN2(N3322));
nor2s1 U1146 (.Q(N3365), .DIN1(N3323), .DIN2(N3324));
nor2s1 U1147 (.Q(N3368), .DIN1(N3325), .DIN2(N3326));
nor2s1 U1148 (.Q(N3371), .DIN1(N3327), .DIN2(N3328));
nor2s1 U1149 (.Q(N3374), .DIN1(N3329), .DIN2(N3330));
nor2s1 U1150 (.Q(N3377), .DIN1(N3331), .DIN2(N3332));
nor2s1 U1151 (.Q(N3380), .DIN1(N3333), .DIN2(N3334));
nor2s1 U1152 (.Q(N3383), .DIN1(N3335), .DIN2(N3336));
nor2s1 U1153 (.Q(N3386), .DIN1(N3337), .DIN2(N3338));
nor2s1 U1154 (.Q(N3389), .DIN1(N3339), .DIN2(N3340));
nor2s1 U1155 (.Q(N3392), .DIN1(N3341), .DIN2(N996));
nor2s1 U1156 (.Q(N3396), .DIN1(N3302), .DIN2(N3344));
nor2s1 U1157 (.Q(N3397), .DIN1(N3344), .DIN2(N1044));
nor2s1 U1158 (.Q(N3398), .DIN1(N3193), .DIN2(N3344));
nor2s1 U1159 (.Q(N3401), .DIN1(N3348), .DIN2(N3349));
nor2s1 U1160 (.Q(N3404), .DIN1(N3353), .DIN2(N3350));
nor2s1 U1161 (.Q(N3408), .DIN1(N3314), .DIN2(N3356));
nor2s1 U1162 (.Q(N3409), .DIN1(N3356), .DIN2(N3311));
nor2s1 U1163 (.Q(N3410), .DIN1(N3360), .DIN2(N3361));
nor2s1 U1164 (.Q(N3413), .DIN1(N3362), .DIN2(N1239));
nor2s1 U1165 (.Q(N3417), .DIN1(N3365), .DIN2(N564));
nor2s1 U1166 (.Q(N3421), .DIN1(N3368), .DIN2(N612));
nor2s1 U1167 (.Q(N3425), .DIN1(N3371), .DIN2(N660));
nor2s1 U1168 (.Q(N3429), .DIN1(N3374), .DIN2(N708));
nor2s1 U1169 (.Q(N3433), .DIN1(N3377), .DIN2(N756));
nor2s1 U1170 (.Q(N3437), .DIN1(N3380), .DIN2(N804));
nor2s1 U1171 (.Q(N3441), .DIN1(N3383), .DIN2(N852));
nor2s1 U1172 (.Q(N3445), .DIN1(N3386), .DIN2(N900));
nor2s1 U1173 (.Q(N3449), .DIN1(N3389), .DIN2(N948));
nor2s1 U1174 (.Q(N3453), .DIN1(N3341), .DIN2(N3392));
nor2s1 U1175 (.Q(N3454), .DIN1(N3392), .DIN2(N996));
nor2s1 U1176 (.Q(N3455), .DIN1(N3239), .DIN2(N3392));
nor2s1 U1177 (.Q(N3458), .DIN1(N3396), .DIN2(N3397));
nor2s1 U1178 (.Q(N3461), .DIN1(N3401), .DIN2(N3398));
nor2s1 U1179 (.Q(N3465), .DIN1(N3353), .DIN2(N3404));
nor2s1 U1180 (.Q(N3466), .DIN1(N3404), .DIN2(N3350));
nor2s1 U1181 (.Q(N3467), .DIN1(N3408), .DIN2(N3409));
nor2s1 U1182 (.Q(N3470), .DIN1(N3410), .DIN2(N1191));
nor2s1 U1183 (.Q(N3474), .DIN1(N3362), .DIN2(N3413));
nor2s1 U1184 (.Q(N3475), .DIN1(N3413), .DIN2(N1239));
nor2s1 U1185 (.Q(N3476), .DIN1(N3260), .DIN2(N3413));
nor2s1 U1186 (.Q(N3479), .DIN1(N3365), .DIN2(N3417));
nor2s1 U1187 (.Q(N3480), .DIN1(N3417), .DIN2(N564));
nor2s1 U1188 (.Q(N3481), .DIN1(N3264), .DIN2(N3417));
nor2s1 U1189 (.Q(N3484), .DIN1(N3368), .DIN2(N3421));
nor2s1 U1190 (.Q(N3485), .DIN1(N3421), .DIN2(N612));
nor2s1 U1191 (.Q(N3486), .DIN1(N3268), .DIN2(N3421));
nor2s1 U1192 (.Q(N3489), .DIN1(N3371), .DIN2(N3425));
nor2s1 U1193 (.Q(N3490), .DIN1(N3425), .DIN2(N660));
nor2s1 U1194 (.Q(N3491), .DIN1(N3272), .DIN2(N3425));
nor2s1 U1195 (.Q(N3494), .DIN1(N3374), .DIN2(N3429));
nor2s1 U1196 (.Q(N3495), .DIN1(N3429), .DIN2(N708));
nor2s1 U1197 (.Q(N3496), .DIN1(N3276), .DIN2(N3429));
nor2s1 U1198 (.Q(N3499), .DIN1(N3377), .DIN2(N3433));
nor2s1 U1199 (.Q(N3500), .DIN1(N3433), .DIN2(N756));
nor2s1 U1200 (.Q(N3501), .DIN1(N3280), .DIN2(N3433));
nor2s1 U1201 (.Q(N3504), .DIN1(N3380), .DIN2(N3437));
nor2s1 U1202 (.Q(N3505), .DIN1(N3437), .DIN2(N804));
nor2s1 U1203 (.Q(N3506), .DIN1(N3284), .DIN2(N3437));
nor2s1 U1204 (.Q(N3509), .DIN1(N3383), .DIN2(N3441));
nor2s1 U1205 (.Q(N3510), .DIN1(N3441), .DIN2(N852));
nor2s1 U1206 (.Q(N3511), .DIN1(N3288), .DIN2(N3441));
nor2s1 U1207 (.Q(N3514), .DIN1(N3386), .DIN2(N3445));
nor2s1 U1208 (.Q(N3515), .DIN1(N3445), .DIN2(N900));
nor2s1 U1209 (.Q(N3516), .DIN1(N3292), .DIN2(N3445));
nor2s1 U1210 (.Q(N3519), .DIN1(N3389), .DIN2(N3449));
nor2s1 U1211 (.Q(N3520), .DIN1(N3449), .DIN2(N948));
nor2s1 U1212 (.Q(N3521), .DIN1(N3296), .DIN2(N3449));
nor2s1 U1213 (.Q(N3524), .DIN1(N3453), .DIN2(N3454));
nor2s1 U1214 (.Q(N3527), .DIN1(N3458), .DIN2(N3455));
nor2s1 U1215 (.Q(N3531), .DIN1(N3401), .DIN2(N3461));
nor2s1 U1216 (.Q(N3532), .DIN1(N3461), .DIN2(N3398));
nor2s1 U1217 (.Q(N3533), .DIN1(N3465), .DIN2(N3466));
nor2s1 U1218 (.Q(N3536), .DIN1(N3467), .DIN2(N1143));
nor2s1 U1219 (.Q(N3540), .DIN1(N3410), .DIN2(N3470));
nor2s1 U1220 (.Q(N3541), .DIN1(N3470), .DIN2(N1191));
nor2s1 U1221 (.Q(N3542), .DIN1(N3317), .DIN2(N3470));
nor2s1 U1222 (.Q(N3545), .DIN1(N3474), .DIN2(N3475));
nor2s1 U1223 (.Q(N3548), .DIN1(N1287), .DIN2(N3476));
nor2s1 U1224 (.Q(N3552), .DIN1(N3479), .DIN2(N3480));
nor2s1 U1225 (.Q(N3553), .DIN1(N3484), .DIN2(N3485));
nor2s1 U1226 (.Q(N3556), .DIN1(N3489), .DIN2(N3490));
nor2s1 U1227 (.Q(N3559), .DIN1(N3494), .DIN2(N3495));
nor2s1 U1228 (.Q(N3562), .DIN1(N3499), .DIN2(N3500));
nor2s1 U1229 (.Q(N3565), .DIN1(N3504), .DIN2(N3505));
nor2s1 U1230 (.Q(N3568), .DIN1(N3509), .DIN2(N3510));
nor2s1 U1231 (.Q(N3571), .DIN1(N3514), .DIN2(N3515));
nor2s1 U1232 (.Q(N3574), .DIN1(N3519), .DIN2(N3520));
nor2s1 U1233 (.Q(N3577), .DIN1(N3524), .DIN2(N3521));
nor2s1 U1234 (.Q(N3581), .DIN1(N3458), .DIN2(N3527));
nor2s1 U1235 (.Q(N3582), .DIN1(N3527), .DIN2(N3455));
nor2s1 U1236 (.Q(N3583), .DIN1(N3531), .DIN2(N3532));
nor2s1 U1237 (.Q(N3586), .DIN1(N3533), .DIN2(N1095));
nor2s1 U1238 (.Q(N3590), .DIN1(N3467), .DIN2(N3536));
nor2s1 U1239 (.Q(N3591), .DIN1(N3536), .DIN2(N1143));
nor2s1 U1240 (.Q(N3592), .DIN1(N3356), .DIN2(N3536));
nor2s1 U1241 (.Q(N3595), .DIN1(N3540), .DIN2(N3541));
nor2s1 U1242 (.Q(N3598), .DIN1(N3545), .DIN2(N3542));
nor2s1 U1243 (.Q(N3602), .DIN1(N1287), .DIN2(N3548));
nor2s1 U1244 (.Q(N3603), .DIN1(N3548), .DIN2(N3476));
nor2s1 U1245 (.Q(N3604), .DIN1(N3553), .DIN2(N3481));
nor2s1 U1246 (.Q(N3608), .DIN1(N3556), .DIN2(N3486));
nor2s1 U1247 (.Q(N3612), .DIN1(N3559), .DIN2(N3491));
nor2s1 U1248 (.Q(N3616), .DIN1(N3562), .DIN2(N3496));
nor2s1 U1249 (.Q(N3620), .DIN1(N3565), .DIN2(N3501));
nor2s1 U1250 (.Q(N3624), .DIN1(N3568), .DIN2(N3506));
nor2s1 U1251 (.Q(N3628), .DIN1(N3571), .DIN2(N3511));
nor2s1 U1252 (.Q(N3632), .DIN1(N3574), .DIN2(N3516));
nor2s1 U1253 (.Q(N3636), .DIN1(N3524), .DIN2(N3577));
nor2s1 U1254 (.Q(N3637), .DIN1(N3577), .DIN2(N3521));
nor2s1 U1255 (.Q(N3638), .DIN1(N3581), .DIN2(N3582));
nor2s1 U1256 (.Q(N3641), .DIN1(N3583), .DIN2(N1047));
nor2s1 U1257 (.Q(N3645), .DIN1(N3533), .DIN2(N3586));
nor2s1 U1258 (.Q(N3646), .DIN1(N3586), .DIN2(N1095));
nor2s1 U1259 (.Q(N3647), .DIN1(N3404), .DIN2(N3586));
nor2s1 U1260 (.Q(N3650), .DIN1(N3590), .DIN2(N3591));
nor2s1 U1261 (.Q(N3653), .DIN1(N3595), .DIN2(N3592));
nor2s1 U1262 (.Q(N3657), .DIN1(N3545), .DIN2(N3598));
nor2s1 U1263 (.Q(N3658), .DIN1(N3598), .DIN2(N3542));
nor2s1 U1264 (.Q(N3659), .DIN1(N3602), .DIN2(N3603));
nor2s1 U1265 (.Q(N3662), .DIN1(N3553), .DIN2(N3604));
nor2s1 U1266 (.Q(N3663), .DIN1(N3604), .DIN2(N3481));
nor2s1 U1267 (.Q(N3664), .DIN1(N3556), .DIN2(N3608));
nor2s1 U1268 (.Q(N3665), .DIN1(N3608), .DIN2(N3486));
nor2s1 U1269 (.Q(N3666), .DIN1(N3559), .DIN2(N3612));
nor2s1 U1270 (.Q(N3667), .DIN1(N3612), .DIN2(N3491));
nor2s1 U1271 (.Q(N3668), .DIN1(N3562), .DIN2(N3616));
nor2s1 U1272 (.Q(N3669), .DIN1(N3616), .DIN2(N3496));
nor2s1 U1273 (.Q(N3670), .DIN1(N3565), .DIN2(N3620));
nor2s1 U1274 (.Q(N3671), .DIN1(N3620), .DIN2(N3501));
nor2s1 U1275 (.Q(N3672), .DIN1(N3568), .DIN2(N3624));
nor2s1 U1276 (.Q(N3673), .DIN1(N3624), .DIN2(N3506));
nor2s1 U1277 (.Q(N3674), .DIN1(N3571), .DIN2(N3628));
nor2s1 U1278 (.Q(N3675), .DIN1(N3628), .DIN2(N3511));
nor2s1 U1279 (.Q(N3676), .DIN1(N3574), .DIN2(N3632));
nor2s1 U1280 (.Q(N3677), .DIN1(N3632), .DIN2(N3516));
nor2s1 U1281 (.Q(N3678), .DIN1(N3636), .DIN2(N3637));
nor2s1 U1282 (.Q(N3681), .DIN1(N3638), .DIN2(N999));
nor2s1 U1283 (.Q(N3685), .DIN1(N3583), .DIN2(N3641));
nor2s1 U1284 (.Q(N3686), .DIN1(N3641), .DIN2(N1047));
nor2s1 U1285 (.Q(N3687), .DIN1(N3461), .DIN2(N3641));
nor2s1 U1286 (.Q(N3690), .DIN1(N3645), .DIN2(N3646));
nor2s1 U1287 (.Q(N3693), .DIN1(N3650), .DIN2(N3647));
nor2s1 U1288 (.Q(N3697), .DIN1(N3595), .DIN2(N3653));
nor2s1 U1289 (.Q(N3698), .DIN1(N3653), .DIN2(N3592));
nor2s1 U1290 (.Q(N3699), .DIN1(N3657), .DIN2(N3658));
nor2s1 U1291 (.Q(N3702), .DIN1(N3659), .DIN2(N1242));
nor2s1 U1292 (.Q(N3706), .DIN1(N3662), .DIN2(N3663));
nor2s1 U1293 (.Q(N3709), .DIN1(N3664), .DIN2(N3665));
nor2s1 U1294 (.Q(N3712), .DIN1(N3666), .DIN2(N3667));
nor2s1 U1295 (.Q(N3715), .DIN1(N3668), .DIN2(N3669));
nor2s1 U1296 (.Q(N3718), .DIN1(N3670), .DIN2(N3671));
nor2s1 U1297 (.Q(N3721), .DIN1(N3672), .DIN2(N3673));
nor2s1 U1298 (.Q(N3724), .DIN1(N3674), .DIN2(N3675));
nor2s1 U1299 (.Q(N3727), .DIN1(N3676), .DIN2(N3677));
nor2s1 U1300 (.Q(N3730), .DIN1(N3678), .DIN2(N951));
nor2s1 U1301 (.Q(N3734), .DIN1(N3638), .DIN2(N3681));
nor2s1 U1302 (.Q(N3735), .DIN1(N3681), .DIN2(N999));
nor2s1 U1303 (.Q(N3736), .DIN1(N3527), .DIN2(N3681));
nor2s1 U1304 (.Q(N3739), .DIN1(N3685), .DIN2(N3686));
nor2s1 U1305 (.Q(N3742), .DIN1(N3690), .DIN2(N3687));
nor2s1 U1306 (.Q(N3746), .DIN1(N3650), .DIN2(N3693));
nor2s1 U1307 (.Q(N3747), .DIN1(N3693), .DIN2(N3647));
nor2s1 U1308 (.Q(N3748), .DIN1(N3697), .DIN2(N3698));
nor2s1 U1309 (.Q(N3751), .DIN1(N3699), .DIN2(N1194));
nor2s1 U1310 (.Q(N3755), .DIN1(N3659), .DIN2(N3702));
nor2s1 U1311 (.Q(N3756), .DIN1(N3702), .DIN2(N1242));
nor2s1 U1312 (.Q(N3757), .DIN1(N3548), .DIN2(N3702));
nor2s1 U1313 (.Q(N3760), .DIN1(N3706), .DIN2(N567));
nor2s1 U1314 (.Q(N3764), .DIN1(N3709), .DIN2(N615));
nor2s1 U1315 (.Q(N3768), .DIN1(N3712), .DIN2(N663));
nor2s1 U1316 (.Q(N3772), .DIN1(N3715), .DIN2(N711));
nor2s1 U1317 (.Q(N3776), .DIN1(N3718), .DIN2(N759));
nor2s1 U1318 (.Q(N3780), .DIN1(N3721), .DIN2(N807));
nor2s1 U1319 (.Q(N3784), .DIN1(N3724), .DIN2(N855));
nor2s1 U1320 (.Q(N3788), .DIN1(N3727), .DIN2(N903));
nor2s1 U1321 (.Q(N3792), .DIN1(N3678), .DIN2(N3730));
nor2s1 U1322 (.Q(N3793), .DIN1(N3730), .DIN2(N951));
nor2s1 U1323 (.Q(N3794), .DIN1(N3577), .DIN2(N3730));
nor2s1 U1324 (.Q(N3797), .DIN1(N3734), .DIN2(N3735));
nor2s1 U1325 (.Q(N3800), .DIN1(N3739), .DIN2(N3736));
nor2s1 U1326 (.Q(N3804), .DIN1(N3690), .DIN2(N3742));
nor2s1 U1327 (.Q(N3805), .DIN1(N3742), .DIN2(N3687));
nor2s1 U1328 (.Q(N3806), .DIN1(N3746), .DIN2(N3747));
nor2s1 U1329 (.Q(N3809), .DIN1(N3748), .DIN2(N1146));
nor2s1 U1330 (.Q(N3813), .DIN1(N3699), .DIN2(N3751));
nor2s1 U1331 (.Q(N3814), .DIN1(N3751), .DIN2(N1194));
nor2s1 U1332 (.Q(N3815), .DIN1(N3598), .DIN2(N3751));
nor2s1 U1333 (.Q(N3818), .DIN1(N3755), .DIN2(N3756));
nor2s1 U1334 (.Q(N3821), .DIN1(N1290), .DIN2(N3757));
nor2s1 U1335 (.Q(N3825), .DIN1(N3706), .DIN2(N3760));
nor2s1 U1336 (.Q(N3826), .DIN1(N3760), .DIN2(N567));
nor2s1 U1337 (.Q(N3827), .DIN1(N3604), .DIN2(N3760));
nor2s1 U1338 (.Q(N3830), .DIN1(N3709), .DIN2(N3764));
nor2s1 U1339 (.Q(N3831), .DIN1(N3764), .DIN2(N615));
nor2s1 U1340 (.Q(N3832), .DIN1(N3608), .DIN2(N3764));
nor2s1 U1341 (.Q(N3835), .DIN1(N3712), .DIN2(N3768));
nor2s1 U1342 (.Q(N3836), .DIN1(N3768), .DIN2(N663));
nor2s1 U1343 (.Q(N3837), .DIN1(N3612), .DIN2(N3768));
nor2s1 U1344 (.Q(N3840), .DIN1(N3715), .DIN2(N3772));
nor2s1 U1345 (.Q(N3841), .DIN1(N3772), .DIN2(N711));
nor2s1 U1346 (.Q(N3842), .DIN1(N3616), .DIN2(N3772));
nor2s1 U1347 (.Q(N3845), .DIN1(N3718), .DIN2(N3776));
nor2s1 U1348 (.Q(N3846), .DIN1(N3776), .DIN2(N759));
nor2s1 U1349 (.Q(N3847), .DIN1(N3620), .DIN2(N3776));
nor2s1 U1350 (.Q(N3850), .DIN1(N3721), .DIN2(N3780));
nor2s1 U1351 (.Q(N3851), .DIN1(N3780), .DIN2(N807));
nor2s1 U1352 (.Q(N3852), .DIN1(N3624), .DIN2(N3780));
nor2s1 U1353 (.Q(N3855), .DIN1(N3724), .DIN2(N3784));
nor2s1 U1354 (.Q(N3856), .DIN1(N3784), .DIN2(N855));
nor2s1 U1355 (.Q(N3857), .DIN1(N3628), .DIN2(N3784));
nor2s1 U1356 (.Q(N3860), .DIN1(N3727), .DIN2(N3788));
nor2s1 U1357 (.Q(N3861), .DIN1(N3788), .DIN2(N903));
nor2s1 U1358 (.Q(N3862), .DIN1(N3632), .DIN2(N3788));
nor2s1 U1359 (.Q(N3865), .DIN1(N3792), .DIN2(N3793));
nor2s1 U1360 (.Q(N3868), .DIN1(N3797), .DIN2(N3794));
nor2s1 U1361 (.Q(N3872), .DIN1(N3739), .DIN2(N3800));
nor2s1 U1362 (.Q(N3873), .DIN1(N3800), .DIN2(N3736));
nor2s1 U1363 (.Q(N3874), .DIN1(N3804), .DIN2(N3805));
nor2s1 U1364 (.Q(N3877), .DIN1(N3806), .DIN2(N1098));
nor2s1 U1365 (.Q(N3881), .DIN1(N3748), .DIN2(N3809));
nor2s1 U1366 (.Q(N3882), .DIN1(N3809), .DIN2(N1146));
nor2s1 U1367 (.Q(N3883), .DIN1(N3653), .DIN2(N3809));
nor2s1 U1368 (.Q(N3886), .DIN1(N3813), .DIN2(N3814));
nor2s1 U1369 (.Q(N3889), .DIN1(N3818), .DIN2(N3815));
nor2s1 U1370 (.Q(N3893), .DIN1(N1290), .DIN2(N3821));
nor2s1 U1371 (.Q(N3894), .DIN1(N3821), .DIN2(N3757));
nor2s1 U1372 (.Q(N3895), .DIN1(N3825), .DIN2(N3826));
nor2s1 U1373 (.Q(N3896), .DIN1(N3830), .DIN2(N3831));
nor2s1 U1374 (.Q(N3899), .DIN1(N3835), .DIN2(N3836));
nor2s1 U1375 (.Q(N3902), .DIN1(N3840), .DIN2(N3841));
nor2s1 U1376 (.Q(N3905), .DIN1(N3845), .DIN2(N3846));
nor2s1 U1377 (.Q(N3908), .DIN1(N3850), .DIN2(N3851));
nor2s1 U1378 (.Q(N3911), .DIN1(N3855), .DIN2(N3856));
nor2s1 U1379 (.Q(N3914), .DIN1(N3860), .DIN2(N3861));
nor2s1 U1380 (.Q(N3917), .DIN1(N3865), .DIN2(N3862));
nor2s1 U1381 (.Q(N3921), .DIN1(N3797), .DIN2(N3868));
nor2s1 U1382 (.Q(N3922), .DIN1(N3868), .DIN2(N3794));
nor2s1 U1383 (.Q(N3923), .DIN1(N3872), .DIN2(N3873));
nor2s1 U1384 (.Q(N3926), .DIN1(N3874), .DIN2(N1050));
nor2s1 U1385 (.Q(N3930), .DIN1(N3806), .DIN2(N3877));
nor2s1 U1386 (.Q(N3931), .DIN1(N3877), .DIN2(N1098));
nor2s1 U1387 (.Q(N3932), .DIN1(N3693), .DIN2(N3877));
nor2s1 U1388 (.Q(N3935), .DIN1(N3881), .DIN2(N3882));
nor2s1 U1389 (.Q(N3938), .DIN1(N3886), .DIN2(N3883));
nor2s1 U1390 (.Q(N3942), .DIN1(N3818), .DIN2(N3889));
nor2s1 U1391 (.Q(N3943), .DIN1(N3889), .DIN2(N3815));
nor2s1 U1392 (.Q(N3944), .DIN1(N3893), .DIN2(N3894));
nor2s1 U1393 (.Q(N3947), .DIN1(N3896), .DIN2(N3827));
nor2s1 U1394 (.Q(N3951), .DIN1(N3899), .DIN2(N3832));
nor2s1 U1395 (.Q(N3955), .DIN1(N3902), .DIN2(N3837));
nor2s1 U1396 (.Q(N3959), .DIN1(N3905), .DIN2(N3842));
nor2s1 U1397 (.Q(N3963), .DIN1(N3908), .DIN2(N3847));
nor2s1 U1398 (.Q(N3967), .DIN1(N3911), .DIN2(N3852));
nor2s1 U1399 (.Q(N3971), .DIN1(N3914), .DIN2(N3857));
nor2s1 U1400 (.Q(N3975), .DIN1(N3865), .DIN2(N3917));
nor2s1 U1401 (.Q(N3976), .DIN1(N3917), .DIN2(N3862));
nor2s1 U1402 (.Q(N3977), .DIN1(N3921), .DIN2(N3922));
nor2s1 U1403 (.Q(N3980), .DIN1(N3923), .DIN2(N1002));
nor2s1 U1404 (.Q(N3984), .DIN1(N3874), .DIN2(N3926));
nor2s1 U1405 (.Q(N3985), .DIN1(N3926), .DIN2(N1050));
nor2s1 U1406 (.Q(N3986), .DIN1(N3742), .DIN2(N3926));
nor2s1 U1407 (.Q(N3989), .DIN1(N3930), .DIN2(N3931));
nor2s1 U1408 (.Q(N3992), .DIN1(N3935), .DIN2(N3932));
nor2s1 U1409 (.Q(N3996), .DIN1(N3886), .DIN2(N3938));
nor2s1 U1410 (.Q(N3997), .DIN1(N3938), .DIN2(N3883));
nor2s1 U1411 (.Q(N3998), .DIN1(N3942), .DIN2(N3943));
nor2s1 U1412 (.Q(N4001), .DIN1(N3944), .DIN2(N1245));
nor2s1 U1413 (.Q(N4005), .DIN1(N3896), .DIN2(N3947));
nor2s1 U1414 (.Q(N4006), .DIN1(N3947), .DIN2(N3827));
nor2s1 U1415 (.Q(N4007), .DIN1(N3899), .DIN2(N3951));
nor2s1 U1416 (.Q(N4008), .DIN1(N3951), .DIN2(N3832));
nor2s1 U1417 (.Q(N4009), .DIN1(N3902), .DIN2(N3955));
nor2s1 U1418 (.Q(N4010), .DIN1(N3955), .DIN2(N3837));
nor2s1 U1419 (.Q(N4011), .DIN1(N3905), .DIN2(N3959));
nor2s1 U1420 (.Q(N4012), .DIN1(N3959), .DIN2(N3842));
nor2s1 U1421 (.Q(N4013), .DIN1(N3908), .DIN2(N3963));
nor2s1 U1422 (.Q(N4014), .DIN1(N3963), .DIN2(N3847));
nor2s1 U1423 (.Q(N4015), .DIN1(N3911), .DIN2(N3967));
nor2s1 U1424 (.Q(N4016), .DIN1(N3967), .DIN2(N3852));
nor2s1 U1425 (.Q(N4017), .DIN1(N3914), .DIN2(N3971));
nor2s1 U1426 (.Q(N4018), .DIN1(N3971), .DIN2(N3857));
nor2s1 U1427 (.Q(N4019), .DIN1(N3975), .DIN2(N3976));
nor2s1 U1428 (.Q(N4022), .DIN1(N3977), .DIN2(N954));
nor2s1 U1429 (.Q(N4026), .DIN1(N3923), .DIN2(N3980));
nor2s1 U1430 (.Q(N4027), .DIN1(N3980), .DIN2(N1002));
nor2s1 U1431 (.Q(N4028), .DIN1(N3800), .DIN2(N3980));
nor2s1 U1432 (.Q(N4031), .DIN1(N3984), .DIN2(N3985));
nor2s1 U1433 (.Q(N4034), .DIN1(N3989), .DIN2(N3986));
nor2s1 U1434 (.Q(N4038), .DIN1(N3935), .DIN2(N3992));
nor2s1 U1435 (.Q(N4039), .DIN1(N3992), .DIN2(N3932));
nor2s1 U1436 (.Q(N4040), .DIN1(N3996), .DIN2(N3997));
nor2s1 U1437 (.Q(N4043), .DIN1(N3998), .DIN2(N1197));
nor2s1 U1438 (.Q(N4047), .DIN1(N3944), .DIN2(N4001));
nor2s1 U1439 (.Q(N4048), .DIN1(N4001), .DIN2(N1245));
nor2s1 U1440 (.Q(N4049), .DIN1(N3821), .DIN2(N4001));
nor2s1 U1441 (.Q(N4052), .DIN1(N4005), .DIN2(N4006));
nor2s1 U1442 (.Q(N4055), .DIN1(N4007), .DIN2(N4008));
nor2s1 U1443 (.Q(N4058), .DIN1(N4009), .DIN2(N4010));
nor2s1 U1444 (.Q(N4061), .DIN1(N4011), .DIN2(N4012));
nor2s1 U1445 (.Q(N4064), .DIN1(N4013), .DIN2(N4014));
nor2s1 U1446 (.Q(N4067), .DIN1(N4015), .DIN2(N4016));
nor2s1 U1447 (.Q(N4070), .DIN1(N4017), .DIN2(N4018));
nor2s1 U1448 (.Q(N4073), .DIN1(N4019), .DIN2(N906));
nor2s1 U1449 (.Q(N4077), .DIN1(N3977), .DIN2(N4022));
nor2s1 U1450 (.Q(N4078), .DIN1(N4022), .DIN2(N954));
nor2s1 U1451 (.Q(N4079), .DIN1(N3868), .DIN2(N4022));
nor2s1 U1452 (.Q(N4082), .DIN1(N4026), .DIN2(N4027));
nor2s1 U1453 (.Q(N4085), .DIN1(N4031), .DIN2(N4028));
nor2s1 U1454 (.Q(N4089), .DIN1(N3989), .DIN2(N4034));
nor2s1 U1455 (.Q(N4090), .DIN1(N4034), .DIN2(N3986));
nor2s1 U1456 (.Q(N4091), .DIN1(N4038), .DIN2(N4039));
nor2s1 U1457 (.Q(N4094), .DIN1(N4040), .DIN2(N1149));
nor2s1 U1458 (.Q(N4098), .DIN1(N3998), .DIN2(N4043));
nor2s1 U1459 (.Q(N4099), .DIN1(N4043), .DIN2(N1197));
nor2s1 U1460 (.Q(N4100), .DIN1(N3889), .DIN2(N4043));
nor2s1 U1461 (.Q(N4103), .DIN1(N4047), .DIN2(N4048));
nor2s1 U1462 (.Q(N4106), .DIN1(N1293), .DIN2(N4049));
nor2s1 U1463 (.Q(N4110), .DIN1(N4052), .DIN2(N570));
nor2s1 U1464 (.Q(N4114), .DIN1(N4055), .DIN2(N618));
nor2s1 U1465 (.Q(N4118), .DIN1(N4058), .DIN2(N666));
nor2s1 U1466 (.Q(N4122), .DIN1(N4061), .DIN2(N714));
nor2s1 U1467 (.Q(N4126), .DIN1(N4064), .DIN2(N762));
nor2s1 U1468 (.Q(N4130), .DIN1(N4067), .DIN2(N810));
nor2s1 U1469 (.Q(N4134), .DIN1(N4070), .DIN2(N858));
nor2s1 U1470 (.Q(N4138), .DIN1(N4019), .DIN2(N4073));
nor2s1 U1471 (.Q(N4139), .DIN1(N4073), .DIN2(N906));
nor2s1 U1472 (.Q(N4140), .DIN1(N3917), .DIN2(N4073));
nor2s1 U1473 (.Q(N4143), .DIN1(N4077), .DIN2(N4078));
nor2s1 U1474 (.Q(N4146), .DIN1(N4082), .DIN2(N4079));
nor2s1 U1475 (.Q(N4150), .DIN1(N4031), .DIN2(N4085));
nor2s1 U1476 (.Q(N4151), .DIN1(N4085), .DIN2(N4028));
nor2s1 U1477 (.Q(N4152), .DIN1(N4089), .DIN2(N4090));
nor2s1 U1478 (.Q(N4155), .DIN1(N4091), .DIN2(N1101));
nor2s1 U1479 (.Q(N4159), .DIN1(N4040), .DIN2(N4094));
nor2s1 U1480 (.Q(N4160), .DIN1(N4094), .DIN2(N1149));
nor2s1 U1481 (.Q(N4161), .DIN1(N3938), .DIN2(N4094));
nor2s1 U1482 (.Q(N4164), .DIN1(N4098), .DIN2(N4099));
nor2s1 U1483 (.Q(N4167), .DIN1(N4103), .DIN2(N4100));
nor2s1 U1484 (.Q(N4171), .DIN1(N1293), .DIN2(N4106));
nor2s1 U1485 (.Q(N4172), .DIN1(N4106), .DIN2(N4049));
nor2s1 U1486 (.Q(N4173), .DIN1(N4052), .DIN2(N4110));
nor2s1 U1487 (.Q(N4174), .DIN1(N4110), .DIN2(N570));
nor2s1 U1488 (.Q(N4175), .DIN1(N3947), .DIN2(N4110));
nor2s1 U1489 (.Q(N4178), .DIN1(N4055), .DIN2(N4114));
nor2s1 U1490 (.Q(N4179), .DIN1(N4114), .DIN2(N618));
nor2s1 U1491 (.Q(N4180), .DIN1(N3951), .DIN2(N4114));
nor2s1 U1492 (.Q(N4183), .DIN1(N4058), .DIN2(N4118));
nor2s1 U1493 (.Q(N4184), .DIN1(N4118), .DIN2(N666));
nor2s1 U1494 (.Q(N4185), .DIN1(N3955), .DIN2(N4118));
nor2s1 U1495 (.Q(N4188), .DIN1(N4061), .DIN2(N4122));
nor2s1 U1496 (.Q(N4189), .DIN1(N4122), .DIN2(N714));
nor2s1 U1497 (.Q(N4190), .DIN1(N3959), .DIN2(N4122));
nor2s1 U1498 (.Q(N4193), .DIN1(N4064), .DIN2(N4126));
nor2s1 U1499 (.Q(N4194), .DIN1(N4126), .DIN2(N762));
nor2s1 U1500 (.Q(N4195), .DIN1(N3963), .DIN2(N4126));
nor2s1 U1501 (.Q(N4198), .DIN1(N4067), .DIN2(N4130));
nor2s1 U1502 (.Q(N4199), .DIN1(N4130), .DIN2(N810));
nor2s1 U1503 (.Q(N4200), .DIN1(N3967), .DIN2(N4130));
nor2s1 U1504 (.Q(N4203), .DIN1(N4070), .DIN2(N4134));
nor2s1 U1505 (.Q(N4204), .DIN1(N4134), .DIN2(N858));
nor2s1 U1506 (.Q(N4205), .DIN1(N3971), .DIN2(N4134));
nor2s1 U1507 (.Q(N4208), .DIN1(N4138), .DIN2(N4139));
nor2s1 U1508 (.Q(N4211), .DIN1(N4143), .DIN2(N4140));
nor2s1 U1509 (.Q(N4215), .DIN1(N4082), .DIN2(N4146));
nor2s1 U1510 (.Q(N4216), .DIN1(N4146), .DIN2(N4079));
nor2s1 U1511 (.Q(N4217), .DIN1(N4150), .DIN2(N4151));
nor2s1 U1512 (.Q(N4220), .DIN1(N4152), .DIN2(N1053));
nor2s1 U1513 (.Q(N4224), .DIN1(N4091), .DIN2(N4155));
nor2s1 U1514 (.Q(N4225), .DIN1(N4155), .DIN2(N1101));
nor2s1 U1515 (.Q(N4226), .DIN1(N3992), .DIN2(N4155));
nor2s1 U1516 (.Q(N4229), .DIN1(N4159), .DIN2(N4160));
nor2s1 U1517 (.Q(N4232), .DIN1(N4164), .DIN2(N4161));
nor2s1 U1518 (.Q(N4236), .DIN1(N4103), .DIN2(N4167));
nor2s1 U1519 (.Q(N4237), .DIN1(N4167), .DIN2(N4100));
nor2s1 U1520 (.Q(N4238), .DIN1(N4171), .DIN2(N4172));
nor2s1 U1521 (.Q(N4241), .DIN1(N4173), .DIN2(N4174));
nor2s1 U1522 (.Q(N4242), .DIN1(N4178), .DIN2(N4179));
nor2s1 U1523 (.Q(N4245), .DIN1(N4183), .DIN2(N4184));
nor2s1 U1524 (.Q(N4248), .DIN1(N4188), .DIN2(N4189));
nor2s1 U1525 (.Q(N4251), .DIN1(N4193), .DIN2(N4194));
nor2s1 U1526 (.Q(N4254), .DIN1(N4198), .DIN2(N4199));
nor2s1 U1527 (.Q(N4257), .DIN1(N4203), .DIN2(N4204));
nor2s1 U1528 (.Q(N4260), .DIN1(N4208), .DIN2(N4205));
nor2s1 U1529 (.Q(N4264), .DIN1(N4143), .DIN2(N4211));
nor2s1 U1530 (.Q(N4265), .DIN1(N4211), .DIN2(N4140));
nor2s1 U1531 (.Q(N4266), .DIN1(N4215), .DIN2(N4216));
nor2s1 U1532 (.Q(N4269), .DIN1(N4217), .DIN2(N1005));
nor2s1 U1533 (.Q(N4273), .DIN1(N4152), .DIN2(N4220));
nor2s1 U1534 (.Q(N4274), .DIN1(N4220), .DIN2(N1053));
nor2s1 U1535 (.Q(N4275), .DIN1(N4034), .DIN2(N4220));
nor2s1 U1536 (.Q(N4278), .DIN1(N4224), .DIN2(N4225));
nor2s1 U1537 (.Q(N4281), .DIN1(N4229), .DIN2(N4226));
nor2s1 U1538 (.Q(N4285), .DIN1(N4164), .DIN2(N4232));
nor2s1 U1539 (.Q(N4286), .DIN1(N4232), .DIN2(N4161));
nor2s1 U1540 (.Q(N4287), .DIN1(N4236), .DIN2(N4237));
nor2s1 U1541 (.Q(N4290), .DIN1(N4238), .DIN2(N1248));
nor2s1 U1542 (.Q(N4294), .DIN1(N4242), .DIN2(N4175));
nor2s1 U1543 (.Q(N4298), .DIN1(N4245), .DIN2(N4180));
nor2s1 U1544 (.Q(N4302), .DIN1(N4248), .DIN2(N4185));
nor2s1 U1545 (.Q(N4306), .DIN1(N4251), .DIN2(N4190));
nor2s1 U1546 (.Q(N4310), .DIN1(N4254), .DIN2(N4195));
nor2s1 U1547 (.Q(N4314), .DIN1(N4257), .DIN2(N4200));
nor2s1 U1548 (.Q(N4318), .DIN1(N4208), .DIN2(N4260));
nor2s1 U1549 (.Q(N4319), .DIN1(N4260), .DIN2(N4205));
nor2s1 U1550 (.Q(N4320), .DIN1(N4264), .DIN2(N4265));
nor2s1 U1551 (.Q(N4323), .DIN1(N4266), .DIN2(N957));
nor2s1 U1552 (.Q(N4327), .DIN1(N4217), .DIN2(N4269));
nor2s1 U1553 (.Q(N4328), .DIN1(N4269), .DIN2(N1005));
nor2s1 U1554 (.Q(N4329), .DIN1(N4085), .DIN2(N4269));
nor2s1 U1555 (.Q(N4332), .DIN1(N4273), .DIN2(N4274));
nor2s1 U1556 (.Q(N4335), .DIN1(N4278), .DIN2(N4275));
nor2s1 U1557 (.Q(N4339), .DIN1(N4229), .DIN2(N4281));
nor2s1 U1558 (.Q(N4340), .DIN1(N4281), .DIN2(N4226));
nor2s1 U1559 (.Q(N4341), .DIN1(N4285), .DIN2(N4286));
nor2s1 U1560 (.Q(N4344), .DIN1(N4287), .DIN2(N1200));
nor2s1 U1561 (.Q(N4348), .DIN1(N4238), .DIN2(N4290));
nor2s1 U1562 (.Q(N4349), .DIN1(N4290), .DIN2(N1248));
nor2s1 U1563 (.Q(N4350), .DIN1(N4106), .DIN2(N4290));
nor2s1 U1564 (.Q(N4353), .DIN1(N4242), .DIN2(N4294));
nor2s1 U1565 (.Q(N4354), .DIN1(N4294), .DIN2(N4175));
nor2s1 U1566 (.Q(N4355), .DIN1(N4245), .DIN2(N4298));
nor2s1 U1567 (.Q(N4356), .DIN1(N4298), .DIN2(N4180));
nor2s1 U1568 (.Q(N4357), .DIN1(N4248), .DIN2(N4302));
nor2s1 U1569 (.Q(N4358), .DIN1(N4302), .DIN2(N4185));
nor2s1 U1570 (.Q(N4359), .DIN1(N4251), .DIN2(N4306));
nor2s1 U1571 (.Q(N4360), .DIN1(N4306), .DIN2(N4190));
nor2s1 U1572 (.Q(N4361), .DIN1(N4254), .DIN2(N4310));
nor2s1 U1573 (.Q(N4362), .DIN1(N4310), .DIN2(N4195));
nor2s1 U1574 (.Q(N4363), .DIN1(N4257), .DIN2(N4314));
nor2s1 U1575 (.Q(N4364), .DIN1(N4314), .DIN2(N4200));
nor2s1 U1576 (.Q(N4365), .DIN1(N4318), .DIN2(N4319));
nor2s1 U1577 (.Q(N4368), .DIN1(N4320), .DIN2(N909));
nor2s1 U1578 (.Q(N4372), .DIN1(N4266), .DIN2(N4323));
nor2s1 U1579 (.Q(N4373), .DIN1(N4323), .DIN2(N957));
nor2s1 U1580 (.Q(N4374), .DIN1(N4146), .DIN2(N4323));
nor2s1 U1581 (.Q(N4377), .DIN1(N4327), .DIN2(N4328));
nor2s1 U1582 (.Q(N4380), .DIN1(N4332), .DIN2(N4329));
nor2s1 U1583 (.Q(N4384), .DIN1(N4278), .DIN2(N4335));
nor2s1 U1584 (.Q(N4385), .DIN1(N4335), .DIN2(N4275));
nor2s1 U1585 (.Q(N4386), .DIN1(N4339), .DIN2(N4340));
nor2s1 U1586 (.Q(N4389), .DIN1(N4341), .DIN2(N1152));
nor2s1 U1587 (.Q(N4393), .DIN1(N4287), .DIN2(N4344));
nor2s1 U1588 (.Q(N4394), .DIN1(N4344), .DIN2(N1200));
nor2s1 U1589 (.Q(N4395), .DIN1(N4167), .DIN2(N4344));
nor2s1 U1590 (.Q(N4398), .DIN1(N4348), .DIN2(N4349));
nor2s1 U1591 (.Q(N4401), .DIN1(N1296), .DIN2(N4350));
nor2s1 U1592 (.Q(N4405), .DIN1(N4353), .DIN2(N4354));
nor2s1 U1593 (.Q(N4408), .DIN1(N4355), .DIN2(N4356));
nor2s1 U1594 (.Q(N4411), .DIN1(N4357), .DIN2(N4358));
nor2s1 U1595 (.Q(N4414), .DIN1(N4359), .DIN2(N4360));
nor2s1 U1596 (.Q(N4417), .DIN1(N4361), .DIN2(N4362));
nor2s1 U1597 (.Q(N4420), .DIN1(N4363), .DIN2(N4364));
nor2s1 U1598 (.Q(N4423), .DIN1(N4365), .DIN2(N861));
nor2s1 U1599 (.Q(N4427), .DIN1(N4320), .DIN2(N4368));
nor2s1 U1600 (.Q(N4428), .DIN1(N4368), .DIN2(N909));
nor2s1 U1601 (.Q(N4429), .DIN1(N4211), .DIN2(N4368));
nor2s1 U1602 (.Q(N4432), .DIN1(N4372), .DIN2(N4373));
nor2s1 U1603 (.Q(N4435), .DIN1(N4377), .DIN2(N4374));
nor2s1 U1604 (.Q(N4439), .DIN1(N4332), .DIN2(N4380));
nor2s1 U1605 (.Q(N4440), .DIN1(N4380), .DIN2(N4329));
nor2s1 U1606 (.Q(N4441), .DIN1(N4384), .DIN2(N4385));
nor2s1 U1607 (.Q(N4444), .DIN1(N4386), .DIN2(N1104));
nor2s1 U1608 (.Q(N4448), .DIN1(N4341), .DIN2(N4389));
nor2s1 U1609 (.Q(N4449), .DIN1(N4389), .DIN2(N1152));
nor2s1 U1610 (.Q(N4450), .DIN1(N4232), .DIN2(N4389));
nor2s1 U1611 (.Q(N4453), .DIN1(N4393), .DIN2(N4394));
nor2s1 U1612 (.Q(N4456), .DIN1(N4398), .DIN2(N4395));
nor2s1 U1613 (.Q(N4460), .DIN1(N1296), .DIN2(N4401));
nor2s1 U1614 (.Q(N4461), .DIN1(N4401), .DIN2(N4350));
nor2s1 U1615 (.Q(N4462), .DIN1(N4405), .DIN2(N573));
nor2s1 U1616 (.Q(N4466), .DIN1(N4408), .DIN2(N621));
nor2s1 U1617 (.Q(N4470), .DIN1(N4411), .DIN2(N669));
nor2s1 U1618 (.Q(N4474), .DIN1(N4414), .DIN2(N717));
nor2s1 U1619 (.Q(N4478), .DIN1(N4417), .DIN2(N765));
nor2s1 U1620 (.Q(N4482), .DIN1(N4420), .DIN2(N813));
nor2s1 U1621 (.Q(N4486), .DIN1(N4365), .DIN2(N4423));
nor2s1 U1622 (.Q(N4487), .DIN1(N4423), .DIN2(N861));
nor2s1 U1623 (.Q(N4488), .DIN1(N4260), .DIN2(N4423));
nor2s1 U1624 (.Q(N4491), .DIN1(N4427), .DIN2(N4428));
nor2s1 U1625 (.Q(N4494), .DIN1(N4432), .DIN2(N4429));
nor2s1 U1626 (.Q(N4498), .DIN1(N4377), .DIN2(N4435));
nor2s1 U1627 (.Q(N4499), .DIN1(N4435), .DIN2(N4374));
nor2s1 U1628 (.Q(N4500), .DIN1(N4439), .DIN2(N4440));
nor2s1 U1629 (.Q(N4503), .DIN1(N4441), .DIN2(N1056));
nor2s1 U1630 (.Q(N4507), .DIN1(N4386), .DIN2(N4444));
nor2s1 U1631 (.Q(N4508), .DIN1(N4444), .DIN2(N1104));
nor2s1 U1632 (.Q(N4509), .DIN1(N4281), .DIN2(N4444));
nor2s1 U1633 (.Q(N4512), .DIN1(N4448), .DIN2(N4449));
nor2s1 U1634 (.Q(N4515), .DIN1(N4453), .DIN2(N4450));
nor2s1 U1635 (.Q(N4519), .DIN1(N4398), .DIN2(N4456));
nor2s1 U1636 (.Q(N4520), .DIN1(N4456), .DIN2(N4395));
nor2s1 U1637 (.Q(N4521), .DIN1(N4460), .DIN2(N4461));
nor2s1 U1638 (.Q(N4524), .DIN1(N4405), .DIN2(N4462));
nor2s1 U1639 (.Q(N4525), .DIN1(N4462), .DIN2(N573));
nor2s1 U1640 (.Q(N4526), .DIN1(N4294), .DIN2(N4462));
nor2s1 U1641 (.Q(N4529), .DIN1(N4408), .DIN2(N4466));
nor2s1 U1642 (.Q(N4530), .DIN1(N4466), .DIN2(N621));
nor2s1 U1643 (.Q(N4531), .DIN1(N4298), .DIN2(N4466));
nor2s1 U1644 (.Q(N4534), .DIN1(N4411), .DIN2(N4470));
nor2s1 U1645 (.Q(N4535), .DIN1(N4470), .DIN2(N669));
nor2s1 U1646 (.Q(N4536), .DIN1(N4302), .DIN2(N4470));
nor2s1 U1647 (.Q(N4539), .DIN1(N4414), .DIN2(N4474));
nor2s1 U1648 (.Q(N4540), .DIN1(N4474), .DIN2(N717));
nor2s1 U1649 (.Q(N4541), .DIN1(N4306), .DIN2(N4474));
nor2s1 U1650 (.Q(N4544), .DIN1(N4417), .DIN2(N4478));
nor2s1 U1651 (.Q(N4545), .DIN1(N4478), .DIN2(N765));
nor2s1 U1652 (.Q(N4546), .DIN1(N4310), .DIN2(N4478));
nor2s1 U1653 (.Q(N4549), .DIN1(N4420), .DIN2(N4482));
nor2s1 U1654 (.Q(N4550), .DIN1(N4482), .DIN2(N813));
nor2s1 U1655 (.Q(N4551), .DIN1(N4314), .DIN2(N4482));
nor2s1 U1656 (.Q(N4554), .DIN1(N4486), .DIN2(N4487));
nor2s1 U1657 (.Q(N4557), .DIN1(N4491), .DIN2(N4488));
nor2s1 U1658 (.Q(N4561), .DIN1(N4432), .DIN2(N4494));
nor2s1 U1659 (.Q(N4562), .DIN1(N4494), .DIN2(N4429));
nor2s1 U1660 (.Q(N4563), .DIN1(N4498), .DIN2(N4499));
nor2s1 U1661 (.Q(N4566), .DIN1(N4500), .DIN2(N1008));
nor2s1 U1662 (.Q(N4570), .DIN1(N4441), .DIN2(N4503));
nor2s1 U1663 (.Q(N4571), .DIN1(N4503), .DIN2(N1056));
nor2s1 U1664 (.Q(N4572), .DIN1(N4335), .DIN2(N4503));
nor2s1 U1665 (.Q(N4575), .DIN1(N4507), .DIN2(N4508));
nor2s1 U1666 (.Q(N4578), .DIN1(N4512), .DIN2(N4509));
nor2s1 U1667 (.Q(N4582), .DIN1(N4453), .DIN2(N4515));
nor2s1 U1668 (.Q(N4583), .DIN1(N4515), .DIN2(N4450));
nor2s1 U1669 (.Q(N4584), .DIN1(N4519), .DIN2(N4520));
nor2s1 U1670 (.Q(N4587), .DIN1(N4521), .DIN2(N1251));
nor2s1 U1671 (.Q(N4591), .DIN1(N4524), .DIN2(N4525));
nor2s1 U1672 (.Q(N4592), .DIN1(N4529), .DIN2(N4530));
nor2s1 U1673 (.Q(N4595), .DIN1(N4534), .DIN2(N4535));
nor2s1 U1674 (.Q(N4598), .DIN1(N4539), .DIN2(N4540));
nor2s1 U1675 (.Q(N4601), .DIN1(N4544), .DIN2(N4545));
nor2s1 U1676 (.Q(N4604), .DIN1(N4549), .DIN2(N4550));
nor2s1 U1677 (.Q(N4607), .DIN1(N4554), .DIN2(N4551));
nor2s1 U1678 (.Q(N4611), .DIN1(N4491), .DIN2(N4557));
nor2s1 U1679 (.Q(N4612), .DIN1(N4557), .DIN2(N4488));
nor2s1 U1680 (.Q(N4613), .DIN1(N4561), .DIN2(N4562));
nor2s1 U1681 (.Q(N4616), .DIN1(N4563), .DIN2(N960));
nor2s1 U1682 (.Q(N4620), .DIN1(N4500), .DIN2(N4566));
nor2s1 U1683 (.Q(N4621), .DIN1(N4566), .DIN2(N1008));
nor2s1 U1684 (.Q(N4622), .DIN1(N4380), .DIN2(N4566));
nor2s1 U1685 (.Q(N4625), .DIN1(N4570), .DIN2(N4571));
nor2s1 U1686 (.Q(N4628), .DIN1(N4575), .DIN2(N4572));
nor2s1 U1687 (.Q(N4632), .DIN1(N4512), .DIN2(N4578));
nor2s1 U1688 (.Q(N4633), .DIN1(N4578), .DIN2(N4509));
nor2s1 U1689 (.Q(N4634), .DIN1(N4582), .DIN2(N4583));
nor2s1 U1690 (.Q(N4637), .DIN1(N4584), .DIN2(N1203));
nor2s1 U1691 (.Q(N4641), .DIN1(N4521), .DIN2(N4587));
nor2s1 U1692 (.Q(N4642), .DIN1(N4587), .DIN2(N1251));
nor2s1 U1693 (.Q(N4643), .DIN1(N4401), .DIN2(N4587));
nor2s1 U1694 (.Q(N4646), .DIN1(N4592), .DIN2(N4526));
nor2s1 U1695 (.Q(N4650), .DIN1(N4595), .DIN2(N4531));
nor2s1 U1696 (.Q(N4654), .DIN1(N4598), .DIN2(N4536));
nor2s1 U1697 (.Q(N4658), .DIN1(N4601), .DIN2(N4541));
nor2s1 U1698 (.Q(N4662), .DIN1(N4604), .DIN2(N4546));
nor2s1 U1699 (.Q(N4666), .DIN1(N4554), .DIN2(N4607));
nor2s1 U1700 (.Q(N4667), .DIN1(N4607), .DIN2(N4551));
nor2s1 U1701 (.Q(N4668), .DIN1(N4611), .DIN2(N4612));
nor2s1 U1702 (.Q(N4671), .DIN1(N4613), .DIN2(N912));
nor2s1 U1703 (.Q(N4675), .DIN1(N4563), .DIN2(N4616));
nor2s1 U1704 (.Q(N4676), .DIN1(N4616), .DIN2(N960));
nor2s1 U1705 (.Q(N4677), .DIN1(N4435), .DIN2(N4616));
nor2s1 U1706 (.Q(N4680), .DIN1(N4620), .DIN2(N4621));
nor2s1 U1707 (.Q(N4683), .DIN1(N4625), .DIN2(N4622));
nor2s1 U1708 (.Q(N4687), .DIN1(N4575), .DIN2(N4628));
nor2s1 U1709 (.Q(N4688), .DIN1(N4628), .DIN2(N4572));
nor2s1 U1710 (.Q(N4689), .DIN1(N4632), .DIN2(N4633));
nor2s1 U1711 (.Q(N4692), .DIN1(N4634), .DIN2(N1155));
nor2s1 U1712 (.Q(N4696), .DIN1(N4584), .DIN2(N4637));
nor2s1 U1713 (.Q(N4697), .DIN1(N4637), .DIN2(N1203));
nor2s1 U1714 (.Q(N4698), .DIN1(N4456), .DIN2(N4637));
nor2s1 U1715 (.Q(N4701), .DIN1(N4641), .DIN2(N4642));
nor2s1 U1716 (.Q(N4704), .DIN1(N1299), .DIN2(N4643));
nor2s1 U1717 (.Q(N4708), .DIN1(N4592), .DIN2(N4646));
nor2s1 U1718 (.Q(N4709), .DIN1(N4646), .DIN2(N4526));
nor2s1 U1719 (.Q(N4710), .DIN1(N4595), .DIN2(N4650));
nor2s1 U1720 (.Q(N4711), .DIN1(N4650), .DIN2(N4531));
nor2s1 U1721 (.Q(N4712), .DIN1(N4598), .DIN2(N4654));
nor2s1 U1722 (.Q(N4713), .DIN1(N4654), .DIN2(N4536));
nor2s1 U1723 (.Q(N4714), .DIN1(N4601), .DIN2(N4658));
nor2s1 U1724 (.Q(N4715), .DIN1(N4658), .DIN2(N4541));
nor2s1 U1725 (.Q(N4716), .DIN1(N4604), .DIN2(N4662));
nor2s1 U1726 (.Q(N4717), .DIN1(N4662), .DIN2(N4546));
nor2s1 U1727 (.Q(N4718), .DIN1(N4666), .DIN2(N4667));
nor2s1 U1728 (.Q(N4721), .DIN1(N4668), .DIN2(N864));
nor2s1 U1729 (.Q(N4725), .DIN1(N4613), .DIN2(N4671));
nor2s1 U1730 (.Q(N4726), .DIN1(N4671), .DIN2(N912));
nor2s1 U1731 (.Q(N4727), .DIN1(N4494), .DIN2(N4671));
nor2s1 U1732 (.Q(N4730), .DIN1(N4675), .DIN2(N4676));
nor2s1 U1733 (.Q(N4733), .DIN1(N4680), .DIN2(N4677));
nor2s1 U1734 (.Q(N4737), .DIN1(N4625), .DIN2(N4683));
nor2s1 U1735 (.Q(N4738), .DIN1(N4683), .DIN2(N4622));
nor2s1 U1736 (.Q(N4739), .DIN1(N4687), .DIN2(N4688));
nor2s1 U1737 (.Q(N4742), .DIN1(N4689), .DIN2(N1107));
nor2s1 U1738 (.Q(N4746), .DIN1(N4634), .DIN2(N4692));
nor2s1 U1739 (.Q(N4747), .DIN1(N4692), .DIN2(N1155));
nor2s1 U1740 (.Q(N4748), .DIN1(N4515), .DIN2(N4692));
nor2s1 U1741 (.Q(N4751), .DIN1(N4696), .DIN2(N4697));
nor2s1 U1742 (.Q(N4754), .DIN1(N4701), .DIN2(N4698));
nor2s1 U1743 (.Q(N4758), .DIN1(N1299), .DIN2(N4704));
nor2s1 U1744 (.Q(N4759), .DIN1(N4704), .DIN2(N4643));
nor2s1 U1745 (.Q(N4760), .DIN1(N4708), .DIN2(N4709));
nor2s1 U1746 (.Q(N4763), .DIN1(N4710), .DIN2(N4711));
nor2s1 U1747 (.Q(N4766), .DIN1(N4712), .DIN2(N4713));
nor2s1 U1748 (.Q(N4769), .DIN1(N4714), .DIN2(N4715));
nor2s1 U1749 (.Q(N4772), .DIN1(N4716), .DIN2(N4717));
nor2s1 U1750 (.Q(N4775), .DIN1(N4718), .DIN2(N816));
nor2s1 U1751 (.Q(N4779), .DIN1(N4668), .DIN2(N4721));
nor2s1 U1752 (.Q(N4780), .DIN1(N4721), .DIN2(N864));
nor2s1 U1753 (.Q(N4781), .DIN1(N4557), .DIN2(N4721));
nor2s1 U1754 (.Q(N4784), .DIN1(N4725), .DIN2(N4726));
nor2s1 U1755 (.Q(N4787), .DIN1(N4730), .DIN2(N4727));
nor2s1 U1756 (.Q(N4791), .DIN1(N4680), .DIN2(N4733));
nor2s1 U1757 (.Q(N4792), .DIN1(N4733), .DIN2(N4677));
nor2s1 U1758 (.Q(N4793), .DIN1(N4737), .DIN2(N4738));
nor2s1 U1759 (.Q(N4796), .DIN1(N4739), .DIN2(N1059));
nor2s1 U1760 (.Q(N4800), .DIN1(N4689), .DIN2(N4742));
nor2s1 U1761 (.Q(N4801), .DIN1(N4742), .DIN2(N1107));
nor2s1 U1762 (.Q(N4802), .DIN1(N4578), .DIN2(N4742));
nor2s1 U1763 (.Q(N4805), .DIN1(N4746), .DIN2(N4747));
nor2s1 U1764 (.Q(N4808), .DIN1(N4751), .DIN2(N4748));
nor2s1 U1765 (.Q(N4812), .DIN1(N4701), .DIN2(N4754));
nor2s1 U1766 (.Q(N4813), .DIN1(N4754), .DIN2(N4698));
nor2s1 U1767 (.Q(N4814), .DIN1(N4758), .DIN2(N4759));
nor2s1 U1768 (.Q(N4817), .DIN1(N4760), .DIN2(N576));
nor2s1 U1769 (.Q(N4821), .DIN1(N4763), .DIN2(N624));
nor2s1 U1770 (.Q(N4825), .DIN1(N4766), .DIN2(N672));
nor2s1 U1771 (.Q(N4829), .DIN1(N4769), .DIN2(N720));
nor2s1 U1772 (.Q(N4833), .DIN1(N4772), .DIN2(N768));
nor2s1 U1773 (.Q(N4837), .DIN1(N4718), .DIN2(N4775));
nor2s1 U1774 (.Q(N4838), .DIN1(N4775), .DIN2(N816));
nor2s1 U1775 (.Q(N4839), .DIN1(N4607), .DIN2(N4775));
nor2s1 U1776 (.Q(N4842), .DIN1(N4779), .DIN2(N4780));
nor2s1 U1777 (.Q(N4845), .DIN1(N4784), .DIN2(N4781));
nor2s1 U1778 (.Q(N4849), .DIN1(N4730), .DIN2(N4787));
nor2s1 U1779 (.Q(N4850), .DIN1(N4787), .DIN2(N4727));
nor2s1 U1780 (.Q(N4851), .DIN1(N4791), .DIN2(N4792));
nor2s1 U1781 (.Q(N4854), .DIN1(N4793), .DIN2(N1011));
nor2s1 U1782 (.Q(N4858), .DIN1(N4739), .DIN2(N4796));
nor2s1 U1783 (.Q(N4859), .DIN1(N4796), .DIN2(N1059));
nor2s1 U1784 (.Q(N4860), .DIN1(N4628), .DIN2(N4796));
nor2s1 U1785 (.Q(N4863), .DIN1(N4800), .DIN2(N4801));
nor2s1 U1786 (.Q(N4866), .DIN1(N4805), .DIN2(N4802));
nor2s1 U1787 (.Q(N4870), .DIN1(N4751), .DIN2(N4808));
nor2s1 U1788 (.Q(N4871), .DIN1(N4808), .DIN2(N4748));
nor2s1 U1789 (.Q(N4872), .DIN1(N4812), .DIN2(N4813));
nor2s1 U1790 (.Q(N4875), .DIN1(N4814), .DIN2(N1254));
nor2s1 U1791 (.Q(N4879), .DIN1(N4760), .DIN2(N4817));
nor2s1 U1792 (.Q(N4880), .DIN1(N4817), .DIN2(N576));
nor2s1 U1793 (.Q(N4881), .DIN1(N4646), .DIN2(N4817));
nor2s1 U1794 (.Q(N4884), .DIN1(N4763), .DIN2(N4821));
nor2s1 U1795 (.Q(N4885), .DIN1(N4821), .DIN2(N624));
nor2s1 U1796 (.Q(N4886), .DIN1(N4650), .DIN2(N4821));
nor2s1 U1797 (.Q(N4889), .DIN1(N4766), .DIN2(N4825));
nor2s1 U1798 (.Q(N4890), .DIN1(N4825), .DIN2(N672));
nor2s1 U1799 (.Q(N4891), .DIN1(N4654), .DIN2(N4825));
nor2s1 U1800 (.Q(N4894), .DIN1(N4769), .DIN2(N4829));
nor2s1 U1801 (.Q(N4895), .DIN1(N4829), .DIN2(N720));
nor2s1 U1802 (.Q(N4896), .DIN1(N4658), .DIN2(N4829));
nor2s1 U1803 (.Q(N4899), .DIN1(N4772), .DIN2(N4833));
nor2s1 U1804 (.Q(N4900), .DIN1(N4833), .DIN2(N768));
nor2s1 U1805 (.Q(N4901), .DIN1(N4662), .DIN2(N4833));
nor2s1 U1806 (.Q(N4904), .DIN1(N4837), .DIN2(N4838));
nor2s1 U1807 (.Q(N4907), .DIN1(N4842), .DIN2(N4839));
nor2s1 U1808 (.Q(N4911), .DIN1(N4784), .DIN2(N4845));
nor2s1 U1809 (.Q(N4912), .DIN1(N4845), .DIN2(N4781));
nor2s1 U1810 (.Q(N4913), .DIN1(N4849), .DIN2(N4850));
nor2s1 U1811 (.Q(N4916), .DIN1(N4851), .DIN2(N963));
nor2s1 U1812 (.Q(N4920), .DIN1(N4793), .DIN2(N4854));
nor2s1 U1813 (.Q(N4921), .DIN1(N4854), .DIN2(N1011));
nor2s1 U1814 (.Q(N4922), .DIN1(N4683), .DIN2(N4854));
nor2s1 U1815 (.Q(N4925), .DIN1(N4858), .DIN2(N4859));
nor2s1 U1816 (.Q(N4928), .DIN1(N4863), .DIN2(N4860));
nor2s1 U1817 (.Q(N4932), .DIN1(N4805), .DIN2(N4866));
nor2s1 U1818 (.Q(N4933), .DIN1(N4866), .DIN2(N4802));
nor2s1 U1819 (.Q(N4934), .DIN1(N4870), .DIN2(N4871));
nor2s1 U1820 (.Q(N4937), .DIN1(N4872), .DIN2(N1206));
nor2s1 U1821 (.Q(N4941), .DIN1(N4814), .DIN2(N4875));
nor2s1 U1822 (.Q(N4942), .DIN1(N4875), .DIN2(N1254));
nor2s1 U1823 (.Q(N4943), .DIN1(N4704), .DIN2(N4875));
nor2s1 U1824 (.Q(N4946), .DIN1(N4879), .DIN2(N4880));
nor2s1 U1825 (.Q(N4947), .DIN1(N4884), .DIN2(N4885));
nor2s1 U1826 (.Q(N4950), .DIN1(N4889), .DIN2(N4890));
nor2s1 U1827 (.Q(N4953), .DIN1(N4894), .DIN2(N4895));
nor2s1 U1828 (.Q(N4956), .DIN1(N4899), .DIN2(N4900));
nor2s1 U1829 (.Q(N4959), .DIN1(N4904), .DIN2(N4901));
nor2s1 U1830 (.Q(N4963), .DIN1(N4842), .DIN2(N4907));
nor2s1 U1831 (.Q(N4964), .DIN1(N4907), .DIN2(N4839));
nor2s1 U1832 (.Q(N4965), .DIN1(N4911), .DIN2(N4912));
nor2s1 U1833 (.Q(N4968), .DIN1(N4913), .DIN2(N915));
nor2s1 U1834 (.Q(N4972), .DIN1(N4851), .DIN2(N4916));
nor2s1 U1835 (.Q(N4973), .DIN1(N4916), .DIN2(N963));
nor2s1 U1836 (.Q(N4974), .DIN1(N4733), .DIN2(N4916));
nor2s1 U1837 (.Q(N4977), .DIN1(N4920), .DIN2(N4921));
nor2s1 U1838 (.Q(N4980), .DIN1(N4925), .DIN2(N4922));
nor2s1 U1839 (.Q(N4984), .DIN1(N4863), .DIN2(N4928));
nor2s1 U1840 (.Q(N4985), .DIN1(N4928), .DIN2(N4860));
nor2s1 U1841 (.Q(N4986), .DIN1(N4932), .DIN2(N4933));
nor2s1 U1842 (.Q(N4989), .DIN1(N4934), .DIN2(N1158));
nor2s1 U1843 (.Q(N4993), .DIN1(N4872), .DIN2(N4937));
nor2s1 U1844 (.Q(N4994), .DIN1(N4937), .DIN2(N1206));
nor2s1 U1845 (.Q(N4995), .DIN1(N4754), .DIN2(N4937));
nor2s1 U1846 (.Q(N4998), .DIN1(N4941), .DIN2(N4942));
nor2s1 U1847 (.Q(N5001), .DIN1(N1302), .DIN2(N4943));
nor2s1 U1848 (.Q(N5005), .DIN1(N4947), .DIN2(N4881));
nor2s1 U1849 (.Q(N5009), .DIN1(N4950), .DIN2(N4886));
nor2s1 U1850 (.Q(N5013), .DIN1(N4953), .DIN2(N4891));
nor2s1 U1851 (.Q(N5017), .DIN1(N4956), .DIN2(N4896));
nor2s1 U1852 (.Q(N5021), .DIN1(N4904), .DIN2(N4959));
nor2s1 U1853 (.Q(N5022), .DIN1(N4959), .DIN2(N4901));
nor2s1 U1854 (.Q(N5023), .DIN1(N4963), .DIN2(N4964));
nor2s1 U1855 (.Q(N5026), .DIN1(N4965), .DIN2(N867));
nor2s1 U1856 (.Q(N5030), .DIN1(N4913), .DIN2(N4968));
nor2s1 U1857 (.Q(N5031), .DIN1(N4968), .DIN2(N915));
nor2s1 U1858 (.Q(N5032), .DIN1(N4787), .DIN2(N4968));
nor2s1 U1859 (.Q(N5035), .DIN1(N4972), .DIN2(N4973));
nor2s1 U1860 (.Q(N5038), .DIN1(N4977), .DIN2(N4974));
nor2s1 U1861 (.Q(N5042), .DIN1(N4925), .DIN2(N4980));
nor2s1 U1862 (.Q(N5043), .DIN1(N4980), .DIN2(N4922));
nor2s1 U1863 (.Q(N5044), .DIN1(N4984), .DIN2(N4985));
nor2s1 U1864 (.Q(N5047), .DIN1(N4986), .DIN2(N1110));
nor2s1 U1865 (.Q(N5051), .DIN1(N4934), .DIN2(N4989));
nor2s1 U1866 (.Q(N5052), .DIN1(N4989), .DIN2(N1158));
nor2s1 U1867 (.Q(N5053), .DIN1(N4808), .DIN2(N4989));
nor2s1 U1868 (.Q(N5056), .DIN1(N4993), .DIN2(N4994));
nor2s1 U1869 (.Q(N5059), .DIN1(N4998), .DIN2(N4995));
nor2s1 U1870 (.Q(N5063), .DIN1(N1302), .DIN2(N5001));
nor2s1 U1871 (.Q(N5064), .DIN1(N5001), .DIN2(N4943));
nor2s1 U1872 (.Q(N5065), .DIN1(N4947), .DIN2(N5005));
nor2s1 U1873 (.Q(N5066), .DIN1(N5005), .DIN2(N4881));
nor2s1 U1874 (.Q(N5067), .DIN1(N4950), .DIN2(N5009));
nor2s1 U1875 (.Q(N5068), .DIN1(N5009), .DIN2(N4886));
nor2s1 U1876 (.Q(N5069), .DIN1(N4953), .DIN2(N5013));
nor2s1 U1877 (.Q(N5070), .DIN1(N5013), .DIN2(N4891));
nor2s1 U1878 (.Q(N5071), .DIN1(N4956), .DIN2(N5017));
nor2s1 U1879 (.Q(N5072), .DIN1(N5017), .DIN2(N4896));
nor2s1 U1880 (.Q(N5073), .DIN1(N5021), .DIN2(N5022));
nor2s1 U1881 (.Q(N5076), .DIN1(N5023), .DIN2(N819));
nor2s1 U1882 (.Q(N5080), .DIN1(N4965), .DIN2(N5026));
nor2s1 U1883 (.Q(N5081), .DIN1(N5026), .DIN2(N867));
nor2s1 U1884 (.Q(N5082), .DIN1(N4845), .DIN2(N5026));
nor2s1 U1885 (.Q(N5085), .DIN1(N5030), .DIN2(N5031));
nor2s1 U1886 (.Q(N5088), .DIN1(N5035), .DIN2(N5032));
nor2s1 U1887 (.Q(N5092), .DIN1(N4977), .DIN2(N5038));
nor2s1 U1888 (.Q(N5093), .DIN1(N5038), .DIN2(N4974));
nor2s1 U1889 (.Q(N5094), .DIN1(N5042), .DIN2(N5043));
nor2s1 U1890 (.Q(N5097), .DIN1(N5044), .DIN2(N1062));
nor2s1 U1891 (.Q(N5101), .DIN1(N4986), .DIN2(N5047));
nor2s1 U1892 (.Q(N5102), .DIN1(N5047), .DIN2(N1110));
nor2s1 U1893 (.Q(N5103), .DIN1(N4866), .DIN2(N5047));
nor2s1 U1894 (.Q(N5106), .DIN1(N5051), .DIN2(N5052));
nor2s1 U1895 (.Q(N5109), .DIN1(N5056), .DIN2(N5053));
nor2s1 U1896 (.Q(N5113), .DIN1(N4998), .DIN2(N5059));
nor2s1 U1897 (.Q(N5114), .DIN1(N5059), .DIN2(N4995));
nor2s1 U1898 (.Q(N5115), .DIN1(N5063), .DIN2(N5064));
nor2s1 U1899 (.Q(N5118), .DIN1(N5065), .DIN2(N5066));
nor2s1 U1900 (.Q(N5121), .DIN1(N5067), .DIN2(N5068));
nor2s1 U1901 (.Q(N5124), .DIN1(N5069), .DIN2(N5070));
nor2s1 U1902 (.Q(N5127), .DIN1(N5071), .DIN2(N5072));
nor2s1 U1903 (.Q(N5130), .DIN1(N5073), .DIN2(N771));
nor2s1 U1904 (.Q(N5134), .DIN1(N5023), .DIN2(N5076));
nor2s1 U1905 (.Q(N5135), .DIN1(N5076), .DIN2(N819));
nor2s1 U1906 (.Q(N5136), .DIN1(N4907), .DIN2(N5076));
nor2s1 U1907 (.Q(N5139), .DIN1(N5080), .DIN2(N5081));
nor2s1 U1908 (.Q(N5142), .DIN1(N5085), .DIN2(N5082));
nor2s1 U1909 (.Q(N5146), .DIN1(N5035), .DIN2(N5088));
nor2s1 U1910 (.Q(N5147), .DIN1(N5088), .DIN2(N5032));
nor2s1 U1911 (.Q(N5148), .DIN1(N5092), .DIN2(N5093));
nor2s1 U1912 (.Q(N5151), .DIN1(N5094), .DIN2(N1014));
nor2s1 U1913 (.Q(N5155), .DIN1(N5044), .DIN2(N5097));
nor2s1 U1914 (.Q(N5156), .DIN1(N5097), .DIN2(N1062));
nor2s1 U1915 (.Q(N5157), .DIN1(N4928), .DIN2(N5097));
nor2s1 U1916 (.Q(N5160), .DIN1(N5101), .DIN2(N5102));
nor2s1 U1917 (.Q(N5163), .DIN1(N5106), .DIN2(N5103));
nor2s1 U1918 (.Q(N5167), .DIN1(N5056), .DIN2(N5109));
nor2s1 U1919 (.Q(N5168), .DIN1(N5109), .DIN2(N5053));
nor2s1 U1920 (.Q(N5169), .DIN1(N5113), .DIN2(N5114));
nor2s1 U1921 (.Q(N5172), .DIN1(N5115), .DIN2(N1257));
nor2s1 U1922 (.Q(N5176), .DIN1(N5118), .DIN2(N579));
nor2s1 U1923 (.Q(N5180), .DIN1(N5121), .DIN2(N627));
nor2s1 U1924 (.Q(N5184), .DIN1(N5124), .DIN2(N675));
nor2s1 U1925 (.Q(N5188), .DIN1(N5127), .DIN2(N723));
nor2s1 U1926 (.Q(N5192), .DIN1(N5073), .DIN2(N5130));
nor2s1 U1927 (.Q(N5193), .DIN1(N5130), .DIN2(N771));
nor2s1 U1928 (.Q(N5194), .DIN1(N4959), .DIN2(N5130));
nor2s1 U1929 (.Q(N5197), .DIN1(N5134), .DIN2(N5135));
nor2s1 U1930 (.Q(N5200), .DIN1(N5139), .DIN2(N5136));
nor2s1 U1931 (.Q(N5204), .DIN1(N5085), .DIN2(N5142));
nor2s1 U1932 (.Q(N5205), .DIN1(N5142), .DIN2(N5082));
nor2s1 U1933 (.Q(N5206), .DIN1(N5146), .DIN2(N5147));
nor2s1 U1934 (.Q(N5209), .DIN1(N5148), .DIN2(N966));
nor2s1 U1935 (.Q(N5213), .DIN1(N5094), .DIN2(N5151));
nor2s1 U1936 (.Q(N5214), .DIN1(N5151), .DIN2(N1014));
nor2s1 U1937 (.Q(N5215), .DIN1(N4980), .DIN2(N5151));
nor2s1 U1938 (.Q(N5218), .DIN1(N5155), .DIN2(N5156));
nor2s1 U1939 (.Q(N5221), .DIN1(N5160), .DIN2(N5157));
nor2s1 U1940 (.Q(N5225), .DIN1(N5106), .DIN2(N5163));
nor2s1 U1941 (.Q(N5226), .DIN1(N5163), .DIN2(N5103));
nor2s1 U1942 (.Q(N5227), .DIN1(N5167), .DIN2(N5168));
nor2s1 U1943 (.Q(N5230), .DIN1(N5169), .DIN2(N1209));
nor2s1 U1944 (.Q(N5234), .DIN1(N5115), .DIN2(N5172));
nor2s1 U1945 (.Q(N5235), .DIN1(N5172), .DIN2(N1257));
nor2s1 U1946 (.Q(N5236), .DIN1(N5001), .DIN2(N5172));
nor2s1 U1947 (.Q(N5239), .DIN1(N5118), .DIN2(N5176));
nor2s1 U1948 (.Q(N5240), .DIN1(N5176), .DIN2(N579));
nor2s1 U1949 (.Q(N5241), .DIN1(N5005), .DIN2(N5176));
nor2s1 U1950 (.Q(N5244), .DIN1(N5121), .DIN2(N5180));
nor2s1 U1951 (.Q(N5245), .DIN1(N5180), .DIN2(N627));
nor2s1 U1952 (.Q(N5246), .DIN1(N5009), .DIN2(N5180));
nor2s1 U1953 (.Q(N5249), .DIN1(N5124), .DIN2(N5184));
nor2s1 U1954 (.Q(N5250), .DIN1(N5184), .DIN2(N675));
nor2s1 U1955 (.Q(N5251), .DIN1(N5013), .DIN2(N5184));
nor2s1 U1956 (.Q(N5254), .DIN1(N5127), .DIN2(N5188));
nor2s1 U1957 (.Q(N5255), .DIN1(N5188), .DIN2(N723));
nor2s1 U1958 (.Q(N5256), .DIN1(N5017), .DIN2(N5188));
nor2s1 U1959 (.Q(N5259), .DIN1(N5192), .DIN2(N5193));
nor2s1 U1960 (.Q(N5262), .DIN1(N5197), .DIN2(N5194));
nor2s1 U1961 (.Q(N5266), .DIN1(N5139), .DIN2(N5200));
nor2s1 U1962 (.Q(N5267), .DIN1(N5200), .DIN2(N5136));
nor2s1 U1963 (.Q(N5268), .DIN1(N5204), .DIN2(N5205));
nor2s1 U1964 (.Q(N5271), .DIN1(N5206), .DIN2(N918));
nor2s1 U1965 (.Q(N5275), .DIN1(N5148), .DIN2(N5209));
nor2s1 U1966 (.Q(N5276), .DIN1(N5209), .DIN2(N966));
nor2s1 U1967 (.Q(N5277), .DIN1(N5038), .DIN2(N5209));
nor2s1 U1968 (.Q(N5280), .DIN1(N5213), .DIN2(N5214));
nor2s1 U1969 (.Q(N5283), .DIN1(N5218), .DIN2(N5215));
nor2s1 U1970 (.Q(N5287), .DIN1(N5160), .DIN2(N5221));
nor2s1 U1971 (.Q(N5288), .DIN1(N5221), .DIN2(N5157));
nor2s1 U1972 (.Q(N5289), .DIN1(N5225), .DIN2(N5226));
nor2s1 U1973 (.Q(N5292), .DIN1(N5227), .DIN2(N1161));
nor2s1 U1974 (.Q(N5296), .DIN1(N5169), .DIN2(N5230));
nor2s1 U1975 (.Q(N5297), .DIN1(N5230), .DIN2(N1209));
nor2s1 U1976 (.Q(N5298), .DIN1(N5059), .DIN2(N5230));
nor2s1 U1977 (.Q(N5301), .DIN1(N5234), .DIN2(N5235));
nor2s1 U1978 (.Q(N5304), .DIN1(N1305), .DIN2(N5236));
nor2s1 U1979 (.Q(N5308), .DIN1(N5239), .DIN2(N5240));
nor2s1 U1980 (.Q(N5309), .DIN1(N5244), .DIN2(N5245));
nor2s1 U1981 (.Q(N5312), .DIN1(N5249), .DIN2(N5250));
nor2s1 U1982 (.Q(N5315), .DIN1(N5254), .DIN2(N5255));
nor2s1 U1983 (.Q(N5318), .DIN1(N5259), .DIN2(N5256));
nor2s1 U1984 (.Q(N5322), .DIN1(N5197), .DIN2(N5262));
nor2s1 U1985 (.Q(N5323), .DIN1(N5262), .DIN2(N5194));
nor2s1 U1986 (.Q(N5324), .DIN1(N5266), .DIN2(N5267));
nor2s1 U1987 (.Q(N5327), .DIN1(N5268), .DIN2(N870));
nor2s1 U1988 (.Q(N5331), .DIN1(N5206), .DIN2(N5271));
nor2s1 U1989 (.Q(N5332), .DIN1(N5271), .DIN2(N918));
nor2s1 U1990 (.Q(N5333), .DIN1(N5088), .DIN2(N5271));
nor2s1 U1991 (.Q(N5336), .DIN1(N5275), .DIN2(N5276));
nor2s1 U1992 (.Q(N5339), .DIN1(N5280), .DIN2(N5277));
nor2s1 U1993 (.Q(N5343), .DIN1(N5218), .DIN2(N5283));
nor2s1 U1994 (.Q(N5344), .DIN1(N5283), .DIN2(N5215));
nor2s1 U1995 (.Q(N5345), .DIN1(N5287), .DIN2(N5288));
nor2s1 U1996 (.Q(N5348), .DIN1(N5289), .DIN2(N1113));
nor2s1 U1997 (.Q(N5352), .DIN1(N5227), .DIN2(N5292));
nor2s1 U1998 (.Q(N5353), .DIN1(N5292), .DIN2(N1161));
nor2s1 U1999 (.Q(N5354), .DIN1(N5109), .DIN2(N5292));
nor2s1 U2000 (.Q(N5357), .DIN1(N5296), .DIN2(N5297));
nor2s1 U2001 (.Q(N5360), .DIN1(N5301), .DIN2(N5298));
nor2s1 U2002 (.Q(N5364), .DIN1(N1305), .DIN2(N5304));
nor2s1 U2003 (.Q(N5365), .DIN1(N5304), .DIN2(N5236));
nor2s1 U2004 (.Q(N5366), .DIN1(N5309), .DIN2(N5241));
nor2s1 U2005 (.Q(N5370), .DIN1(N5312), .DIN2(N5246));
nor2s1 U2006 (.Q(N5374), .DIN1(N5315), .DIN2(N5251));
nor2s1 U2007 (.Q(N5378), .DIN1(N5259), .DIN2(N5318));
nor2s1 U2008 (.Q(N5379), .DIN1(N5318), .DIN2(N5256));
nor2s1 U2009 (.Q(N5380), .DIN1(N5322), .DIN2(N5323));
nor2s1 U2010 (.Q(N5383), .DIN1(N5324), .DIN2(N822));
nor2s1 U2011 (.Q(N5387), .DIN1(N5268), .DIN2(N5327));
nor2s1 U2012 (.Q(N5388), .DIN1(N5327), .DIN2(N870));
nor2s1 U2013 (.Q(N5389), .DIN1(N5142), .DIN2(N5327));
nor2s1 U2014 (.Q(N5392), .DIN1(N5331), .DIN2(N5332));
nor2s1 U2015 (.Q(N5395), .DIN1(N5336), .DIN2(N5333));
nor2s1 U2016 (.Q(N5399), .DIN1(N5280), .DIN2(N5339));
nor2s1 U2017 (.Q(N5400), .DIN1(N5339), .DIN2(N5277));
nor2s1 U2018 (.Q(N5401), .DIN1(N5343), .DIN2(N5344));
nor2s1 U2019 (.Q(N5404), .DIN1(N5345), .DIN2(N1065));
nor2s1 U2020 (.Q(N5408), .DIN1(N5289), .DIN2(N5348));
nor2s1 U2021 (.Q(N5409), .DIN1(N5348), .DIN2(N1113));
nor2s1 U2022 (.Q(N5410), .DIN1(N5163), .DIN2(N5348));
nor2s1 U2023 (.Q(N5413), .DIN1(N5352), .DIN2(N5353));
nor2s1 U2024 (.Q(N5416), .DIN1(N5357), .DIN2(N5354));
nor2s1 U2025 (.Q(N5420), .DIN1(N5301), .DIN2(N5360));
nor2s1 U2026 (.Q(N5421), .DIN1(N5360), .DIN2(N5298));
nor2s1 U2027 (.Q(N5422), .DIN1(N5364), .DIN2(N5365));
nor2s1 U2028 (.Q(N5425), .DIN1(N5309), .DIN2(N5366));
nor2s1 U2029 (.Q(N5426), .DIN1(N5366), .DIN2(N5241));
nor2s1 U2030 (.Q(N5427), .DIN1(N5312), .DIN2(N5370));
nor2s1 U2031 (.Q(N5428), .DIN1(N5370), .DIN2(N5246));
nor2s1 U2032 (.Q(N5429), .DIN1(N5315), .DIN2(N5374));
nor2s1 U2033 (.Q(N5430), .DIN1(N5374), .DIN2(N5251));
nor2s1 U2034 (.Q(N5431), .DIN1(N5378), .DIN2(N5379));
nor2s1 U2035 (.Q(N5434), .DIN1(N5380), .DIN2(N774));
nor2s1 U2036 (.Q(N5438), .DIN1(N5324), .DIN2(N5383));
nor2s1 U2037 (.Q(N5439), .DIN1(N5383), .DIN2(N822));
nor2s1 U2038 (.Q(N5440), .DIN1(N5200), .DIN2(N5383));
nor2s1 U2039 (.Q(N5443), .DIN1(N5387), .DIN2(N5388));
nor2s1 U2040 (.Q(N5446), .DIN1(N5392), .DIN2(N5389));
nor2s1 U2041 (.Q(N5450), .DIN1(N5336), .DIN2(N5395));
nor2s1 U2042 (.Q(N5451), .DIN1(N5395), .DIN2(N5333));
nor2s1 U2043 (.Q(N5452), .DIN1(N5399), .DIN2(N5400));
nor2s1 U2044 (.Q(N5455), .DIN1(N5401), .DIN2(N1017));
nor2s1 U2045 (.Q(N5459), .DIN1(N5345), .DIN2(N5404));
nor2s1 U2046 (.Q(N5460), .DIN1(N5404), .DIN2(N1065));
nor2s1 U2047 (.Q(N5461), .DIN1(N5221), .DIN2(N5404));
nor2s1 U2048 (.Q(N5464), .DIN1(N5408), .DIN2(N5409));
nor2s1 U2049 (.Q(N5467), .DIN1(N5413), .DIN2(N5410));
nor2s1 U2050 (.Q(N5471), .DIN1(N5357), .DIN2(N5416));
nor2s1 U2051 (.Q(N5472), .DIN1(N5416), .DIN2(N5354));
nor2s1 U2052 (.Q(N5473), .DIN1(N5420), .DIN2(N5421));
nor2s1 U2053 (.Q(N5476), .DIN1(N5422), .DIN2(N1260));
nor2s1 U2054 (.Q(N5480), .DIN1(N5425), .DIN2(N5426));
nor2s1 U2055 (.Q(N5483), .DIN1(N5427), .DIN2(N5428));
nor2s1 U2056 (.Q(N5486), .DIN1(N5429), .DIN2(N5430));
nor2s1 U2057 (.Q(N5489), .DIN1(N5431), .DIN2(N726));
nor2s1 U2058 (.Q(N5493), .DIN1(N5380), .DIN2(N5434));
nor2s1 U2059 (.Q(N5494), .DIN1(N5434), .DIN2(N774));
nor2s1 U2060 (.Q(N5495), .DIN1(N5262), .DIN2(N5434));
nor2s1 U2061 (.Q(N5498), .DIN1(N5438), .DIN2(N5439));
nor2s1 U2062 (.Q(N5501), .DIN1(N5443), .DIN2(N5440));
nor2s1 U2063 (.Q(N5505), .DIN1(N5392), .DIN2(N5446));
nor2s1 U2064 (.Q(N5506), .DIN1(N5446), .DIN2(N5389));
nor2s1 U2065 (.Q(N5507), .DIN1(N5450), .DIN2(N5451));
nor2s1 U2066 (.Q(N5510), .DIN1(N5452), .DIN2(N969));
nor2s1 U2067 (.Q(N5514), .DIN1(N5401), .DIN2(N5455));
nor2s1 U2068 (.Q(N5515), .DIN1(N5455), .DIN2(N1017));
nor2s1 U2069 (.Q(N5516), .DIN1(N5283), .DIN2(N5455));
nor2s1 U2070 (.Q(N5519), .DIN1(N5459), .DIN2(N5460));
nor2s1 U2071 (.Q(N5522), .DIN1(N5464), .DIN2(N5461));
nor2s1 U2072 (.Q(N5526), .DIN1(N5413), .DIN2(N5467));
nor2s1 U2073 (.Q(N5527), .DIN1(N5467), .DIN2(N5410));
nor2s1 U2074 (.Q(N5528), .DIN1(N5471), .DIN2(N5472));
nor2s1 U2075 (.Q(N5531), .DIN1(N5473), .DIN2(N1212));
nor2s1 U2076 (.Q(N5535), .DIN1(N5422), .DIN2(N5476));
nor2s1 U2077 (.Q(N5536), .DIN1(N5476), .DIN2(N1260));
nor2s1 U2078 (.Q(N5537), .DIN1(N5304), .DIN2(N5476));
nor2s1 U2079 (.Q(N5540), .DIN1(N5480), .DIN2(N582));
nor2s1 U2080 (.Q(N5544), .DIN1(N5483), .DIN2(N630));
nor2s1 U2081 (.Q(N5548), .DIN1(N5486), .DIN2(N678));
nor2s1 U2082 (.Q(N5552), .DIN1(N5431), .DIN2(N5489));
nor2s1 U2083 (.Q(N5553), .DIN1(N5489), .DIN2(N726));
nor2s1 U2084 (.Q(N5554), .DIN1(N5318), .DIN2(N5489));
nor2s1 U2085 (.Q(N5557), .DIN1(N5493), .DIN2(N5494));
nor2s1 U2086 (.Q(N5560), .DIN1(N5498), .DIN2(N5495));
nor2s1 U2087 (.Q(N5564), .DIN1(N5443), .DIN2(N5501));
nor2s1 U2088 (.Q(N5565), .DIN1(N5501), .DIN2(N5440));
nor2s1 U2089 (.Q(N5566), .DIN1(N5505), .DIN2(N5506));
nor2s1 U2090 (.Q(N5569), .DIN1(N5507), .DIN2(N921));
nor2s1 U2091 (.Q(N5573), .DIN1(N5452), .DIN2(N5510));
nor2s1 U2092 (.Q(N5574), .DIN1(N5510), .DIN2(N969));
nor2s1 U2093 (.Q(N5575), .DIN1(N5339), .DIN2(N5510));
nor2s1 U2094 (.Q(N5578), .DIN1(N5514), .DIN2(N5515));
nor2s1 U2095 (.Q(N5581), .DIN1(N5519), .DIN2(N5516));
nor2s1 U2096 (.Q(N5585), .DIN1(N5464), .DIN2(N5522));
nor2s1 U2097 (.Q(N5586), .DIN1(N5522), .DIN2(N5461));
nor2s1 U2098 (.Q(N5587), .DIN1(N5526), .DIN2(N5527));
nor2s1 U2099 (.Q(N5590), .DIN1(N5528), .DIN2(N1164));
nor2s1 U2100 (.Q(N5594), .DIN1(N5473), .DIN2(N5531));
nor2s1 U2101 (.Q(N5595), .DIN1(N5531), .DIN2(N1212));
nor2s1 U2102 (.Q(N5596), .DIN1(N5360), .DIN2(N5531));
nor2s1 U2103 (.Q(N5599), .DIN1(N5535), .DIN2(N5536));
nor2s1 U2104 (.Q(N5602), .DIN1(N1308), .DIN2(N5537));
nor2s1 U2105 (.Q(N5606), .DIN1(N5480), .DIN2(N5540));
nor2s1 U2106 (.Q(N5607), .DIN1(N5540), .DIN2(N582));
nor2s1 U2107 (.Q(N5608), .DIN1(N5366), .DIN2(N5540));
nor2s1 U2108 (.Q(N5611), .DIN1(N5483), .DIN2(N5544));
nor2s1 U2109 (.Q(N5612), .DIN1(N5544), .DIN2(N630));
nor2s1 U2110 (.Q(N5613), .DIN1(N5370), .DIN2(N5544));
nor2s1 U2111 (.Q(N5616), .DIN1(N5486), .DIN2(N5548));
nor2s1 U2112 (.Q(N5617), .DIN1(N5548), .DIN2(N678));
nor2s1 U2113 (.Q(N5618), .DIN1(N5374), .DIN2(N5548));
nor2s1 U2114 (.Q(N5621), .DIN1(N5552), .DIN2(N5553));
nor2s1 U2115 (.Q(N5624), .DIN1(N5557), .DIN2(N5554));
nor2s1 U2116 (.Q(N5628), .DIN1(N5498), .DIN2(N5560));
nor2s1 U2117 (.Q(N5629), .DIN1(N5560), .DIN2(N5495));
nor2s1 U2118 (.Q(N5630), .DIN1(N5564), .DIN2(N5565));
nor2s1 U2119 (.Q(N5633), .DIN1(N5566), .DIN2(N873));
nor2s1 U2120 (.Q(N5637), .DIN1(N5507), .DIN2(N5569));
nor2s1 U2121 (.Q(N5638), .DIN1(N5569), .DIN2(N921));
nor2s1 U2122 (.Q(N5639), .DIN1(N5395), .DIN2(N5569));
nor2s1 U2123 (.Q(N5642), .DIN1(N5573), .DIN2(N5574));
nor2s1 U2124 (.Q(N5645), .DIN1(N5578), .DIN2(N5575));
nor2s1 U2125 (.Q(N5649), .DIN1(N5519), .DIN2(N5581));
nor2s1 U2126 (.Q(N5650), .DIN1(N5581), .DIN2(N5516));
nor2s1 U2127 (.Q(N5651), .DIN1(N5585), .DIN2(N5586));
nor2s1 U2128 (.Q(N5654), .DIN1(N5587), .DIN2(N1116));
nor2s1 U2129 (.Q(N5658), .DIN1(N5528), .DIN2(N5590));
nor2s1 U2130 (.Q(N5659), .DIN1(N5590), .DIN2(N1164));
nor2s1 U2131 (.Q(N5660), .DIN1(N5416), .DIN2(N5590));
nor2s1 U2132 (.Q(N5663), .DIN1(N5594), .DIN2(N5595));
nor2s1 U2133 (.Q(N5666), .DIN1(N5599), .DIN2(N5596));
nor2s1 U2134 (.Q(N5670), .DIN1(N1308), .DIN2(N5602));
nor2s1 U2135 (.Q(N5671), .DIN1(N5602), .DIN2(N5537));
nor2s1 U2136 (.Q(N5672), .DIN1(N5606), .DIN2(N5607));
nor2s1 U2137 (.Q(N5673), .DIN1(N5611), .DIN2(N5612));
nor2s1 U2138 (.Q(N5676), .DIN1(N5616), .DIN2(N5617));
nor2s1 U2139 (.Q(N5679), .DIN1(N5621), .DIN2(N5618));
nor2s1 U2140 (.Q(N5683), .DIN1(N5557), .DIN2(N5624));
nor2s1 U2141 (.Q(N5684), .DIN1(N5624), .DIN2(N5554));
nor2s1 U2142 (.Q(N5685), .DIN1(N5628), .DIN2(N5629));
nor2s1 U2143 (.Q(N5688), .DIN1(N5630), .DIN2(N825));
nor2s1 U2144 (.Q(N5692), .DIN1(N5566), .DIN2(N5633));
nor2s1 U2145 (.Q(N5693), .DIN1(N5633), .DIN2(N873));
nor2s1 U2146 (.Q(N5694), .DIN1(N5446), .DIN2(N5633));
nor2s1 U2147 (.Q(N5697), .DIN1(N5637), .DIN2(N5638));
nor2s1 U2148 (.Q(N5700), .DIN1(N5642), .DIN2(N5639));
nor2s1 U2149 (.Q(N5704), .DIN1(N5578), .DIN2(N5645));
nor2s1 U2150 (.Q(N5705), .DIN1(N5645), .DIN2(N5575));
nor2s1 U2151 (.Q(N5706), .DIN1(N5649), .DIN2(N5650));
nor2s1 U2152 (.Q(N5709), .DIN1(N5651), .DIN2(N1068));
nor2s1 U2153 (.Q(N5713), .DIN1(N5587), .DIN2(N5654));
nor2s1 U2154 (.Q(N5714), .DIN1(N5654), .DIN2(N1116));
nor2s1 U2155 (.Q(N5715), .DIN1(N5467), .DIN2(N5654));
nor2s1 U2156 (.Q(N5718), .DIN1(N5658), .DIN2(N5659));
nor2s1 U2157 (.Q(N5721), .DIN1(N5663), .DIN2(N5660));
nor2s1 U2158 (.Q(N5725), .DIN1(N5599), .DIN2(N5666));
nor2s1 U2159 (.Q(N5726), .DIN1(N5666), .DIN2(N5596));
nor2s1 U2160 (.Q(N5727), .DIN1(N5670), .DIN2(N5671));
nor2s1 U2161 (.Q(N5730), .DIN1(N5673), .DIN2(N5608));
nor2s1 U2162 (.Q(N5734), .DIN1(N5676), .DIN2(N5613));
nor2s1 U2163 (.Q(N5738), .DIN1(N5621), .DIN2(N5679));
nor2s1 U2164 (.Q(N5739), .DIN1(N5679), .DIN2(N5618));
nor2s1 U2165 (.Q(N5740), .DIN1(N5683), .DIN2(N5684));
nor2s1 U2166 (.Q(N5743), .DIN1(N5685), .DIN2(N777));
nor2s1 U2167 (.Q(N5747), .DIN1(N5630), .DIN2(N5688));
nor2s1 U2168 (.Q(N5748), .DIN1(N5688), .DIN2(N825));
nor2s1 U2169 (.Q(N5749), .DIN1(N5501), .DIN2(N5688));
nor2s1 U2170 (.Q(N5752), .DIN1(N5692), .DIN2(N5693));
nor2s1 U2171 (.Q(N5755), .DIN1(N5697), .DIN2(N5694));
nor2s1 U2172 (.Q(N5759), .DIN1(N5642), .DIN2(N5700));
nor2s1 U2173 (.Q(N5760), .DIN1(N5700), .DIN2(N5639));
nor2s1 U2174 (.Q(N5761), .DIN1(N5704), .DIN2(N5705));
nor2s1 U2175 (.Q(N5764), .DIN1(N5706), .DIN2(N1020));
nor2s1 U2176 (.Q(N5768), .DIN1(N5651), .DIN2(N5709));
nor2s1 U2177 (.Q(N5769), .DIN1(N5709), .DIN2(N1068));
nor2s1 U2178 (.Q(N5770), .DIN1(N5522), .DIN2(N5709));
nor2s1 U2179 (.Q(N5773), .DIN1(N5713), .DIN2(N5714));
nor2s1 U2180 (.Q(N5776), .DIN1(N5718), .DIN2(N5715));
nor2s1 U2181 (.Q(N5780), .DIN1(N5663), .DIN2(N5721));
nor2s1 U2182 (.Q(N5781), .DIN1(N5721), .DIN2(N5660));
nor2s1 U2183 (.Q(N5782), .DIN1(N5725), .DIN2(N5726));
nor2s1 U2184 (.Q(N5785), .DIN1(N5673), .DIN2(N5730));
nor2s1 U2185 (.Q(N5786), .DIN1(N5730), .DIN2(N5608));
nor2s1 U2186 (.Q(N5787), .DIN1(N5676), .DIN2(N5734));
nor2s1 U2187 (.Q(N5788), .DIN1(N5734), .DIN2(N5613));
nor2s1 U2188 (.Q(N5789), .DIN1(N5738), .DIN2(N5739));
nor2s1 U2189 (.Q(N5792), .DIN1(N5740), .DIN2(N729));
nor2s1 U2190 (.Q(N5796), .DIN1(N5685), .DIN2(N5743));
nor2s1 U2191 (.Q(N5797), .DIN1(N5743), .DIN2(N777));
nor2s1 U2192 (.Q(N5798), .DIN1(N5560), .DIN2(N5743));
nor2s1 U2193 (.Q(N5801), .DIN1(N5747), .DIN2(N5748));
nor2s1 U2194 (.Q(N5804), .DIN1(N5752), .DIN2(N5749));
nor2s1 U2195 (.Q(N5808), .DIN1(N5697), .DIN2(N5755));
nor2s1 U2196 (.Q(N5809), .DIN1(N5755), .DIN2(N5694));
nor2s1 U2197 (.Q(N5810), .DIN1(N5759), .DIN2(N5760));
nor2s1 U2198 (.Q(N5813), .DIN1(N5761), .DIN2(N972));
nor2s1 U2199 (.Q(N5817), .DIN1(N5706), .DIN2(N5764));
nor2s1 U2200 (.Q(N5818), .DIN1(N5764), .DIN2(N1020));
nor2s1 U2201 (.Q(N5819), .DIN1(N5581), .DIN2(N5764));
nor2s1 U2202 (.Q(N5822), .DIN1(N5768), .DIN2(N5769));
nor2s1 U2203 (.Q(N5825), .DIN1(N5773), .DIN2(N5770));
nor2s1 U2204 (.Q(N5829), .DIN1(N5718), .DIN2(N5776));
nor2s1 U2205 (.Q(N5830), .DIN1(N5776), .DIN2(N5715));
nor2s1 U2206 (.Q(N5831), .DIN1(N5780), .DIN2(N5781));
nor2s1 U2207 (.Q(N5834), .DIN1(N5785), .DIN2(N5786));
nor2s1 U2208 (.Q(N5837), .DIN1(N5787), .DIN2(N5788));
nor2s1 U2209 (.Q(N5840), .DIN1(N5789), .DIN2(N681));
nor2s1 U2210 (.Q(N5844), .DIN1(N5740), .DIN2(N5792));
nor2s1 U2211 (.Q(N5845), .DIN1(N5792), .DIN2(N729));
nor2s1 U2212 (.Q(N5846), .DIN1(N5624), .DIN2(N5792));
nor2s1 U2213 (.Q(N5849), .DIN1(N5796), .DIN2(N5797));
nor2s1 U2214 (.Q(N5852), .DIN1(N5801), .DIN2(N5798));
nor2s1 U2215 (.Q(N5856), .DIN1(N5752), .DIN2(N5804));
nor2s1 U2216 (.Q(N5857), .DIN1(N5804), .DIN2(N5749));
nor2s1 U2217 (.Q(N5858), .DIN1(N5808), .DIN2(N5809));
nor2s1 U2218 (.Q(N5861), .DIN1(N5810), .DIN2(N924));
nor2s1 U2219 (.Q(N5865), .DIN1(N5761), .DIN2(N5813));
nor2s1 U2220 (.Q(N5866), .DIN1(N5813), .DIN2(N972));
nor2s1 U2221 (.Q(N5867), .DIN1(N5645), .DIN2(N5813));
nor2s1 U2222 (.Q(N5870), .DIN1(N5817), .DIN2(N5818));
nor2s1 U2223 (.Q(N5873), .DIN1(N5822), .DIN2(N5819));
nor2s1 U2224 (.Q(N5877), .DIN1(N5773), .DIN2(N5825));
nor2s1 U2225 (.Q(N5878), .DIN1(N5825), .DIN2(N5770));
nor2s1 U2226 (.Q(N5879), .DIN1(N5829), .DIN2(N5830));
nor2s1 U2227 (.Q(N5882), .DIN1(N5834), .DIN2(N585));
nor2s1 U2228 (.Q(N5886), .DIN1(N5837), .DIN2(N633));
nor2s1 U2229 (.Q(N5890), .DIN1(N5789), .DIN2(N5840));
nor2s1 U2230 (.Q(N5891), .DIN1(N5840), .DIN2(N681));
nor2s1 U2231 (.Q(N5892), .DIN1(N5679), .DIN2(N5840));
nor2s1 U2232 (.Q(N5895), .DIN1(N5844), .DIN2(N5845));
nor2s1 U2233 (.Q(N5898), .DIN1(N5849), .DIN2(N5846));
nor2s1 U2234 (.Q(N5902), .DIN1(N5801), .DIN2(N5852));
nor2s1 U2235 (.Q(N5903), .DIN1(N5852), .DIN2(N5798));
nor2s1 U2236 (.Q(N5904), .DIN1(N5856), .DIN2(N5857));
nor2s1 U2237 (.Q(N5907), .DIN1(N5858), .DIN2(N876));
nor2s1 U2238 (.Q(N5911), .DIN1(N5810), .DIN2(N5861));
nor2s1 U2239 (.Q(N5912), .DIN1(N5861), .DIN2(N924));
nor2s1 U2240 (.Q(N5913), .DIN1(N5700), .DIN2(N5861));
nor2s1 U2241 (.Q(N5916), .DIN1(N5865), .DIN2(N5866));
nor2s1 U2242 (.Q(N5919), .DIN1(N5870), .DIN2(N5867));
nor2s1 U2243 (.Q(N5923), .DIN1(N5822), .DIN2(N5873));
nor2s1 U2244 (.Q(N5924), .DIN1(N5873), .DIN2(N5819));
nor2s1 U2245 (.Q(N5925), .DIN1(N5877), .DIN2(N5878));
nor2s1 U2246 (.Q(N5928), .DIN1(N5834), .DIN2(N5882));
nor2s1 U2247 (.Q(N5929), .DIN1(N5882), .DIN2(N585));
nor2s1 U2248 (.Q(N5930), .DIN1(N5730), .DIN2(N5882));
nor2s1 U2249 (.Q(N5933), .DIN1(N5837), .DIN2(N5886));
nor2s1 U2250 (.Q(N5934), .DIN1(N5886), .DIN2(N633));
nor2s1 U2251 (.Q(N5935), .DIN1(N5734), .DIN2(N5886));
nor2s1 U2252 (.Q(N5938), .DIN1(N5890), .DIN2(N5891));
nor2s1 U2253 (.Q(N5941), .DIN1(N5895), .DIN2(N5892));
nor2s1 U2254 (.Q(N5945), .DIN1(N5849), .DIN2(N5898));
nor2s1 U2255 (.Q(N5946), .DIN1(N5898), .DIN2(N5846));
nor2s1 U2256 (.Q(N5947), .DIN1(N5902), .DIN2(N5903));
nor2s1 U2257 (.Q(N5950), .DIN1(N5904), .DIN2(N828));
nor2s1 U2258 (.Q(N5954), .DIN1(N5858), .DIN2(N5907));
nor2s1 U2259 (.Q(N5955), .DIN1(N5907), .DIN2(N876));
nor2s1 U2260 (.Q(N5956), .DIN1(N5755), .DIN2(N5907));
nor2s1 U2261 (.Q(N5959), .DIN1(N5911), .DIN2(N5912));
nor2s1 U2262 (.Q(N5962), .DIN1(N5916), .DIN2(N5913));
nor2s1 U2263 (.Q(N5966), .DIN1(N5870), .DIN2(N5919));
nor2s1 U2264 (.Q(N5967), .DIN1(N5919), .DIN2(N5867));
nor2s1 U2265 (.Q(N5968), .DIN1(N5923), .DIN2(N5924));
nor2s1 U2266 (.Q(N5971), .DIN1(N5928), .DIN2(N5929));
nor2s1 U2267 (.Q(N5972), .DIN1(N5933), .DIN2(N5934));
nor2s1 U2268 (.Q(N5975), .DIN1(N5938), .DIN2(N5935));
nor2s1 U2269 (.Q(N5979), .DIN1(N5895), .DIN2(N5941));
nor2s1 U2270 (.Q(N5980), .DIN1(N5941), .DIN2(N5892));
nor2s1 U2271 (.Q(N5981), .DIN1(N5945), .DIN2(N5946));
nor2s1 U2272 (.Q(N5984), .DIN1(N5947), .DIN2(N780));
nor2s1 U2273 (.Q(N5988), .DIN1(N5904), .DIN2(N5950));
nor2s1 U2274 (.Q(N5989), .DIN1(N5950), .DIN2(N828));
nor2s1 U2275 (.Q(N5990), .DIN1(N5804), .DIN2(N5950));
nor2s1 U2276 (.Q(N5993), .DIN1(N5954), .DIN2(N5955));
nor2s1 U2277 (.Q(N5996), .DIN1(N5959), .DIN2(N5956));
nor2s1 U2278 (.Q(N6000), .DIN1(N5916), .DIN2(N5962));
nor2s1 U2279 (.Q(N6001), .DIN1(N5962), .DIN2(N5913));
nor2s1 U2280 (.Q(N6002), .DIN1(N5966), .DIN2(N5967));
nor2s1 U2281 (.Q(N6005), .DIN1(N5972), .DIN2(N5930));
nor2s1 U2282 (.Q(N6009), .DIN1(N5938), .DIN2(N5975));
nor2s1 U2283 (.Q(N6010), .DIN1(N5975), .DIN2(N5935));
nor2s1 U2284 (.Q(N6011), .DIN1(N5979), .DIN2(N5980));
nor2s1 U2285 (.Q(N6014), .DIN1(N5981), .DIN2(N732));
nor2s1 U2286 (.Q(N6018), .DIN1(N5947), .DIN2(N5984));
nor2s1 U2287 (.Q(N6019), .DIN1(N5984), .DIN2(N780));
nor2s1 U2288 (.Q(N6020), .DIN1(N5852), .DIN2(N5984));
nor2s1 U2289 (.Q(N6023), .DIN1(N5988), .DIN2(N5989));
nor2s1 U2290 (.Q(N6026), .DIN1(N5993), .DIN2(N5990));
nor2s1 U2291 (.Q(N6030), .DIN1(N5959), .DIN2(N5996));
nor2s1 U2292 (.Q(N6031), .DIN1(N5996), .DIN2(N5956));
nor2s1 U2293 (.Q(N6032), .DIN1(N6000), .DIN2(N6001));
nor2s1 U2294 (.Q(N6035), .DIN1(N5972), .DIN2(N6005));
nor2s1 U2295 (.Q(N6036), .DIN1(N6005), .DIN2(N5930));
nor2s1 U2296 (.Q(N6037), .DIN1(N6009), .DIN2(N6010));
nor2s1 U2297 (.Q(N6040), .DIN1(N6011), .DIN2(N684));
nor2s1 U2298 (.Q(N6044), .DIN1(N5981), .DIN2(N6014));
nor2s1 U2299 (.Q(N6045), .DIN1(N6014), .DIN2(N732));
nor2s1 U2300 (.Q(N6046), .DIN1(N5898), .DIN2(N6014));
nor2s1 U2301 (.Q(N6049), .DIN1(N6018), .DIN2(N6019));
nor2s1 U2302 (.Q(N6052), .DIN1(N6023), .DIN2(N6020));
nor2s1 U2303 (.Q(N6056), .DIN1(N5993), .DIN2(N6026));
nor2s1 U2304 (.Q(N6057), .DIN1(N6026), .DIN2(N5990));
nor2s1 U2305 (.Q(N6058), .DIN1(N6030), .DIN2(N6031));
nor2s1 U2306 (.Q(N6061), .DIN1(N6035), .DIN2(N6036));
nor2s1 U2307 (.Q(N6064), .DIN1(N6037), .DIN2(N636));
nor2s1 U2308 (.Q(N6068), .DIN1(N6011), .DIN2(N6040));
nor2s1 U2309 (.Q(N6069), .DIN1(N6040), .DIN2(N684));
nor2s1 U2310 (.Q(N6070), .DIN1(N5941), .DIN2(N6040));
nor2s1 U2311 (.Q(N6073), .DIN1(N6044), .DIN2(N6045));
nor2s1 U2312 (.Q(N6076), .DIN1(N6049), .DIN2(N6046));
nor2s1 U2313 (.Q(N6080), .DIN1(N6023), .DIN2(N6052));
nor2s1 U2314 (.Q(N6081), .DIN1(N6052), .DIN2(N6020));
nor2s1 U2315 (.Q(N6082), .DIN1(N6056), .DIN2(N6057));
nor2s1 U2316 (.Q(N6085), .DIN1(N6061), .DIN2(N588));
nor2s1 U2317 (.Q(N6089), .DIN1(N6037), .DIN2(N6064));
nor2s1 U2318 (.Q(N6090), .DIN1(N6064), .DIN2(N636));
nor2s1 U2319 (.Q(N6091), .DIN1(N5975), .DIN2(N6064));
nor2s1 U2320 (.Q(N6094), .DIN1(N6068), .DIN2(N6069));
nor2s1 U2321 (.Q(N6097), .DIN1(N6073), .DIN2(N6070));
nor2s1 U2322 (.Q(N6101), .DIN1(N6049), .DIN2(N6076));
nor2s1 U2323 (.Q(N6102), .DIN1(N6076), .DIN2(N6046));
nor2s1 U2324 (.Q(N6103), .DIN1(N6080), .DIN2(N6081));
nor2s1 U2325 (.Q(N6106), .DIN1(N6061), .DIN2(N6085));
nor2s1 U2326 (.Q(N6107), .DIN1(N6085), .DIN2(N588));
nor2s1 U2327 (.Q(N6108), .DIN1(N6005), .DIN2(N6085));
nor2s1 U2328 (.Q(N6111), .DIN1(N6089), .DIN2(N6090));
nor2s1 U2329 (.Q(N6114), .DIN1(N6094), .DIN2(N6091));
nor2s1 U2330 (.Q(N6118), .DIN1(N6073), .DIN2(N6097));
nor2s1 U2331 (.Q(N6119), .DIN1(N6097), .DIN2(N6070));
nor2s1 U2332 (.Q(N6120), .DIN1(N6101), .DIN2(N6102));
nor2s1 U2333 (.Q(N6123), .DIN1(N6106), .DIN2(N6107));
nor2s1 U2334 (.Q(N6124), .DIN1(N6111), .DIN2(N6108));
nor2s1 U2335 (.Q(N6128), .DIN1(N6094), .DIN2(N6114));
nor2s1 U2336 (.Q(N6129), .DIN1(N6114), .DIN2(N6091));
nor2s1 U2337 (.Q(N6130), .DIN1(N6118), .DIN2(N6119));
nor2s1 U2338 (.Q(N6133), .DIN1(N6111), .DIN2(N6124));
nor2s1 U2339 (.Q(N6134), .DIN1(N6124), .DIN2(N6108));
nor2s1 U2340 (.Q(N6135), .DIN1(N6128), .DIN2(N6129));
nor2s1 U2341 (.Q(N6138), .DIN1(N6133), .DIN2(N6134));
hi1s1 U2342 (.Q(N6141), .DIN(N6138));
nor2s1 U2343 (.Q(N6145), .DIN1(N6138), .DIN2(N6141));
hi1s1 U2344 (.Q(N6146), .DIN(N6141));
nor2s1 U2345 (.Q(N6147), .DIN1(N6124), .DIN2(N6141));
nor2s1 U2346 (.Q(N6150), .DIN1(N6145), .DIN2(N6146));
nor2s1 U2347 (.Q(N6151), .DIN1(N6135), .DIN2(N6147));
nor2s1 U2348 (.Q(N6155), .DIN1(N6135), .DIN2(N6151));
nor2s1 U2349 (.Q(N6156), .DIN1(N6151), .DIN2(N6147));
nor2s1 U2350 (.Q(N6157), .DIN1(N6114), .DIN2(N6151));
nor2s1 U2351 (.Q(N6160), .DIN1(N6155), .DIN2(N6156));
nor2s1 U2352 (.Q(N6161), .DIN1(N6130), .DIN2(N6157));
nor2s1 U2353 (.Q(N6165), .DIN1(N6130), .DIN2(N6161));
nor2s1 U2354 (.Q(N6166), .DIN1(N6161), .DIN2(N6157));
nor2s1 U2355 (.Q(N6167), .DIN1(N6097), .DIN2(N6161));
nor2s1 U2356 (.Q(N6170), .DIN1(N6165), .DIN2(N6166));
nor2s1 U2357 (.Q(N6171), .DIN1(N6120), .DIN2(N6167));
nor2s1 U2358 (.Q(N6175), .DIN1(N6120), .DIN2(N6171));
nor2s1 U2359 (.Q(N6176), .DIN1(N6171), .DIN2(N6167));
nor2s1 U2360 (.Q(N6177), .DIN1(N6076), .DIN2(N6171));
nor2s1 U2361 (.Q(N6180), .DIN1(N6175), .DIN2(N6176));
nor2s1 U2362 (.Q(N6181), .DIN1(N6103), .DIN2(N6177));
nor2s1 U2363 (.Q(N6185), .DIN1(N6103), .DIN2(N6181));
nor2s1 U2364 (.Q(N6186), .DIN1(N6181), .DIN2(N6177));
nor2s1 U2365 (.Q(N6187), .DIN1(N6052), .DIN2(N6181));
nor2s1 U2366 (.Q(N6190), .DIN1(N6185), .DIN2(N6186));
nor2s1 U2367 (.Q(N6191), .DIN1(N6082), .DIN2(N6187));
nor2s1 U2368 (.Q(N6195), .DIN1(N6082), .DIN2(N6191));
nor2s1 U2369 (.Q(N6196), .DIN1(N6191), .DIN2(N6187));
nor2s1 U2370 (.Q(N6197), .DIN1(N6026), .DIN2(N6191));
nor2s1 U2371 (.Q(N6200), .DIN1(N6195), .DIN2(N6196));
nor2s1 U2372 (.Q(N6201), .DIN1(N6058), .DIN2(N6197));
nor2s1 U2373 (.Q(N6205), .DIN1(N6058), .DIN2(N6201));
nor2s1 U2374 (.Q(N6206), .DIN1(N6201), .DIN2(N6197));
nor2s1 U2375 (.Q(N6207), .DIN1(N5996), .DIN2(N6201));
nor2s1 U2376 (.Q(N6210), .DIN1(N6205), .DIN2(N6206));
nor2s1 U2377 (.Q(N6211), .DIN1(N6032), .DIN2(N6207));
nor2s1 U2378 (.Q(N6215), .DIN1(N6032), .DIN2(N6211));
nor2s1 U2379 (.Q(N6216), .DIN1(N6211), .DIN2(N6207));
nor2s1 U2380 (.Q(N6217), .DIN1(N5962), .DIN2(N6211));
nor2s1 U2381 (.Q(N6220), .DIN1(N6215), .DIN2(N6216));
nor2s1 U2382 (.Q(N6221), .DIN1(N6002), .DIN2(N6217));
nor2s1 U2383 (.Q(N6225), .DIN1(N6002), .DIN2(N6221));
nor2s1 U2384 (.Q(N6226), .DIN1(N6221), .DIN2(N6217));
nor2s1 U2385 (.Q(N6227), .DIN1(N5919), .DIN2(N6221));
nor2s1 U2386 (.Q(N6230), .DIN1(N6225), .DIN2(N6226));
nor2s1 U2387 (.Q(N6231), .DIN1(N5968), .DIN2(N6227));
nor2s1 U2388 (.Q(N6235), .DIN1(N5968), .DIN2(N6231));
nor2s1 U2389 (.Q(N6236), .DIN1(N6231), .DIN2(N6227));
nor2s1 U2390 (.Q(N6237), .DIN1(N5873), .DIN2(N6231));
nor2s1 U2391 (.Q(N6240), .DIN1(N6235), .DIN2(N6236));
nor2s1 U2392 (.Q(N6241), .DIN1(N5925), .DIN2(N6237));
nor2s1 U2393 (.Q(N6245), .DIN1(N5925), .DIN2(N6241));
nor2s1 U2394 (.Q(N6246), .DIN1(N6241), .DIN2(N6237));
nor2s1 U2395 (.Q(N6247), .DIN1(N5825), .DIN2(N6241));
nor2s1 U2396 (.Q(N6250), .DIN1(N6245), .DIN2(N6246));
nor2s1 U2397 (.Q(N6251), .DIN1(N5879), .DIN2(N6247));
nor2s1 U2398 (.Q(N6255), .DIN1(N5879), .DIN2(N6251));
nor2s1 U2399 (.Q(N6256), .DIN1(N6251), .DIN2(N6247));
nor2s1 U2400 (.Q(N6257), .DIN1(N5776), .DIN2(N6251));
nor2s1 U2401 (.Q(N6260), .DIN1(N6255), .DIN2(N6256));
nor2s1 U2402 (.Q(N6261), .DIN1(N5831), .DIN2(N6257));
nor2s1 U2403 (.Q( tempN6265 ), .DIN1(N5831), .DIN2(N6261));
nor2s1 U2404 (.Q(N6266), .DIN1(N6261), .DIN2(N6257));
nor2s1 U2405 (.Q(N6267), .DIN1(N5721), .DIN2(N6261));
nor2s1 U2406 (.Q(N6270), .DIN1(N6265), .DIN2(N6266));
nor2s1 U2407 (.Q(N6271), .DIN1(N5782), .DIN2(N6267));
nor2s1 U2408 (.Q(N6275), .DIN1(N5782), .DIN2(N6271));
nor2s1 U2409 (.Q(N6276), .DIN1(N6271), .DIN2(N6267));
nor2s1 U2410 (.Q(N6277), .DIN1(N5666), .DIN2(N6271));
nor2s1 U2411 (.Q(N6280), .DIN1(N6275), .DIN2(N6276));
nor2s1 U2412 (.Q(N6281), .DIN1(N5727), .DIN2(N6277));
nor2s1 U2413 (.Q(N6285), .DIN1(N5727), .DIN2(N6281));
nor2s1 U2414 (.Q(N6286), .DIN1(N6281), .DIN2(N6277));
nor2s1 U2415 (.Q(N6287), .DIN1(N5602), .DIN2(N6281));
nor2s1 U2416 (.Q(N6288), .DIN1(N6285), .DIN2(N6286));
  nor2s1 troj65_0U1 ( .DIN1(troj65_0n1), .DIN2(troj65_0n2), .Q(Trigger_en65_0) );
  nnd4s1 troj65_0U2 ( .DIN1(N6128), .DIN2(N5038), .DIN3(N6205), .DIN4(troj65_0n3), .Q(troj65_0n2) );
  nor2s1 troj65_0U3 ( .DIN1(troj65_0n4), .DIN2(troj65_0n5), .Q(troj65_0n3) );
  nnd2s1 troj65_0U4 ( .DIN1(N5009), .DIN2(N4937), .Q(troj65_0n5) );
  nnd2s1 troj65_0U5 ( .DIN1(N4571), .DIN2(N4094), .Q(troj65_0n4) );
  nnd4s1 troj65_0U6 ( .DIN1(N2281), .DIN2(N2081), .DIN3(N3301), .DIN4(troj65_0n6), .Q(troj65_0n1) );
  nor3s1 troj65_0U7 ( .DIN1(troj65_0n7), .DIN2(N2545), .DIN3(troj65_0n8), .Q(troj65_0n6) );
  i1s1 troj65_0U8 ( .DIN(N1490), .Q(troj65_0n8) );
  nnd2s1 troj65_0U9 ( .DIN1(N1542), .DIN2(N1531), .Q(troj65_0n7) );
    xor2s1 trojan65_0  (.DIN1(tempN6265), .DIN2(Trigger_en65_0), .Q(N6265) );

endmodule
