
module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si, test_so );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so;
  wire   g2355, g4191, g4192, g4193, g4194, g4195, g4196, g4197, g4198, g4199,
         g4200, g4201, g4202, g4203, g4204, g4205, g4206, g4207, g4208, g4209,
         g4210, g4211, g4212, g4213, g4214, g4215, g4216, g4887, g4888, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g7744, g8061, g8062, g8271, g8561, g8562, g8563, g8564,
         g8565, g8566, g8984, g9961, n2061, n2074, g9930, n1975, n1982, g9895,
         n1948, n1983, g9827, n1980, g9826, n1953, g9825, g9824, g9823, g9822,
         g9821, g9820, n1978, n1987, g9819, g9818, n1985, g9356, n2008, g9355,
         n1993, n1954, g9354, g9353, n2028, n1932, n1957, g9352, g9351, g9350,
         n2010, n1956, n1935, g9349, g9348, n1989, g9347, n2009, g9346, n1994,
         n1955, g9345, g9344, n2029, n1933, n1958, g9343, g9342, g9341, n1968,
         n2039, n1936, g9340, g9339, g9338, n1981, g8993, g8992, g8991, g8990,
         g8989, g8988, g8987, g8874, n1974, g8873, n1976, n1929, g8872, g8871,
         n1949, g8870, g8869, g8868, g8782, g8781, g4190, g4187, g4186, g4189,
         g4188, g4185, g4184, g2613, g5656, g8780, g8695, g8694, g8573, g8572,
         n2045, g8571, n2046, g8570, n2007, g8569, n2047, \DFF_436/net723 ,
         g8568, n2043, g8567, n2055, g8450, g8449, g8448, g8447, g8446, g8445,
         g8444, g8443, g8442, g8441, g8440, g8439, g8438, n1991, g8437, g8436,
         g8435, g8434, g8433, g8432, g8431, g8430, g8429, g8428, g8427, n1937,
         g7750, g8426, n1992, g7752, g8425, n1959, g7753, g8424, g7754, g8423,
         g7755, g8422, n1960, g7756, g8421, n1996, g7757, g8420, n1961, g7758,
         g8419, n1938, g7759, g8418, g7751, g8288, g8287, g8286, g8285, g8284,
         g8283, g8282, g8281, g8280, n1952, g8279, g8278, g8277, g8276, g8274,
         n2049, g8273, n2056, g8272, n1925, n1926, g7749, n2017, n2023, n2034,
         n2018, n2035, n2019, n2036, n2020, n2037, n2021, n2038, n2022, g8080,
         g8079, g7329, g8078, g7335, g8077, g8076, g8067, g8066, g8065, g8064,
         g8063, n1951, g7817, g7816, g7815, g7814, g7813, n1984, g7812, g7811,
         g7810, g7809, \DFF_452/net739 , g7808, g7807, g7806, g7805, g7804,
         g7803, g7802, g7801, g7800, g7799, g7798, g7786, n2050, g7785, n2057,
         g7784, g7783, g7782, g7781, g7780, g7779, g7778, g7777, g7776, g7775,
         g7774, g7773, g7772, g7771, g7770, g7769, g7768, g7767, g7766, g7765,
         g7764, g7763, g7762, g7761, g7760, g7746, g7748, g7747, g7745, g7366,
         g7365, g7364, g7363, g7362, g7361, g7360, g7359, g7358, g7357, g7356,
         g7355, g7354, g7353, g7352, g7351, g7350, g7349, g7348, g7347, g7346,
         g7345, g7344, g7343, g7342, g7341, g7340, g7339, g7338, g7337, g7336,
         g7334, g7333, g7332, g7331, g7330, g7328, g7326, g7327, n2012, g7325,
         g7324, n1963, g7323, g7322, n1946, g7321, g6825, g7319, g7318, n2041,
         g7317, g7316, n2001, g7315, g7314, n1962, g7313, g7312, n1972, g7311,
         n2040, g7310, g7309, g7308, n1947, g7307, n1939, g7306, g7305, n2002,
         g7304, g6836, n1995, g7303, g7302, g7301, g7300, g7299, g7298, g7297,
         g7296, g7295, g7294, g7293, g7292, g7291, g7290, g7289, g7288, g7287,
         g7285, g6845, g6844, g4907, g6843, g4901, g6837, g6835, g6818, n2011,
         g6817, g6816, g6815, g6814, \DFF_126/net413 , g6813, g6812, g6811,
         g6810, g6809, g6808, g6807, g6806, g6805, g6804, g6803, g6802, g6800,
         n1990, n1999, g4183, g4182, g6801, g2639, g745, g6799, n2058, g6798,
         n2051, g6797, g6339, n2025, g6337, g6336, g1710, g6330, g6313, g6312,
         n1970, g6311, n1944, g6310, n2013, g6309, n1971, g6308, n1945, g6307,
         n2014, g6306, n2015, g6305, n2016, g6304, n1988, g6303, g6302, g6301,
         g6300, g6299, n1969, g5673, g4906, \DFF_489/net776 , g5671,
         \DFF_330/net617 , g5670, \DFF_385/net672 , g5669, g5668, g5667, g5666,
         g5665, g5664, g5663, g5662, g5661, g5660, g5657, g4894,
         \DFF_157/net444 , g632, g5655, \DFF_136/net423 , g5654,
         \DFF_336/net623 , \DFF_275/net562 , g4897, g4895, g3329, g1737,
         g11657, n2000, g4898, g11656, g11655, g11654, g11653, g11642, n1930,
         n1977, n1950, g11635, g11634, g11633, g11632, g11631, g11630, g11629,
         g11628, g11627, g1317, g11611, g11594, g11513, n2073, g11512, g11511,
         g11510, g11509, g11508, g11507, g11506, g11505, g11473, g11472, n2044,
         g11471, g11470, g11469, g11468, g11467, g11466, \DFF_441/net728 ,
         g11443, n2048, n2031, n2052, g11442, g11441, g11440, g11439, g11409,
         g10774, g11408, g2731, g5672, g1850, n1986, g11406, g11405, g11404,
         g11403, g11402, g11401, g11400, g11399, g11398, g11338, g11337,
         g11336, g11335, g11334, g11333, g11332, g11331, g11330, g11329,
         g11328, g11327, g11326, g11325, g11324, n2032, n2053, g11270, g11269,
         g11268, g11267, g11266, g11265, g11264, g11263, g11262, g11261,
         g11260, g11259, g11258, g11257, g11256, g11185, g11184, g11183,
         g11182, g11181, g11180, n2033, n2054, g11052, g11051, g11050, g11049,
         g11048, g11047, g11044, g11043, g11042, g11041, g11040, g11039,
         g11038, g11037, g11036, g11035, n1979, g11034, g11033, g10882, g10881,
         g10880, g10879, g10878, g10877, g10876, g10875, g10874, n2030,
         \DFF_194/net481 , g6846, g1765, g757, \DFF_121/net408 ,
         \DFF_93/net380 , g16, g37, g7, g17, g8, \DFF_228/net515 ,
         \DFF_242/net529 , \DFF_384/net671 , \DFF_319/net606 , g1360, g5645,
         g5647, g5648, g755, g5649, g874, g113, g875, g5643, g5646, g2044,
         g2638, g1217, g1955, g5644, g5652, g5650, g1356, g5651, g1956, g1736,
         n514, n516, n517, n518, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n872, n873, n874, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1927, n1928, n1931, n1934, n1940, n1941, n1942, n1943,
         n1964, n1965, n1966, n1967, n1973, n1997, n1998, n2003, n2004, n2005,
         n2006, n2024, n2026, n2027, n2042, n2059, n2060, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277;

wire Trojan_out0,  troj12_0counter_0_,  troj12_0N1,  troj12_0N2,  troj12_0N3,  troj12_0N6,  troj12_0n1,  troj12_0n2,  troj12_0n3,  troj12_0n4,  troj12_0n5,  troj12_0n6,  troj12_0n7,  troj12_0n8,  troj12_0n9,  troj12_0n10,  Trigger_en0_0,  trig50_0n1,  trig50_0n2,  trig50_0n3,  trig50_0n4,  trig50_0n5,  tempn1458;

  assign g11489 = 1'b0;
  assign g2355 = g18;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g4196 = g925;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g4204 = g922;
  assign g4205 = g1170;
  assign g4206 = g1197;
  assign g4207 = g1200;
  assign g4208 = g1203;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4887 = g1961;
  assign g4888 = g1960;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g6270 = g88;
  assign g6271 = g89;
  assign g6272 = g90;
  assign g6273 = g91;
  assign g6274 = g92;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g6285 = g28;
  assign g7744 = g27;
  assign g5101 = g8061;
  assign g8061 = g872;
  assign g5105 = g8062;
  assign g8062 = g873;
  assign g5816 = g8271;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign test_so = g8984;
  assign g9451 = g9961;

  xor2s3 U2 ( .DIN1(n907), .DIN2(n2575), .Q(n2826) );
  or3s3 U3 ( .DIN1(g6254), .DIN2(g6255), .DIN3(n908), .Q(g9961) );
  nor2s3 U4 ( .DIN1(n909), .DIN2(n2861), .Q(g9930) );
  xor2s3 U5 ( .DIN1(n910), .DIN2(n1975), .Q(n909) );
  nnd2s3 U6 ( .DIN1(n911), .DIN2(n912), .Q(n910) );
  nnd2s3 U7 ( .DIN1(n542), .DIN2(n913), .Q(n912) );
  nnd2s3 U8 ( .DIN1(n1982), .DIN2(n914), .Q(n913) );
  nnd2s3 U9 ( .DIN1(n662), .DIN2(n915), .Q(n914) );
  and3s3 U10 ( .DIN1(n916), .DIN2(n917), .DIN3(g2355), .Q(g9895) );
  nnd2s3 U11 ( .DIN1(n1948), .DIN2(n918), .Q(n917) );
  nnd3s3 U12 ( .DIN1(n919), .DIN2(n589), .DIN3(n920), .Q(n916) );
  nnd2s3 U13 ( .DIN1(n1983), .DIN2(n921), .Q(n919) );
  or2s3 U14 ( .DIN1(n922), .DIN2(n923), .Q(n921) );
  and3s3 U15 ( .DIN1(n924), .DIN2(n925), .DIN3(g2355), .Q(g9827) );
  nnd3s3 U16 ( .DIN1(n926), .DIN2(n927), .DIN3(n1980), .Q(n925) );
  or2s3 U17 ( .DIN1(n926), .DIN2(n1980), .Q(n924) );
  nnd3s3 U18 ( .DIN1(n928), .DIN2(n929), .DIN3(n923), .Q(n926) );
  nnd2s3 U19 ( .DIN1(n930), .DIN2(n702), .Q(n929) );
  nnd2s3 U20 ( .DIN1(n652), .DIN2(n698), .Q(n930) );
  nnd2s3 U21 ( .DIN1(n931), .DIN2(n652), .Q(n928) );
  nor2s3 U22 ( .DIN1(n2861), .DIN2(n932), .Q(g9826) );
  xor2s3 U23 ( .DIN1(n698), .DIN2(n933), .Q(n932) );
  nnd2s3 U24 ( .DIN1(n923), .DIN2(n934), .Q(n933) );
  nnd2s3 U25 ( .DIN1(n935), .DIN2(n936), .Q(n934) );
  nor2s3 U26 ( .DIN1(n2861), .DIN2(n937), .Q(g9825) );
  xor2s3 U27 ( .DIN1(n702), .DIN2(n938), .Q(n937) );
  nnd2s3 U28 ( .DIN1(n923), .DIN2(n939), .Q(n938) );
  nnd2s3 U29 ( .DIN1(n940), .DIN2(n922), .Q(n939) );
  nnd2s3 U30 ( .DIN1(n941), .DIN2(n942), .Q(n940) );
  nnd2s3 U31 ( .DIN1(n936), .DIN2(n702), .Q(n942) );
  nnd2s3 U32 ( .DIN1(n1986), .DIN2(n1953), .Q(n941) );
  nnd4s2 U33 ( .DIN1(n943), .DIN2(g6262), .DIN3(n897), .DIN4(n901), .Q(g9824)
         );
  nnd2s3 U34 ( .DIN1(n895), .DIN2(g6262), .Q(g9823) );
  nnd2s3 U35 ( .DIN1(n944), .DIN2(g6257), .Q(g9822) );
  nnd2s3 U36 ( .DIN1(n944), .DIN2(n897), .Q(g9821) );
  and3s3 U37 ( .DIN1(g6261), .DIN2(n902), .DIN3(n943), .Q(n944) );
  and3s3 U38 ( .DIN1(n945), .DIN2(n946), .DIN3(g2355), .Q(g9820) );
  nnd3s3 U39 ( .DIN1(n947), .DIN2(n948), .DIN3(n1978), .Q(n946) );
  nnd2s3 U40 ( .DIN1(n539), .DIN2(n949), .Q(n947) );
  nnd3s3 U41 ( .DIN1(n949), .DIN2(n660), .DIN3(n539), .Q(n945) );
  nnd3s3 U42 ( .DIN1(n950), .DIN2(n951), .DIN3(n952), .Q(n949) );
  nnd2s3 U43 ( .DIN1(n658), .DIN2(n691), .Q(n951) );
  nnd2s3 U44 ( .DIN1(n1987), .DIN2(n662), .Q(n950) );
  nor2s3 U45 ( .DIN1(n2861), .DIN2(n953), .Q(g9819) );
  xor2s3 U46 ( .DIN1(n691), .DIN2(n954), .Q(n953) );
  nnd2s3 U47 ( .DIN1(n539), .DIN2(n955), .Q(n954) );
  nnd2s3 U48 ( .DIN1(n956), .DIN2(n957), .Q(n955) );
  nnd2s3 U49 ( .DIN1(n958), .DIN2(n959), .Q(n956) );
  nnd2s3 U50 ( .DIN1(n1985), .DIN2(n960), .Q(n959) );
  nnd2s3 U51 ( .DIN1(n660), .DIN2(n691), .Q(n958) );
  nor2s3 U52 ( .DIN1(n2861), .DIN2(n961), .Q(g9818) );
  xor2s3 U53 ( .DIN1(n663), .DIN2(n962), .Q(n961) );
  nnd2s3 U54 ( .DIN1(n539), .DIN2(n963), .Q(n962) );
  nnd3s3 U55 ( .DIN1(n964), .DIN2(n965), .DIN3(n966), .Q(n963) );
  nnd2s3 U56 ( .DIN1(n658), .DIN2(n1985), .Q(n966) );
  nnd2s3 U57 ( .DIN1(n967), .DIN2(n968), .Q(g9356) );
  nnd2s3 U58 ( .DIN1(n969), .DIN2(n970), .Q(n968) );
  xor2s3 U59 ( .DIN1(n971), .DIN2(n2008), .Q(n969) );
  nnd3s3 U60 ( .DIN1(n972), .DIN2(n973), .DIN3(n974), .Q(n971) );
  nnd2s3 U61 ( .DIN1(n2502), .DIN2(n975), .Q(n974) );
  nnd3s3 U62 ( .DIN1(n976), .DIN2(n977), .DIN3(n586), .Q(n972) );
  nnd2s3 U63 ( .DIN1(n967), .DIN2(n978), .Q(g9355) );
  nnd2s3 U64 ( .DIN1(n979), .DIN2(n970), .Q(n978) );
  xor2s3 U65 ( .DIN1(n980), .DIN2(n1993), .Q(n979) );
  nnd3s3 U66 ( .DIN1(n981), .DIN2(n973), .DIN3(n982), .Q(n980) );
  nnd2s3 U67 ( .DIN1(n2503), .DIN2(n975), .Q(n982) );
  nnd3s3 U68 ( .DIN1(n983), .DIN2(n984), .DIN3(n586), .Q(n981) );
  nnd4s2 U69 ( .DIN1(n985), .DIN2(n849), .DIN3(n581), .DIN4(n699), .Q(n984) );
  nnd4s2 U70 ( .DIN1(n2028), .DIN2(n1957), .DIN3(n1954), .DIN4(n986), .Q(n983)
         );
  nnd2s3 U71 ( .DIN1(n967), .DIN2(n987), .Q(g9354) );
  nnd2s3 U72 ( .DIN1(n988), .DIN2(n970), .Q(n987) );
  xor2s3 U73 ( .DIN1(n989), .DIN2(n1954), .Q(n988) );
  nnd3s3 U74 ( .DIN1(n990), .DIN2(n973), .DIN3(n991), .Q(n989) );
  nnd2s3 U75 ( .DIN1(n2504), .DIN2(n975), .Q(n991) );
  nnd3s3 U76 ( .DIN1(n992), .DIN2(n993), .DIN3(n586), .Q(n990) );
  nnd3s3 U77 ( .DIN1(n581), .DIN2(n699), .DIN3(n985), .Q(n993) );
  nnd3s3 U78 ( .DIN1(n1957), .DIN2(n986), .DIN3(n2028), .Q(n992) );
  nnd2s3 U79 ( .DIN1(n967), .DIN2(n994), .Q(g9353) );
  nnd2s3 U80 ( .DIN1(n995), .DIN2(n970), .Q(n994) );
  xor2s3 U81 ( .DIN1(n996), .DIN2(n2028), .Q(n995) );
  nnd3s3 U82 ( .DIN1(n997), .DIN2(n973), .DIN3(n998), .Q(n996) );
  nnd2s3 U83 ( .DIN1(n2505), .DIN2(n975), .Q(n998) );
  nnd2s3 U84 ( .DIN1(n586), .DIN2(n999), .Q(n997) );
  nnd2s3 U85 ( .DIN1(n1000), .DIN2(n1001), .Q(n999) );
  nnd2s3 U86 ( .DIN1(n595), .DIN2(n581), .Q(n1001) );
  nnd2s3 U87 ( .DIN1(n1957), .DIN2(n596), .Q(n1000) );
  nnd2s3 U88 ( .DIN1(n967), .DIN2(n1002), .Q(g9352) );
  nnd2s3 U89 ( .DIN1(n1003), .DIN2(n970), .Q(n1002) );
  xor2s3 U90 ( .DIN1(n1004), .DIN2(n1957), .Q(n1003) );
  nnd3s3 U91 ( .DIN1(n1005), .DIN2(n973), .DIN3(n1006), .Q(n1004) );
  nnd2s3 U92 ( .DIN1(n2506), .DIN2(n975), .Q(n1006) );
  nnd2s3 U93 ( .DIN1(n586), .DIN2(n1007), .Q(n1005) );
  nnd2s3 U94 ( .DIN1(n1008), .DIN2(n1009), .Q(n1007) );
  nnd2s3 U95 ( .DIN1(n1010), .DIN2(n675), .Q(n1009) );
  nnd2s3 U96 ( .DIN1(n1932), .DIN2(n1011), .Q(n1008) );
  nnd2s3 U97 ( .DIN1(n967), .DIN2(n1012), .Q(g9351) );
  nnd2s3 U98 ( .DIN1(n1013), .DIN2(n970), .Q(n1012) );
  xor2s3 U99 ( .DIN1(n1014), .DIN2(n1932), .Q(n1013) );
  nnd3s3 U100 ( .DIN1(n1015), .DIN2(n973), .DIN3(n1016), .Q(n1014) );
  nnd2s3 U101 ( .DIN1(n2507), .DIN2(n975), .Q(n1016) );
  nnd3s3 U102 ( .DIN1(n1010), .DIN2(n1011), .DIN3(n586), .Q(n1015) );
  nnd2s3 U103 ( .DIN1(n967), .DIN2(n1017), .Q(g9350) );
  nnd2s3 U104 ( .DIN1(n1018), .DIN2(n970), .Q(n1017) );
  xor2s3 U105 ( .DIN1(n1019), .DIN2(n2010), .Q(n1018) );
  nnd3s3 U106 ( .DIN1(n1020), .DIN2(n973), .DIN3(n1021), .Q(n1019) );
  nnd2s3 U107 ( .DIN1(n2508), .DIN2(n975), .Q(n1021) );
  nnd2s3 U108 ( .DIN1(n586), .DIN2(n1022), .Q(n1020) );
  nnd3s3 U109 ( .DIN1(n1023), .DIN2(n1024), .DIN3(n1025), .Q(n1022) );
  or2s3 U110 ( .DIN1(n594), .DIN2(n1935), .Q(n1025) );
  nnd2s3 U111 ( .DIN1(n651), .DIN2(n594), .Q(n1024) );
  nnd2s3 U112 ( .DIN1(n1935), .DIN2(n1026), .Q(n1023) );
  nnd2s3 U113 ( .DIN1(n967), .DIN2(n1027), .Q(g9349) );
  nnd2s3 U114 ( .DIN1(n1028), .DIN2(n970), .Q(n1027) );
  xor2s3 U115 ( .DIN1(n1029), .DIN2(n1935), .Q(n1028) );
  nnd3s3 U116 ( .DIN1(n1030), .DIN2(n973), .DIN3(n1031), .Q(n1029) );
  nnd2s3 U117 ( .DIN1(n2509), .DIN2(n975), .Q(n1031) );
  nnd2s3 U118 ( .DIN1(n586), .DIN2(n1032), .Q(n1030) );
  xor2s3 U119 ( .DIN1(n594), .DIN2(n1026), .Q(n1032) );
  nnd2s3 U120 ( .DIN1(n967), .DIN2(n1033), .Q(g9348) );
  nnd2s3 U121 ( .DIN1(n1034), .DIN2(n970), .Q(n1033) );
  xor2s3 U122 ( .DIN1(n1035), .DIN2(n1956), .Q(n1034) );
  nnd2s3 U123 ( .DIN1(n973), .DIN2(n1036), .Q(n1035) );
  nnd2s3 U124 ( .DIN1(n2510), .DIN2(n975), .Q(n1036) );
  nnd2s3 U125 ( .DIN1(n586), .DIN2(n1037), .Q(n973) );
  nnd2s3 U126 ( .DIN1(n1038), .DIN2(n918), .Q(n975) );
  nnd2s3 U127 ( .DIN1(n920), .DIN2(n747), .Q(n918) );
  nor2s3 U129 ( .DIN1(n591), .DIN2(n923), .Q(n970) );
  and3s3 U130 ( .DIN1(n1039), .DIN2(n1040), .DIN3(n588), .Q(n923) );
  nnd2s3 U131 ( .DIN1(n920), .DIN2(n1041), .Q(n1037) );
  nnd2s3 U132 ( .DIN1(n1042), .DIN2(n922), .Q(n1041) );
  or2s3 U133 ( .DIN1(n1989), .DIN2(n1043), .Q(n1042) );
  nnd2s3 U134 ( .DIN1(n976), .DIN2(n721), .Q(n1040) );
  or5s3 U135 ( .DIN1(n2028), .DIN2(n1993), .DIN3(n1957), .DIN4(n1954), .DIN5(
        n595), .Q(n976) );
  nor2s3 U136 ( .DIN1(n1010), .DIN2(n1932), .Q(n985) );
  or4s3 U137 ( .DIN1(n651), .DIN2(n1935), .DIN3(n1956), .DIN4(n2010), .Q(n1010) );
  nnd2s3 U138 ( .DIN1(n2008), .DIN2(n977), .Q(n1039) );
  or5s3 U139 ( .DIN1(n596), .DIN2(n849), .DIN3(n581), .DIN4(n752), .DIN5(n699), 
        .Q(n977) );
  nor2s3 U140 ( .DIN1(n675), .DIN2(n1011), .Q(n986) );
  nnd4s2 U141 ( .DIN1(n2010), .DIN2(n1956), .DIN3(n1935), .DIN4(n651), .Q(
        n1011) );
  nnd2s3 U142 ( .DIN1(n698), .DIN2(n1044), .Q(n1026) );
  nnd2s3 U143 ( .DIN1(n1986), .DIN2(n1980), .Q(n1044) );
  nnd3s3 U144 ( .DIN1(n589), .DIN2(n702), .DIN3(n1983), .Q(n922) );
  nnd2s3 U145 ( .DIN1(n1045), .DIN2(n1046), .Q(g9347) );
  nnd2s3 U146 ( .DIN1(n1047), .DIN2(n540), .Q(n1046) );
  xor2s3 U147 ( .DIN1(n1048), .DIN2(n2009), .Q(n1047) );
  nnd3s3 U148 ( .DIN1(n1049), .DIN2(n1050), .DIN3(n1051), .Q(n1048) );
  nnd2s3 U149 ( .DIN1(n2493), .DIN2(n1052), .Q(n1051) );
  nnd3s3 U150 ( .DIN1(n1053), .DIN2(n1054), .DIN3(n538), .Q(n1049) );
  nnd2s3 U151 ( .DIN1(n1045), .DIN2(n1055), .Q(g9346) );
  nnd2s3 U152 ( .DIN1(n1056), .DIN2(n540), .Q(n1055) );
  xor2s3 U153 ( .DIN1(n1057), .DIN2(n1994), .Q(n1056) );
  nnd3s3 U154 ( .DIN1(n1058), .DIN2(n1050), .DIN3(n1059), .Q(n1057) );
  nnd2s3 U155 ( .DIN1(n2494), .DIN2(n1052), .Q(n1059) );
  nnd3s3 U156 ( .DIN1(n1060), .DIN2(n1061), .DIN3(n538), .Q(n1058) );
  nnd4s2 U157 ( .DIN1(n1062), .DIN2(n867), .DIN3(n866), .DIN4(n838), .Q(n1061)
         );
  nnd4s2 U158 ( .DIN1(n2029), .DIN2(n1958), .DIN3(n1955), .DIN4(n1063), .Q(
        n1060) );
  nnd2s3 U159 ( .DIN1(n1045), .DIN2(n1064), .Q(g9345) );
  nnd2s3 U160 ( .DIN1(n1065), .DIN2(n540), .Q(n1064) );
  xor2s3 U161 ( .DIN1(n1066), .DIN2(n1955), .Q(n1065) );
  nnd3s3 U162 ( .DIN1(n1067), .DIN2(n1050), .DIN3(n1068), .Q(n1066) );
  nnd2s3 U163 ( .DIN1(n2495), .DIN2(n1052), .Q(n1068) );
  nnd3s3 U164 ( .DIN1(n1069), .DIN2(n1070), .DIN3(n538), .Q(n1067) );
  nnd3s3 U165 ( .DIN1(n866), .DIN2(n838), .DIN3(n1062), .Q(n1070) );
  nnd3s3 U166 ( .DIN1(n1958), .DIN2(n1063), .DIN3(n2029), .Q(n1069) );
  nnd2s3 U167 ( .DIN1(n1045), .DIN2(n1071), .Q(g9344) );
  nnd2s3 U168 ( .DIN1(n1072), .DIN2(n540), .Q(n1071) );
  xor2s3 U169 ( .DIN1(n1073), .DIN2(n2029), .Q(n1072) );
  nnd3s3 U170 ( .DIN1(n1074), .DIN2(n1050), .DIN3(n1075), .Q(n1073) );
  nnd2s3 U171 ( .DIN1(n2496), .DIN2(n1052), .Q(n1075) );
  nnd2s3 U172 ( .DIN1(n538), .DIN2(n1076), .Q(n1074) );
  nnd2s3 U173 ( .DIN1(n1077), .DIN2(n1078), .Q(n1076) );
  nnd2s3 U174 ( .DIN1(n592), .DIN2(n866), .Q(n1078) );
  nnd2s3 U175 ( .DIN1(n1958), .DIN2(n593), .Q(n1077) );
  nnd2s3 U176 ( .DIN1(n1045), .DIN2(n1079), .Q(g9343) );
  nnd2s3 U177 ( .DIN1(n1080), .DIN2(n540), .Q(n1079) );
  xor2s3 U178 ( .DIN1(n1081), .DIN2(n1958), .Q(n1080) );
  nnd3s3 U179 ( .DIN1(n1082), .DIN2(n1050), .DIN3(n1083), .Q(n1081) );
  nnd2s3 U180 ( .DIN1(n2497), .DIN2(n1052), .Q(n1083) );
  nnd2s3 U181 ( .DIN1(n538), .DIN2(n1084), .Q(n1082) );
  nnd2s3 U182 ( .DIN1(n1085), .DIN2(n1086), .Q(n1084) );
  nnd2s3 U183 ( .DIN1(n1087), .DIN2(n687), .Q(n1086) );
  nnd2s3 U184 ( .DIN1(n1933), .DIN2(n1088), .Q(n1085) );
  nnd2s3 U185 ( .DIN1(n1045), .DIN2(n1089), .Q(g9342) );
  nnd2s3 U186 ( .DIN1(n1090), .DIN2(n540), .Q(n1089) );
  xor2s3 U187 ( .DIN1(n1091), .DIN2(n1933), .Q(n1090) );
  nnd3s3 U188 ( .DIN1(n1092), .DIN2(n1050), .DIN3(n1093), .Q(n1091) );
  nnd2s3 U189 ( .DIN1(n2498), .DIN2(n1052), .Q(n1093) );
  nnd3s3 U190 ( .DIN1(n1087), .DIN2(n1088), .DIN3(n538), .Q(n1092) );
  nnd2s3 U191 ( .DIN1(n1045), .DIN2(n1094), .Q(g9341) );
  nnd2s3 U192 ( .DIN1(n1095), .DIN2(n540), .Q(n1094) );
  xor2s3 U193 ( .DIN1(n1096), .DIN2(n1968), .Q(n1095) );
  nnd3s3 U194 ( .DIN1(n1097), .DIN2(n1050), .DIN3(n1098), .Q(n1096) );
  nnd2s3 U195 ( .DIN1(n2499), .DIN2(n1052), .Q(n1098) );
  nnd2s3 U196 ( .DIN1(n538), .DIN2(n1099), .Q(n1097) );
  nnd3s3 U197 ( .DIN1(n1100), .DIN2(n1101), .DIN3(n1102), .Q(n1099) );
  nnd2s3 U198 ( .DIN1(n2039), .DIN2(n638), .Q(n1102) );
  or2s3 U199 ( .DIN1(n1103), .DIN2(n2039), .Q(n1101) );
  nnd2s3 U200 ( .DIN1(n1936), .DIN2(n1103), .Q(n1100) );
  nnd2s3 U201 ( .DIN1(n1045), .DIN2(n1104), .Q(g9340) );
  nnd2s3 U202 ( .DIN1(n1105), .DIN2(n540), .Q(n1104) );
  xor2s3 U203 ( .DIN1(n1106), .DIN2(n1936), .Q(n1105) );
  nnd3s3 U204 ( .DIN1(n1107), .DIN2(n1050), .DIN3(n1108), .Q(n1106) );
  nnd2s3 U205 ( .DIN1(n2500), .DIN2(n1052), .Q(n1108) );
  nnd2s3 U206 ( .DIN1(n538), .DIN2(n1109), .Q(n1107) );
  xor2s3 U207 ( .DIN1(n2039), .DIN2(n659), .Q(n1109) );
  nnd2s3 U208 ( .DIN1(n1045), .DIN2(n1110), .Q(g9339) );
  nnd2s3 U209 ( .DIN1(n1111), .DIN2(n540), .Q(n1110) );
  xor2s3 U210 ( .DIN1(n1113), .DIN2(n2039), .Q(n1111) );
  nnd2s3 U211 ( .DIN1(n1050), .DIN2(n1114), .Q(n1113) );
  nnd2s3 U212 ( .DIN1(n2501), .DIN2(n1052), .Q(n1114) );
  nnd2s3 U213 ( .DIN1(n538), .DIN2(n1115), .Q(n1050) );
  nnd2s3 U214 ( .DIN1(n1116), .DIN2(n1117), .Q(n1052) );
  nnd2s3 U215 ( .DIN1(n542), .DIN2(n728), .Q(n1117) );
  nnd4s2 U216 ( .DIN1(n1118), .DIN2(n948), .DIN3(n964), .DIN4(n1112), .Q(n1045) );
  nnd2s3 U217 ( .DIN1(n911), .DIN2(n1119), .Q(g9338) );
  nnd2s3 U218 ( .DIN1(n1120), .DIN2(n850), .Q(n1119) );
  nnd2s3 U219 ( .DIN1(n1112), .DIN2(n1121), .Q(n1120) );
  nnd2s3 U220 ( .DIN1(n948), .DIN2(n964), .Q(n1121) );
  nnd2s3 U221 ( .DIN1(n948), .DIN2(n915), .Q(n1112) );
  nnd3s3 U222 ( .DIN1(n539), .DIN2(n662), .DIN3(n1987), .Q(n911) );
  nnd3s3 U223 ( .DIN1(n1122), .DIN2(n1123), .DIN3(n541), .Q(n915) );
  nnd2s3 U224 ( .DIN1(n542), .DIN2(n1124), .Q(n1115) );
  nnd2s3 U225 ( .DIN1(n1125), .DIN2(n964), .Q(n1124) );
  nnd3s3 U226 ( .DIN1(n663), .DIN2(n797), .DIN3(n1982), .Q(n964) );
  or2s3 U227 ( .DIN1(n1981), .DIN2(n1126), .Q(n1125) );
  nnd2s3 U228 ( .DIN1(n1053), .DIN2(n661), .Q(n1123) );
  or5s3 U229 ( .DIN1(n2029), .DIN2(n1994), .DIN3(n1958), .DIN4(n1955), .DIN5(
        n592), .Q(n1053) );
  nor2s3 U230 ( .DIN1(n1087), .DIN2(n1933), .Q(n1062) );
  or4s3 U231 ( .DIN1(n659), .DIN2(n1936), .DIN3(n1968), .DIN4(n2039), .Q(n1087) );
  nnd2s3 U232 ( .DIN1(n2009), .DIN2(n1054), .Q(n1122) );
  or5s3 U233 ( .DIN1(n593), .DIN2(n867), .DIN3(n866), .DIN4(n710), .DIN5(n838), 
        .Q(n1054) );
  nor2s3 U234 ( .DIN1(n687), .DIN2(n1088), .Q(n1063) );
  nnd4s2 U235 ( .DIN1(n2039), .DIN2(n1968), .DIN3(n1936), .DIN4(n659), .Q(
        n1088) );
  nnd2s3 U236 ( .DIN1(n952), .DIN2(n691), .Q(n1103) );
  and2s3 U237 ( .DIN1(n957), .DIN2(n1127), .Q(n952) );
  or2s3 U238 ( .DIN1(n965), .DIN2(n660), .Q(n1127) );
  nor2s3 U239 ( .DIN1(n1128), .DIN2(n2865), .Q(g8993) );
  xor2s3 U240 ( .DIN1(n1129), .DIN2(n2527), .Q(n1128) );
  nor2s3 U241 ( .DIN1(n1130), .DIN2(n2865), .Q(g8992) );
  xor2s3 U242 ( .DIN1(n1131), .DIN2(n2526), .Q(n1130) );
  nor2s3 U243 ( .DIN1(n1132), .DIN2(n2865), .Q(g8991) );
  xor2s3 U244 ( .DIN1(n1133), .DIN2(n2525), .Q(n1132) );
  nor2s3 U245 ( .DIN1(n1134), .DIN2(n2865), .Q(g8990) );
  xor2s3 U246 ( .DIN1(n2524), .DIN2(n1135), .Q(n1134) );
  nor2s3 U247 ( .DIN1(n1136), .DIN2(n2865), .Q(g8989) );
  xor2s3 U248 ( .DIN1(n1137), .DIN2(n2523), .Q(n1136) );
  nor2s3 U249 ( .DIN1(n1138), .DIN2(n2865), .Q(g8988) );
  xor2s3 U250 ( .DIN1(n1139), .DIN2(n2522), .Q(n1138) );
  nor2s3 U251 ( .DIN1(n1140), .DIN2(n2865), .Q(g8987) );
  xor2s3 U252 ( .DIN1(n1141), .DIN2(n2588), .Q(n1140) );
  nnd2s3 U253 ( .DIN1(n1142), .DIN2(n1143), .Q(g8874) );
  nnd2s3 U254 ( .DIN1(n2848), .DIN2(n1141), .Q(n1143) );
  nnd2s3 U255 ( .DIN1(n1144), .DIN2(n1145), .Q(n1141) );
  nnd2s3 U256 ( .DIN1(n1146), .DIN2(n2863), .Q(n1145) );
  xor2s3 U257 ( .DIN1(n1147), .DIN2(n1970), .Q(n1146) );
  nnd3s3 U258 ( .DIN1(n1148), .DIN2(n717), .DIN3(n1976), .Q(n1147) );
  nnd2s3 U259 ( .DIN1(n2854), .DIN2(n628), .Q(n1142) );
  nnd2s3 U260 ( .DIN1(n1150), .DIN2(n1151), .Q(g8873) );
  nnd2s3 U261 ( .DIN1(n2848), .DIN2(n1139), .Q(n1151) );
  nnd2s3 U262 ( .DIN1(n1152), .DIN2(n1153), .Q(n1139) );
  nnd2s3 U263 ( .DIN1(n1154), .DIN2(n2863), .Q(n1153) );
  xor2s3 U264 ( .DIN1(n1155), .DIN2(n1944), .Q(n1154) );
  nnd2s3 U265 ( .DIN1(n1156), .DIN2(n1976), .Q(n1155) );
  nnd2s3 U266 ( .DIN1(n2852), .DIN2(n764), .Q(n1150) );
  nnd2s3 U267 ( .DIN1(n1157), .DIN2(n1158), .Q(g8872) );
  nnd2s3 U268 ( .DIN1(n2848), .DIN2(n1137), .Q(n1158) );
  nnd3s3 U269 ( .DIN1(n1159), .DIN2(n1160), .DIN3(n1161), .Q(n1137) );
  nnd3s3 U270 ( .DIN1(n2861), .DIN2(n665), .DIN3(n1162), .Q(n1161) );
  nnd3s3 U271 ( .DIN1(n620), .DIN2(n787), .DIN3(n1163), .Q(n1162) );
  nnd4s2 U272 ( .DIN1(n2013), .DIN2(n1164), .DIN3(n620), .DIN4(n787), .Q(n1159) );
  nnd2s3 U273 ( .DIN1(n2852), .DIN2(n558), .Q(n1157) );
  nnd2s3 U274 ( .DIN1(n1165), .DIN2(n1166), .Q(g8871) );
  nnd2s3 U275 ( .DIN1(n2849), .DIN2(n1135), .Q(n1166) );
  nnd3s3 U276 ( .DIN1(n1167), .DIN2(n1168), .DIN3(n1169), .Q(n1135) );
  nnd4s2 U277 ( .DIN1(n1971), .DIN2(n1974), .DIN3(n1164), .DIN4(n620), .Q(
        n1168) );
  nnd3s3 U278 ( .DIN1(n2861), .DIN2(n794), .DIN3(n1170), .Q(n1167) );
  nnd3s3 U279 ( .DIN1(n1163), .DIN2(n620), .DIN3(n1974), .Q(n1170) );
  nnd2s3 U280 ( .DIN1(n2852), .DIN2(n735), .Q(n1165) );
  nnd2s3 U281 ( .DIN1(n1171), .DIN2(n1172), .Q(g8870) );
  nnd2s3 U282 ( .DIN1(n2848), .DIN2(n1133), .Q(n1172) );
  nnd2s3 U283 ( .DIN1(n1173), .DIN2(n1174), .Q(n1133) );
  nnd2s3 U284 ( .DIN1(n1175), .DIN2(n2863), .Q(n1174) );
  xnr2s3 U285 ( .DIN1(n1945), .DIN2(n1176), .Q(n1175) );
  nor2s3 U286 ( .DIN1(n1974), .DIN2(n1177), .Q(n1176) );
  nnd2s3 U287 ( .DIN1(n2852), .DIN2(n643), .Q(n1171) );
  nnd2s3 U288 ( .DIN1(n1178), .DIN2(n1179), .Q(g8869) );
  nnd2s3 U289 ( .DIN1(n2848), .DIN2(n1131), .Q(n1179) );
  nnd2s3 U290 ( .DIN1(n1180), .DIN2(n1181), .Q(n1131) );
  nnd2s3 U291 ( .DIN1(n1182), .DIN2(n2862), .Q(n1181) );
  xor2s3 U292 ( .DIN1(n1183), .DIN2(n2014), .Q(n1182) );
  or2s3 U293 ( .DIN1(n787), .DIN2(n1177), .Q(n1183) );
  nnd3s3 U294 ( .DIN1(n1949), .DIN2(n620), .DIN3(n1976), .Q(n1177) );
  or2s3 U295 ( .DIN1(n2850), .DIN2(n2705), .Q(n1178) );
  nnd2s3 U296 ( .DIN1(n1184), .DIN2(n1185), .Q(g8868) );
  nnd2s3 U297 ( .DIN1(n2849), .DIN2(n1129), .Q(n1185) );
  nnd3s3 U298 ( .DIN1(n1186), .DIN2(n1187), .DIN3(n1188), .Q(n1129) );
  nnd3s3 U299 ( .DIN1(n2861), .DIN2(n585), .DIN3(n1189), .Q(n1188) );
  nnd2s3 U300 ( .DIN1(n1148), .DIN2(n1163), .Q(n1189) );
  nnd3s3 U301 ( .DIN1(n1164), .DIN2(n1148), .DIN3(n2015), .Q(n1186) );
  and2s3 U302 ( .DIN1(n1163), .DIN2(n2863), .Q(n1164) );
  or2s3 U303 ( .DIN1(n2849), .DIN2(n2707), .Q(n1184) );
  nnd3s3 U304 ( .DIN1(n1190), .DIN2(n948), .DIN3(n1191), .Q(g8782) );
  nnd2s3 U305 ( .DIN1(n1192), .DIN2(n774), .Q(n1191) );
  nnd2s3 U306 ( .DIN1(n1193), .DIN2(n1194), .Q(g8781) );
  nnd2s3 U307 ( .DIN1(n1195), .DIN2(n948), .Q(n1194) );
  nnd2s3 U308 ( .DIN1(n1196), .DIN2(n1197), .Q(n1195) );
  nnd2s3 U309 ( .DIN1(n1198), .DIN2(g2613), .Q(n1197) );
  nnd3s3 U310 ( .DIN1(g5656), .DIN2(n1199), .DIN3(n1200), .Q(n1198) );
  xor2s3 U311 ( .DIN1(n1201), .DIN2(n1202), .Q(n1200) );
  nor2s3 U312 ( .DIN1(n1203), .DIN2(n1204), .Q(n1202) );
  nor2s3 U313 ( .DIN1(n1981), .DIN2(n965), .Q(n1204) );
  nor2s3 U314 ( .DIN1(n1205), .DIN2(n830), .Q(n1203) );
  nor2s3 U315 ( .DIN1(n658), .DIN2(n797), .Q(n1205) );
  nnd2s3 U316 ( .DIN1(g5644), .DIN2(n850), .Q(n1201) );
  nnd3s3 U317 ( .DIN1(n1206), .DIN2(n965), .DIN3(n1975), .Q(n1199) );
  nnd2s3 U318 ( .DIN1(n663), .DIN2(n1207), .Q(n1206) );
  nnd2s3 U319 ( .DIN1(n1126), .DIN2(n728), .Q(n1207) );
  or2s3 U320 ( .DIN1(n957), .DIN2(n850), .Q(n1196) );
  nnd2s3 U321 ( .DIN1(n657), .DIN2(n1208), .Q(n1193) );
  nnd3s3 U322 ( .DIN1(n1209), .DIN2(n669), .DIN3(n1210), .Q(n1208) );
  nnd2s3 U323 ( .DIN1(n1211), .DIN2(n1212), .Q(n1210) );
  or2s3 U324 ( .DIN1(n2556), .DIN2(n1999), .Q(n1211) );
  nnd2s3 U325 ( .DIN1(n1213), .DIN2(n1214), .Q(n1209) );
  or2s3 U326 ( .DIN1(n2512), .DIN2(n2050), .Q(n1214) );
  or2s3 U327 ( .DIN1(n2049), .DIN2(n2043), .Q(n1213) );
  nor2s3 U328 ( .DIN1(n1215), .DIN2(n2861), .Q(g8780) );
  xor2s3 U329 ( .DIN1(n1216), .DIN2(n1982), .Q(n1215) );
  nnd2s3 U330 ( .DIN1(n1190), .DIN2(n1217), .Q(n1216) );
  or2s3 U331 ( .DIN1(n1116), .DIN2(n728), .Q(n1217) );
  nnd4s2 U332 ( .DIN1(n1126), .DIN2(n1975), .DIN3(n542), .DIN4(n663), .Q(n1116) );
  nnd2s3 U333 ( .DIN1(n537), .DIN2(n820), .Q(n1190) );
  nnd3s3 U334 ( .DIN1(n1218), .DIN2(n927), .DIN3(n1219), .Q(g8695) );
  nnd2s3 U335 ( .DIN1(n1220), .DIN2(n514), .Q(n1219) );
  nor2s3 U336 ( .DIN1(n1221), .DIN2(n2861), .Q(g8694) );
  xor2s3 U337 ( .DIN1(n1222), .DIN2(n1983), .Q(n1221) );
  nnd2s3 U338 ( .DIN1(n1218), .DIN2(n1223), .Q(n1222) );
  or2s3 U339 ( .DIN1(n1038), .DIN2(n747), .Q(n1223) );
  nnd4s2 U340 ( .DIN1(n1043), .DIN2(n1948), .DIN3(n920), .DIN4(n702), .Q(n1038) );
  nnd2s3 U341 ( .DIN1(n587), .DIN2(n788), .Q(n1218) );
  nor2s3 U342 ( .DIN1(n778), .DIN2(n1224), .Q(g8573) );
  xor2s3 U343 ( .DIN1(n670), .DIN2(n1225), .Q(n1224) );
  nor2s3 U344 ( .DIN1(n2045), .DIN2(n1226), .Q(g8572) );
  nor2s3 U345 ( .DIN1(n2046), .DIN2(n1226), .Q(g8571) );
  nor2s3 U346 ( .DIN1(n2007), .DIN2(n1226), .Q(g8570) );
  nor2s3 U347 ( .DIN1(n2047), .DIN2(n1226), .Q(g8569) );
  nnd2s3 U348 ( .DIN1(g109), .DIN2(n1227), .Q(n1226) );
  nnd3s3 U349 ( .DIN1(n905), .DIN2(\DFF_436/net723 ), .DIN3(n1228), .Q(n1227)
         );
  nor2s3 U350 ( .DIN1(n1229), .DIN2(n1230), .Q(g8568) );
  xor2s3 U351 ( .DIN1(n669), .DIN2(n1231), .Q(n1230) );
  and3s3 U352 ( .DIN1(n1232), .DIN2(n907), .DIN3(n841), .Q(g8567) );
  or3s3 U353 ( .DIN1(n2055), .DIN2(n2511), .DIN3(n1233), .Q(n907) );
  nnd2s3 U354 ( .DIN1(n2055), .DIN2(n1234), .Q(n1232) );
  or2s3 U355 ( .DIN1(n1233), .DIN2(n2511), .Q(n1234) );
  nnd2s3 U356 ( .DIN1(n1235), .DIN2(n1236), .Q(g8566) );
  nnd2s3 U357 ( .DIN1(n718), .DIN2(n579), .Q(n1236) );
  nnd2s3 U359 ( .DIN1(n1237), .DIN2(n1238), .Q(g8565) );
  nnd2s3 U360 ( .DIN1(n718), .DIN2(n829), .Q(n1238) );
  nnd2s3 U362 ( .DIN1(n1239), .DIN2(n1240), .Q(g8564) );
  nnd2s3 U363 ( .DIN1(n718), .DIN2(n758), .Q(n1240) );
  nnd2s3 U365 ( .DIN1(n1241), .DIN2(n1242), .Q(g8563) );
  nnd2s3 U366 ( .DIN1(n718), .DIN2(n815), .Q(n1242) );
  nnd2s3 U368 ( .DIN1(n1243), .DIN2(n1244), .Q(g8562) );
  nnd2s3 U369 ( .DIN1(n718), .DIN2(n832), .Q(n1244) );
  nnd2s3 U371 ( .DIN1(n1245), .DIN2(n1246), .Q(g8561) );
  nnd2s3 U372 ( .DIN1(n718), .DIN2(n858), .Q(n1246) );
  and3s3 U374 ( .DIN1(n1225), .DIN2(n2061), .DIN3(n1247), .Q(g8450) );
  nnd2s3 U375 ( .DIN1(n2623), .DIN2(n531), .Q(n1247) );
  nnd2s3 U376 ( .DIN1(n1248), .DIN2(n812), .Q(n1225) );
  nnd2s3 U377 ( .DIN1(n1249), .DIN2(n1250), .Q(g8449) );
  nnd2s3 U378 ( .DIN1(n2849), .DIN2(n1251), .Q(n1250) );
  xnr2s3 U379 ( .DIN1(n2585), .DIN2(n1252), .Q(n1251) );
  nnd2s3 U380 ( .DIN1(n1156), .DIN2(n855), .Q(n1252) );
  and2s3 U381 ( .DIN1(n1253), .DIN2(n717), .Q(n1156) );
  nnd2s3 U382 ( .DIN1(n2853), .DIN2(n604), .Q(n1249) );
  nnd2s3 U383 ( .DIN1(n1254), .DIN2(n1255), .Q(g8448) );
  nnd2s3 U384 ( .DIN1(n1256), .DIN2(n2849), .Q(n1255) );
  xor2s3 U385 ( .DIN1(n1257), .DIN2(n1969), .Q(n1256) );
  nnd2s3 U386 ( .DIN1(n1253), .DIN2(n1163), .Q(n1257) );
  nor2s3 U387 ( .DIN1(n717), .DIN2(n1976), .Q(n1163) );
  nor2s3 U388 ( .DIN1(n787), .DIN2(n620), .Q(n1253) );
  or2s3 U389 ( .DIN1(n2849), .DIN2(n2709), .Q(n1254) );
  nor2s3 U390 ( .DIN1(n1258), .DIN2(n2865), .Q(g8447) );
  xor2s3 U391 ( .DIN1(n1259), .DIN2(n2542), .Q(n1258) );
  nor2s3 U392 ( .DIN1(n2870), .DIN2(n1260), .Q(g8446) );
  xor2s3 U393 ( .DIN1(n603), .DIN2(n1261), .Q(n1260) );
  nor2s3 U394 ( .DIN1(n2870), .DIN2(n1262), .Q(g8445) );
  xnr2s3 U395 ( .DIN1(n2534), .DIN2(n1263), .Q(n1262) );
  nor2s3 U396 ( .DIN1(n2870), .DIN2(n1264), .Q(g8444) );
  xnr2s3 U397 ( .DIN1(n2533), .DIN2(n1265), .Q(n1264) );
  nor2s3 U398 ( .DIN1(n1266), .DIN2(n2868), .Q(g8443) );
  xor2s3 U399 ( .DIN1(n1267), .DIN2(n2532), .Q(n1266) );
  nor2s3 U400 ( .DIN1(n1268), .DIN2(n2868), .Q(g8442) );
  xor2s3 U401 ( .DIN1(n1269), .DIN2(n2531), .Q(n1268) );
  nor2s3 U402 ( .DIN1(n1270), .DIN2(n2868), .Q(g8441) );
  xor2s3 U403 ( .DIN1(n1271), .DIN2(n2530), .Q(n1270) );
  nor2s3 U404 ( .DIN1(n1272), .DIN2(n2868), .Q(g8440) );
  xor2s3 U405 ( .DIN1(n1273), .DIN2(n2529), .Q(n1272) );
  nor2s3 U406 ( .DIN1(n1274), .DIN2(n2869), .Q(g8439) );
  xor2s3 U407 ( .DIN1(n1275), .DIN2(n2528), .Q(n1274) );
  nor2s3 U408 ( .DIN1(n1276), .DIN2(n2867), .Q(g8438) );
  xor2s3 U409 ( .DIN1(n1277), .DIN2(n1991), .Q(n1276) );
  and3s3 U410 ( .DIN1(n1278), .DIN2(n1231), .DIN3(n695), .Q(g8437) );
  or2s3 U411 ( .DIN1(n1279), .DIN2(n2043), .Q(n1231) );
  nnd2s3 U412 ( .DIN1(n2043), .DIN2(n1279), .Q(n1278) );
  nor2s3 U413 ( .DIN1(n1280), .DIN2(n1281), .Q(g8436) );
  xnr2s3 U414 ( .DIN1(n2511), .DIN2(n1233), .Q(n1281) );
  nnd2s3 U415 ( .DIN1(n1282), .DIN2(n1283), .Q(g8435) );
  nnd2s3 U416 ( .DIN1(n1284), .DIN2(n820), .Q(n1283) );
  nnd2s3 U417 ( .DIN1(n537), .DIN2(n610), .Q(n1282) );
  nnd2s3 U418 ( .DIN1(n1285), .DIN2(n1286), .Q(g8434) );
  nnd2s3 U419 ( .DIN1(n1284), .DIN2(n610), .Q(n1286) );
  nnd2s3 U420 ( .DIN1(n537), .DIN2(n845), .Q(n1285) );
  nnd2s3 U421 ( .DIN1(n1287), .DIN2(n1288), .Q(g8433) );
  nnd2s3 U422 ( .DIN1(n1284), .DIN2(n845), .Q(n1288) );
  nnd2s3 U423 ( .DIN1(n537), .DIN2(n864), .Q(n1287) );
  nnd2s3 U424 ( .DIN1(n1289), .DIN2(n1290), .Q(g8432) );
  nnd2s3 U425 ( .DIN1(n1284), .DIN2(n864), .Q(n1290) );
  nnd2s3 U426 ( .DIN1(n537), .DIN2(n715), .Q(n1289) );
  nnd2s3 U427 ( .DIN1(n1291), .DIN2(n1292), .Q(g8431) );
  nnd2s3 U428 ( .DIN1(n1284), .DIN2(n715), .Q(n1292) );
  nnd2s3 U429 ( .DIN1(n537), .DIN2(n534), .Q(n1291) );
  nnd2s3 U430 ( .DIN1(n1293), .DIN2(n1294), .Q(g8430) );
  nnd2s3 U431 ( .DIN1(n1284), .DIN2(n534), .Q(n1294) );
  nnd2s3 U432 ( .DIN1(n537), .DIN2(n835), .Q(n1293) );
  nnd2s3 U433 ( .DIN1(n1295), .DIN2(n1296), .Q(g8429) );
  nnd2s3 U434 ( .DIN1(n1284), .DIN2(n835), .Q(n1296) );
  nnd2s3 U435 ( .DIN1(n537), .DIN2(n563), .Q(n1295) );
  nnd2s3 U436 ( .DIN1(n1297), .DIN2(n1298), .Q(g8428) );
  nnd2s3 U437 ( .DIN1(n1284), .DIN2(n563), .Q(n1298) );
  nor2s3 U438 ( .DIN1(n537), .DIN2(n657), .Q(n1284) );
  nnd2s3 U439 ( .DIN1(n537), .DIN2(n774), .Q(n1297) );
  nnd3s3 U440 ( .DIN1(n542), .DIN2(n728), .DIN3(n1975), .Q(n1192) );
  nor2s3 U441 ( .DIN1(n1299), .DIN2(n2868), .Q(g8427) );
  xor2s3 U442 ( .DIN1(g7750), .DIN2(n1937), .Q(n1299) );
  nor2s3 U443 ( .DIN1(n1300), .DIN2(n2869), .Q(g8426) );
  xor2s3 U444 ( .DIN1(g7752), .DIN2(n1992), .Q(n1300) );
  nor2s3 U445 ( .DIN1(n1301), .DIN2(n2869), .Q(g8425) );
  xor2s3 U446 ( .DIN1(g7753), .DIN2(n1959), .Q(n1301) );
  nor2s3 U447 ( .DIN1(n1302), .DIN2(n2869), .Q(g8424) );
  xor2s3 U448 ( .DIN1(g7754), .DIN2(n2520), .Q(n1302) );
  nor2s3 U449 ( .DIN1(n1303), .DIN2(n2869), .Q(g8423) );
  xor2s3 U450 ( .DIN1(g7755), .DIN2(n2519), .Q(n1303) );
  nor2s3 U451 ( .DIN1(n1304), .DIN2(n2869), .Q(g8422) );
  xor2s3 U452 ( .DIN1(g7756), .DIN2(n1960), .Q(n1304) );
  nor2s3 U453 ( .DIN1(n1305), .DIN2(n2869), .Q(g8421) );
  xor2s3 U454 ( .DIN1(g7757), .DIN2(n1996), .Q(n1305) );
  nor2s3 U455 ( .DIN1(n1306), .DIN2(n2869), .Q(g8420) );
  xor2s3 U456 ( .DIN1(g7758), .DIN2(n1961), .Q(n1306) );
  nor2s3 U457 ( .DIN1(n1307), .DIN2(n2869), .Q(g8419) );
  xor2s3 U458 ( .DIN1(g7759), .DIN2(n1938), .Q(n1307) );
  nor2s3 U459 ( .DIN1(n1308), .DIN2(n2869), .Q(g8418) );
  xor2s3 U460 ( .DIN1(g7751), .DIN2(n2518), .Q(n1308) );
  nnd2s3 U461 ( .DIN1(n2022), .DIN2(n904), .Q(g8352) );
  nnd2s3 U462 ( .DIN1(n2023), .DIN2(n904), .Q(g8349) );
  nnd2s3 U463 ( .DIN1(n2038), .DIN2(n904), .Q(g8347) );
  nnd2s3 U464 ( .DIN1(n2034), .DIN2(n904), .Q(g8340) );
  nnd2s3 U465 ( .DIN1(n2018), .DIN2(n904), .Q(g8335) );
  nnd2s3 U466 ( .DIN1(n2035), .DIN2(n904), .Q(g8331) );
  nnd2s3 U467 ( .DIN1(n2019), .DIN2(n904), .Q(g8328) );
  nnd2s3 U468 ( .DIN1(n2036), .DIN2(n904), .Q(g8323) );
  nnd2s3 U469 ( .DIN1(n2020), .DIN2(n904), .Q(g8318) );
  nnd2s3 U470 ( .DIN1(n2037), .DIN2(n904), .Q(g8316) );
  nnd2s3 U471 ( .DIN1(n2021), .DIN2(n904), .Q(g8313) );
  nnd2s3 U472 ( .DIN1(n1309), .DIN2(n1310), .Q(g8288) );
  nnd2s3 U473 ( .DIN1(n1311), .DIN2(n788), .Q(n1310) );
  nnd2s3 U474 ( .DIN1(n587), .DIN2(n689), .Q(n1309) );
  nnd2s3 U475 ( .DIN1(n1312), .DIN2(n1313), .Q(g8287) );
  nnd2s3 U476 ( .DIN1(n1311), .DIN2(n689), .Q(n1313) );
  nnd2s3 U477 ( .DIN1(n587), .DIN2(n644), .Q(n1312) );
  nnd2s3 U478 ( .DIN1(n1314), .DIN2(n1315), .Q(g8286) );
  nnd2s3 U479 ( .DIN1(n1311), .DIN2(n644), .Q(n1315) );
  nnd2s3 U480 ( .DIN1(n587), .DIN2(n672), .Q(n1314) );
  nnd2s3 U481 ( .DIN1(n1316), .DIN2(n1317), .Q(g8285) );
  nnd2s3 U482 ( .DIN1(n1311), .DIN2(n672), .Q(n1317) );
  nnd2s3 U483 ( .DIN1(n587), .DIN2(n755), .Q(n1316) );
  nnd2s3 U484 ( .DIN1(n1318), .DIN2(n1319), .Q(g8284) );
  nnd2s3 U485 ( .DIN1(n1311), .DIN2(n755), .Q(n1319) );
  nnd2s3 U486 ( .DIN1(n587), .DIN2(n560), .Q(n1318) );
  nnd2s3 U487 ( .DIN1(n1320), .DIN2(n1321), .Q(g8283) );
  nnd2s3 U488 ( .DIN1(n1311), .DIN2(n560), .Q(n1321) );
  nnd2s3 U489 ( .DIN1(n587), .DIN2(n821), .Q(n1320) );
  nnd2s3 U490 ( .DIN1(n1322), .DIN2(n1323), .Q(g8282) );
  nnd2s3 U491 ( .DIN1(n1311), .DIN2(n821), .Q(n1323) );
  nnd2s3 U492 ( .DIN1(n587), .DIN2(n668), .Q(n1322) );
  nnd2s3 U493 ( .DIN1(n1324), .DIN2(n1325), .Q(g8281) );
  nnd2s3 U494 ( .DIN1(n1311), .DIN2(n668), .Q(n1325) );
  nor2s3 U495 ( .DIN1(n587), .DIN2(n591), .Q(n1311) );
  nnd2s3 U496 ( .DIN1(n587), .DIN2(n514), .Q(n1324) );
  nnd3s3 U497 ( .DIN1(n920), .DIN2(n747), .DIN3(n1948), .Q(n1220) );
  and3s3 U498 ( .DIN1(n531), .DIN2(n2061), .DIN3(n1326), .Q(g8280) );
  nnd2s3 U499 ( .DIN1(n1952), .DIN2(n1327), .Q(n1326) );
  nor2s3 U500 ( .DIN1(n1327), .DIN2(n1952), .Q(n1248) );
  nor2s3 U501 ( .DIN1(n1328), .DIN2(n1329), .Q(g8279) );
  nor2s3 U502 ( .DIN1(n1330), .DIN2(n856), .Q(n1328) );
  nor2s3 U503 ( .DIN1(n1331), .DIN2(n1329), .Q(g8278) );
  nor2s3 U504 ( .DIN1(n1332), .DIN2(n1333), .Q(n1331) );
  nor2s3 U505 ( .DIN1(n2601), .DIN2(n1330), .Q(n1333) );
  nor2s3 U506 ( .DIN1(n1334), .DIN2(n2601), .Q(n1330) );
  nor2s3 U507 ( .DIN1(n1335), .DIN2(n1334), .Q(n1332) );
  and3s3 U508 ( .DIN1(n1336), .DIN2(n1334), .DIN3(n700), .Q(g8277) );
  or2s3 U509 ( .DIN1(n1337), .DIN2(n2603), .Q(n1334) );
  nnd2s3 U510 ( .DIN1(n2603), .DIN2(n1337), .Q(n1336) );
  or2s3 U511 ( .DIN1(n1338), .DIN2(n2602), .Q(n1337) );
  nor2s3 U512 ( .DIN1(n1329), .DIN2(n1339), .Q(g8276) );
  xnr2s3 U513 ( .DIN1(n2602), .DIN2(n1338), .Q(n1339) );
  nnd2s3 U514 ( .DIN1(n649), .DIN2(n1340), .Q(n1338) );
  nnd2s3 U515 ( .DIN1(n2578), .DIN2(g109), .Q(n1329) );
  and3s3 U516 ( .DIN1(n1341), .DIN2(n1279), .DIN3(n695), .Q(g8274) );
  or3s3 U517 ( .DIN1(n2049), .DIN2(n2512), .DIN3(n1342), .Q(n1279) );
  nnd2s3 U518 ( .DIN1(n2049), .DIN2(n1343), .Q(n1341) );
  or2s3 U519 ( .DIN1(n1342), .DIN2(n2512), .Q(n1343) );
  and3s3 U520 ( .DIN1(n1344), .DIN2(n1233), .DIN3(n841), .Q(g8273) );
  or3s3 U521 ( .DIN1(n2056), .DIN2(n2513), .DIN3(n1345), .Q(n1233) );
  nnd2s3 U522 ( .DIN1(n2056), .DIN2(n1346), .Q(n1344) );
  or2s3 U523 ( .DIN1(n1345), .DIN2(n2513), .Q(n1346) );
  nnd2s3 U524 ( .DIN1(n1347), .DIN2(n1348), .Q(g8272) );
  or4s3 U525 ( .DIN1(n1349), .DIN2(n1350), .DIN3(n1351), .DIN4(n1352), .Q(
        n1348) );
  nnd4s2 U526 ( .DIN1(n1960), .DIN2(n1959), .DIN3(n1992), .DIN4(n1937), .Q(
        n1352) );
  nnd4s2 U527 ( .DIN1(n656), .DIN2(n814), .DIN3(n688), .DIN4(n749), .Q(n1351)
         );
  nnd4s2 U528 ( .DIN1(n2017), .DIN2(n1926), .DIN3(n1925), .DIN4(g7749), .Q(
        n1350) );
  nnd4s2 U529 ( .DIN1(n1353), .DIN2(n1938), .DIN3(n1961), .DIN4(n1996), .Q(
        n1349) );
  nnd2s3 U530 ( .DIN1(g109), .DIN2(n869), .Q(n1347) );
  and2s3 U531 ( .DIN1(n1354), .DIN2(n2061), .Q(g8080) );
  nnd2s3 U532 ( .DIN1(n1355), .DIN2(n1356), .Q(n1354) );
  nnd3s3 U533 ( .DIN1(n1357), .DIN2(n836), .DIN3(n2025), .Q(n1356) );
  nnd2s3 U534 ( .DIN1(n1327), .DIN2(n828), .Q(n1355) );
  nnd3s3 U535 ( .DIN1(n828), .DIN2(n836), .DIN3(n1357), .Q(n1327) );
  or2s3 U536 ( .DIN1(n1358), .DIN2(n1359), .Q(g8079) );
  nor2s3 U537 ( .DIN1(n2775), .DIN2(n2869), .Q(n1359) );
  nor6s3 U538 ( .DIN1(n1360), .DIN2(n1361), .DIN3(n1362), .DIN4(n852), .DIN5(
        n1363), .DIN6(n817), .Q(n1358) );
  nnd4s2 U539 ( .DIN1(n1991), .DIN2(n2529), .DIN3(n2533), .DIN4(n2534), .Q(
        n1362) );
  nnd4s2 U540 ( .DIN1(n741), .DIN2(n763), .DIN3(n536), .DIN4(n603), .Q(n1361)
         );
  nnd4s2 U541 ( .DIN1(n719), .DIN2(n780), .DIN3(n816), .DIN4(n694), .Q(n1360)
         );
  or2s3 U542 ( .DIN1(n1364), .DIN2(n1365), .Q(g8078) );
  nor2s3 U543 ( .DIN1(n2764), .DIN2(n2869), .Q(n1365) );
  nor6s3 U544 ( .DIN1(n1366), .DIN2(n1367), .DIN3(n1368), .DIN4(n783), .DIN5(
        n805), .DIN6(n810), .Q(n1364) );
  nnd4s2 U545 ( .DIN1(g7335), .DIN2(n516), .DIN3(n2526), .DIN4(n559), .Q(n1368) );
  nnd4s2 U546 ( .DIN1(n795), .DIN2(n819), .DIN3(n859), .DIN4(n801), .Q(n1367)
         );
  nnd4s2 U547 ( .DIN1(n742), .DIN2(n846), .DIN3(n555), .DIN4(n851), .Q(n1366)
         );
  nor2s3 U548 ( .DIN1(n1229), .DIN2(n1369), .Q(g8077) );
  xnr2s3 U549 ( .DIN1(n2512), .DIN2(n1342), .Q(n1369) );
  nor2s3 U550 ( .DIN1(n1280), .DIN2(n1370), .Q(g8076) );
  xnr2s3 U551 ( .DIN1(n2513), .DIN2(n1345), .Q(n1370) );
  nnd3s3 U552 ( .DIN1(n948), .DIN2(n1371), .DIN3(n1372), .Q(g8067) );
  nnd2s3 U553 ( .DIN1(n1373), .DIN2(n766), .Q(n1372) );
  nnd2s3 U554 ( .DIN1(n543), .DIN2(n629), .Q(n1373) );
  and3s3 U555 ( .DIN1(n948), .DIN2(n1371), .DIN3(n1374), .Q(g8066) );
  xor2s3 U556 ( .DIN1(n2515), .DIN2(n543), .Q(n1374) );
  and3s3 U557 ( .DIN1(n948), .DIN2(n1371), .DIN3(n1375), .Q(g8065) );
  nnd2s3 U558 ( .DIN1(n1376), .DIN2(n1377), .Q(n1375) );
  nnd2s3 U559 ( .DIN1(n1378), .DIN2(n833), .Q(n1377) );
  nnd2s3 U560 ( .DIN1(n2517), .DIN2(n2558), .Q(n1378) );
  nnd2s3 U561 ( .DIN1(n1379), .DIN2(n948), .Q(g8064) );
  xor2s3 U562 ( .DIN1(n2517), .DIN2(n2558), .Q(n1379) );
  nnd3s3 U563 ( .DIN1(n1380), .DIN2(n948), .DIN3(n1381), .Q(g8063) );
  nnd2s3 U564 ( .DIN1(n1371), .DIN2(n830), .Q(n1381) );
  nnd3s3 U565 ( .DIN1(n542), .DIN2(n1382), .DIN3(n1981), .Q(n1380) );
  nnd3s3 U566 ( .DIN1(n960), .DIN2(n965), .DIN3(n1118), .Q(n1382) );
  and2s3 U567 ( .DIN1(n957), .DIN2(n1383), .Q(n1118) );
  nnd2s3 U568 ( .DIN1(n1978), .DIN2(n691), .Q(n1383) );
  nnd3s3 U569 ( .DIN1(n1985), .DIN2(n660), .DIN3(n1951), .Q(n957) );
  nnd2s3 U570 ( .DIN1(n1951), .DIN2(n691), .Q(n965) );
  nnd2s3 U571 ( .DIN1(n660), .DIN2(n663), .Q(n960) );
  nnd3s3 U572 ( .DIN1(n543), .DIN2(n629), .DIN3(n2514), .Q(n1371) );
  nnd3s3 U573 ( .DIN1(n2517), .DIN2(n2558), .DIN3(n2516), .Q(n1376) );
  nnd2s3 U574 ( .DIN1(n1384), .DIN2(n1385), .Q(g7817) );
  nnd2s3 U575 ( .DIN1(n1386), .DIN2(n809), .Q(n1385) );
  nor2s3 U576 ( .DIN1(n1387), .DIN2(n590), .Q(g7816) );
  nor2s3 U577 ( .DIN1(n1388), .DIN2(n666), .Q(n1387) );
  nor2s3 U578 ( .DIN1(n1389), .DIN2(n862), .Q(n1388) );
  nor2s3 U579 ( .DIN1(n590), .DIN2(n1390), .Q(g7815) );
  xor2s3 U580 ( .DIN1(n2626), .DIN2(n2627), .Q(n1390) );
  nor2s3 U581 ( .DIN1(n778), .DIN2(n1391), .Q(g7814) );
  xor2s3 U582 ( .DIN1(n836), .DIN2(n530), .Q(n1391) );
  and3s3 U583 ( .DIN1(n530), .DIN2(n2061), .DIN3(n1392), .Q(g7813) );
  nnd2s3 U584 ( .DIN1(n1984), .DIN2(n1393), .Q(n1392) );
  nor2s3 U585 ( .DIN1(n1393), .DIN2(n1984), .Q(n1357) );
  and2s3 U586 ( .DIN1(n1394), .DIN2(n2061), .Q(g7812) );
  nnd2s3 U587 ( .DIN1(n1395), .DIN2(n1396), .Q(n1394) );
  nnd3s3 U588 ( .DIN1(n1397), .DIN2(n722), .DIN3(n645), .Q(n1396) );
  nnd2s3 U589 ( .DIN1(n1393), .DIN2(n532), .Q(n1395) );
  or2s3 U590 ( .DIN1(n1398), .DIN2(n1397), .Q(n1393) );
  nor2s3 U591 ( .DIN1(n778), .DIN2(n1399), .Q(g7811) );
  xor2s3 U592 ( .DIN1(n2620), .DIN2(n645), .Q(n1399) );
  nnd2s3 U593 ( .DIN1(n1401), .DIN2(n2061), .Q(g7810) );
  nnd2s3 U594 ( .DIN1(n1402), .DIN2(n1400), .Q(n1401) );
  nnd2s3 U595 ( .DIN1(n646), .DIN2(n813), .Q(n1400) );
  nnd2s3 U596 ( .DIN1(n2619), .DIN2(n1398), .Q(n1402) );
  and3s3 U597 ( .DIN1(n1403), .DIN2(n575), .DIN3(g109), .Q(g7809) );
  nnd2s3 U598 ( .DIN1(\DFF_452/net739 ), .DIN2(n708), .Q(n1403) );
  nnd2s3 U599 ( .DIN1(n1404), .DIN2(n1405), .Q(g7808) );
  or2s3 U600 ( .DIN1(n2849), .DIN2(n2652), .Q(n1405) );
  nnd2s3 U601 ( .DIN1(n2849), .DIN2(n782), .Q(n1404) );
  nnd2s3 U602 ( .DIN1(n1406), .DIN2(n1407), .Q(g7807) );
  or2s3 U603 ( .DIN1(n2849), .DIN2(n2647), .Q(n1407) );
  nnd2s3 U604 ( .DIN1(n2849), .DIN2(n822), .Q(n1406) );
  nnd2s3 U605 ( .DIN1(n1408), .DIN2(n1409), .Q(g7806) );
  or2s3 U606 ( .DIN1(n2849), .DIN2(n2650), .Q(n1409) );
  nnd2s3 U607 ( .DIN1(n2849), .DIN2(n839), .Q(n1408) );
  nnd2s3 U608 ( .DIN1(n1410), .DIN2(n1411), .Q(g7805) );
  or2s3 U609 ( .DIN1(n2849), .DIN2(n2651), .Q(n1411) );
  nnd2s3 U610 ( .DIN1(n2849), .DIN2(n863), .Q(n1410) );
  nnd2s3 U611 ( .DIN1(n1412), .DIN2(n1413), .Q(g7804) );
  or2s3 U612 ( .DIN1(n2849), .DIN2(n2655), .Q(n1413) );
  nnd2s3 U613 ( .DIN1(n2849), .DIN2(n707), .Q(n1412) );
  nnd2s3 U614 ( .DIN1(n1414), .DIN2(n1415), .Q(g7803) );
  or2s3 U615 ( .DIN1(n2849), .DIN2(n2649), .Q(n1415) );
  nnd2s3 U616 ( .DIN1(n2849), .DIN2(n818), .Q(n1414) );
  nnd2s3 U617 ( .DIN1(n1416), .DIN2(n1417), .Q(g7802) );
  or2s3 U618 ( .DIN1(n2849), .DIN2(n2648), .Q(n1417) );
  nnd2s3 U619 ( .DIN1(n2849), .DIN2(n630), .Q(n1416) );
  nnd2s3 U620 ( .DIN1(n1418), .DIN2(n1419), .Q(g7801) );
  or2s3 U621 ( .DIN1(n2849), .DIN2(n2654), .Q(n1419) );
  nnd2s3 U622 ( .DIN1(n2849), .DIN2(n779), .Q(n1418) );
  nnd2s3 U623 ( .DIN1(n1420), .DIN2(n1421), .Q(g7800) );
  nnd2s3 U624 ( .DIN1(n2853), .DIN2(n743), .Q(n1421) );
  nnd2s3 U625 ( .DIN1(n2849), .DIN2(n857), .Q(n1420) );
  nnd2s3 U626 ( .DIN1(n1422), .DIN2(n1423), .Q(g7799) );
  or2s3 U627 ( .DIN1(n2849), .DIN2(n2653), .Q(n1423) );
  nnd2s3 U628 ( .DIN1(n2848), .DIN2(n705), .Q(n1422) );
  nnd2s3 U629 ( .DIN1(n1424), .DIN2(n1425), .Q(g7798) );
  nnd2s3 U630 ( .DIN1(n2853), .DIN2(n621), .Q(n1425) );
  nnd2s3 U631 ( .DIN1(n2848), .DIN2(n642), .Q(n1424) );
  and3s3 U632 ( .DIN1(n1426), .DIN2(n1342), .DIN3(n695), .Q(g7786) );
  nnd3s3 U633 ( .DIN1(n635), .DIN2(n802), .DIN3(n1427), .Q(n1342) );
  nnd2s3 U634 ( .DIN1(n2050), .DIN2(n1428), .Q(n1426) );
  nnd2s3 U635 ( .DIN1(n1427), .DIN2(n802), .Q(n1428) );
  and3s3 U636 ( .DIN1(n1429), .DIN2(n1345), .DIN3(n841), .Q(g7785) );
  or3s3 U637 ( .DIN1(n2057), .DIN2(n2557), .DIN3(n1430), .Q(n1345) );
  nnd2s3 U638 ( .DIN1(n2057), .DIN2(n1431), .Q(n1429) );
  or2s3 U639 ( .DIN1(n1430), .DIN2(n2557), .Q(n1431) );
  nnd2s3 U640 ( .DIN1(n2034), .DIN2(n1432), .Q(g7784) );
  nor2s3 U641 ( .DIN1(n2018), .DIN2(n608), .Q(g7783) );
  nnd2s3 U642 ( .DIN1(n2035), .DIN2(n1432), .Q(g7782) );
  nor2s3 U643 ( .DIN1(n2019), .DIN2(n608), .Q(g7781) );
  nnd2s3 U644 ( .DIN1(n2036), .DIN2(n1432), .Q(g7780) );
  nor2s3 U645 ( .DIN1(n2020), .DIN2(n608), .Q(g7779) );
  nnd2s3 U646 ( .DIN1(n2037), .DIN2(n1432), .Q(g7778) );
  nor2s3 U647 ( .DIN1(n2021), .DIN2(n608), .Q(g7777) );
  nor2s3 U648 ( .DIN1(n2022), .DIN2(n608), .Q(g7776) );
  nor2s3 U649 ( .DIN1(n2023), .DIN2(n608), .Q(g7775) );
  nnd2s3 U650 ( .DIN1(n2038), .DIN2(n1432), .Q(g7774) );
  nnd2s3 U651 ( .DIN1(n1433), .DIN2(n1434), .Q(g7773) );
  or2s3 U652 ( .DIN1(n1435), .DIN2(n2733), .Q(n1434) );
  or2s3 U653 ( .DIN1(n574), .DIN2(n1925), .Q(n1433) );
  nnd2s3 U654 ( .DIN1(n1436), .DIN2(n1437), .Q(g7772) );
  or2s3 U655 ( .DIN1(n1435), .DIN2(n2745), .Q(n1437) );
  nnd2s3 U656 ( .DIN1(n1435), .DIN2(n749), .Q(n1436) );
  nnd2s3 U657 ( .DIN1(n1438), .DIN2(n1439), .Q(g7771) );
  or2s3 U658 ( .DIN1(n1435), .DIN2(n2754), .Q(n1439) );
  or2s3 U659 ( .DIN1(n574), .DIN2(n1938), .Q(n1438) );
  nnd2s3 U660 ( .DIN1(n1440), .DIN2(n1441), .Q(g7770) );
  or2s3 U661 ( .DIN1(n1435), .DIN2(n2768), .Q(n1441) );
  or2s3 U662 ( .DIN1(n574), .DIN2(n1961), .Q(n1440) );
  nnd2s3 U663 ( .DIN1(n1442), .DIN2(n1443), .Q(g7769) );
  or2s3 U664 ( .DIN1(n1435), .DIN2(n2780), .Q(n1443) );
  or2s3 U665 ( .DIN1(n574), .DIN2(n1996), .Q(n1442) );
  nnd2s3 U666 ( .DIN1(n1444), .DIN2(n1445), .Q(g7768) );
  or2s3 U667 ( .DIN1(n1435), .DIN2(n2794), .Q(n1445) );
  or2s3 U668 ( .DIN1(n574), .DIN2(n1960), .Q(n1444) );
  nnd2s3 U669 ( .DIN1(n1446), .DIN2(n1447), .Q(g7767) );
  or2s3 U670 ( .DIN1(n1435), .DIN2(n2804), .Q(n1447) );
  nnd2s3 U671 ( .DIN1(n1435), .DIN2(n688), .Q(n1446) );
  nnd2s3 U672 ( .DIN1(n1448), .DIN2(n1449), .Q(g7766) );
  or2s3 U673 ( .DIN1(n1435), .DIN2(n2815), .Q(n1449) );
  nnd2s3 U674 ( .DIN1(n1435), .DIN2(n814), .Q(n1448) );
  nnd2s3 U675 ( .DIN1(n1450), .DIN2(n1451), .Q(g7765) );
  nnd2s3 U676 ( .DIN1(n574), .DIN2(n847), .Q(n1451) );
  or2s3 U677 ( .DIN1(n574), .DIN2(n1959), .Q(n1450) );
  nnd2s3 U678 ( .DIN1(n1452), .DIN2(n1453), .Q(g7764) );
  nnd2s3 U679 ( .DIN1(n574), .DIN2(n636), .Q(n1453) );
  or2s3 U680 ( .DIN1(n574), .DIN2(n1992), .Q(n1452) );
  nnd2s3 U681 ( .DIN1(n1454), .DIN2(n1455), .Q(g7763) );
  or2s3 U682 ( .DIN1(n1435), .DIN2(n2753), .Q(n1455) );
  nnd2s3 U683 ( .DIN1(n1435), .DIN2(n792), .Q(n1454) );
  nnd2s3 U684 ( .DIN1(n1456), .DIN2(n1457), .Q(g7762) );
  or2s3 U685 ( .DIN1(n1435), .DIN2(n2767), .Q(n1457) );
  or2s3 U686 ( .DIN1(n574), .DIN2(n1926), .Q(n1456) );
  nnd2s3 U687 ( .DIN1(n1458), .DIN2(n1459), .Q(g7761) );
  or2s3 U688 ( .DIN1(n1435), .DIN2(n2779), .Q(n1459) );
  or2s3 U689 ( .DIN1(n574), .DIN2(n2521), .Q( tempn1458 ) );
  nnd2s3 U690 ( .DIN1(n1460), .DIN2(n1461), .Q(g7760) );
  or2s3 U691 ( .DIN1(n1435), .DIN2(n2793), .Q(n1461) );
  nnd2s3 U692 ( .DIN1(n1435), .DIN2(n656), .Q(n1460) );
  nnd2s3 U693 ( .DIN1(g109), .DIN2(n1462), .Q(n1435) );
  nnd2s3 U694 ( .DIN1(n2017), .DIN2(n1353), .Q(n1462) );
  nnd2s3 U695 ( .DIN1(n1463), .DIN2(n1464), .Q(g7759) );
  nnd2s3 U696 ( .DIN1(n2861), .DIN2(n753), .Q(n1464) );
  nnd2s3 U697 ( .DIN1(n1465), .DIN2(n1466), .Q(g7758) );
  nnd2s3 U698 ( .DIN1(n2861), .DIN2(n784), .Q(n1466) );
  nnd2s3 U699 ( .DIN1(n1144), .DIN2(n1467), .Q(g7757) );
  nnd2s3 U700 ( .DIN1(n2862), .DIN2(n529), .Q(n1467) );
  nnd2s3 U701 ( .DIN1(n1152), .DIN2(n1468), .Q(g7756) );
  nnd2s3 U702 ( .DIN1(n2862), .DIN2(n709), .Q(n1468) );
  nnd2s3 U703 ( .DIN1(n1160), .DIN2(n1469), .Q(g7755) );
  nnd2s3 U704 ( .DIN1(n2862), .DIN2(n756), .Q(n1469) );
  nnd2s3 U705 ( .DIN1(n1169), .DIN2(n1470), .Q(g7754) );
  nnd2s3 U706 ( .DIN1(n2862), .DIN2(n729), .Q(n1470) );
  nnd2s3 U707 ( .DIN1(g2355), .DIN2(n803), .Q(n1169) );
  nnd2s3 U708 ( .DIN1(n1173), .DIN2(n1471), .Q(g7753) );
  nnd2s3 U709 ( .DIN1(n2862), .DIN2(n771), .Q(n1471) );
  nnd2s3 U710 ( .DIN1(g2355), .DIN2(n677), .Q(n1173) );
  nnd2s3 U711 ( .DIN1(n1180), .DIN2(n1472), .Q(g7752) );
  nnd2s3 U712 ( .DIN1(n2862), .DIN2(n844), .Q(n1472) );
  nnd2s3 U713 ( .DIN1(g2355), .DIN2(n868), .Q(n1180) );
  nnd2s3 U714 ( .DIN1(n1473), .DIN2(n1474), .Q(g7751) );
  nnd2s3 U715 ( .DIN1(n2862), .DIN2(n786), .Q(n1474) );
  nnd2s3 U716 ( .DIN1(n1187), .DIN2(n1475), .Q(g7750) );
  nnd2s3 U717 ( .DIN1(n2862), .DIN2(n582), .Q(n1475) );
  nor2s3 U718 ( .DIN1(n2870), .DIN2(n2521), .Q(g7749) );
  nnd2s3 U719 ( .DIN1(n1476), .DIN2(n1477), .Q(g7746) );
  nnd2s3 U720 ( .DIN1(g7748), .DIN2(n1478), .Q(n1477) );
  xor2s3 U721 ( .DIN1(n1925), .DIN2(n1479), .Q(n1478) );
  nor2s3 U722 ( .DIN1(n2870), .DIN2(n1926), .Q(g7748) );
  nnd2s3 U723 ( .DIN1(n1926), .DIN2(n1480), .Q(n1476) );
  nnd2s3 U724 ( .DIN1(n1481), .DIN2(n1482), .Q(n1480) );
  nnd3s3 U725 ( .DIN1(g109), .DIN2(n1479), .DIN3(n1925), .Q(n1482) );
  nnd2s3 U726 ( .DIN1(g7747), .DIN2(n655), .Q(n1481) );
  xnr2s3 U727 ( .DIN1(n656), .DIN2(n1937), .Q(n1479) );
  nor2s3 U728 ( .DIN1(n2870), .DIN2(n1925), .Q(g7747) );
  nnd2s3 U729 ( .DIN1(n1483), .DIN2(n1484), .Q(g7745) );
  nnd2s3 U730 ( .DIN1(g109), .DIN2(n639), .Q(n1484) );
  or2s3 U731 ( .DIN1(g4906), .DIN2(n2627), .Q(g7366) );
  nnd2s3 U732 ( .DIN1(n1485), .DIN2(n1486), .Q(g7365) );
  nnd2s3 U733 ( .DIN1(n2840), .DIN2(n795), .Q(n1486) );
  nnd2s3 U734 ( .DIN1(n2845), .DIN2(n572), .Q(n1485) );
  nnd2s3 U735 ( .DIN1(n1488), .DIN2(n1489), .Q(g7364) );
  nnd2s3 U736 ( .DIN1(n2840), .DIN2(n851), .Q(n1489) );
  nnd2s3 U737 ( .DIN1(n2844), .DIN2(n823), .Q(n1488) );
  nnd2s3 U738 ( .DIN1(n1490), .DIN2(n1491), .Q(g7363) );
  nnd2s3 U739 ( .DIN1(n2840), .DIN2(n555), .Q(n1491) );
  or2s3 U740 ( .DIN1(n2842), .DIN2(n2755), .Q(n1490) );
  nnd2s3 U741 ( .DIN1(n1492), .DIN2(n1493), .Q(g7362) );
  nnd2s3 U742 ( .DIN1(n2840), .DIN2(n846), .Q(n1493) );
  or2s3 U743 ( .DIN1(n2842), .DIN2(n2769), .Q(n1492) );
  nnd2s3 U744 ( .DIN1(n1494), .DIN2(n1495), .Q(g7361) );
  nnd2s3 U745 ( .DIN1(n2840), .DIN2(n742), .Q(n1495) );
  nnd2s3 U746 ( .DIN1(n2844), .DIN2(n612), .Q(n1494) );
  nnd2s3 U747 ( .DIN1(n1496), .DIN2(n1497), .Q(g7360) );
  or2s3 U748 ( .DIN1(n2847), .DIN2(n2526), .Q(n1497) );
  or2s3 U749 ( .DIN1(n2842), .DIN2(n2798), .Q(n1496) );
  nnd2s3 U750 ( .DIN1(n1498), .DIN2(n1499), .Q(g7359) );
  nnd2s3 U751 ( .DIN1(n2840), .DIN2(n801), .Q(n1499) );
  or2s3 U752 ( .DIN1(n2842), .DIN2(n2802), .Q(n1498) );
  nnd2s3 U753 ( .DIN1(n1500), .DIN2(n1501), .Q(g7358) );
  nnd2s3 U754 ( .DIN1(n2840), .DIN2(n810), .Q(n1501) );
  nnd2s3 U755 ( .DIN1(n2844), .DIN2(n578), .Q(n1500) );
  nnd2s3 U756 ( .DIN1(n1502), .DIN2(n1503), .Q(g7357) );
  nnd2s3 U757 ( .DIN1(n2840), .DIN2(n859), .Q(n1503) );
  nnd2s3 U758 ( .DIN1(n2844), .DIN2(n732), .Q(n1502) );
  nnd2s3 U759 ( .DIN1(n1504), .DIN2(n1505), .Q(g7356) );
  nnd2s3 U760 ( .DIN1(n2840), .DIN2(n783), .Q(n1505) );
  nnd2s3 U761 ( .DIN1(n2844), .DIN2(n861), .Q(n1504) );
  nnd2s3 U762 ( .DIN1(n1506), .DIN2(n1507), .Q(g7355) );
  nnd2s3 U763 ( .DIN1(n2840), .DIN2(n819), .Q(n1507) );
  or2s3 U764 ( .DIN1(n2841), .DIN2(n2756), .Q(n1506) );
  nnd2s3 U765 ( .DIN1(n1508), .DIN2(n1509), .Q(g7354) );
  nnd2s3 U766 ( .DIN1(n2840), .DIN2(n559), .Q(n1509) );
  or2s3 U767 ( .DIN1(n2841), .DIN2(n2770), .Q(n1508) );
  nnd2s3 U768 ( .DIN1(n1510), .DIN2(n1511), .Q(g7353) );
  or2s3 U769 ( .DIN1(n2846), .DIN2(n2537), .Q(n1511) );
  nnd2s3 U770 ( .DIN1(n2845), .DIN2(n796), .Q(n1510) );
  nnd2s3 U771 ( .DIN1(n1512), .DIN2(n1513), .Q(g7352) );
  nnd2s3 U772 ( .DIN1(n2840), .DIN2(n805), .Q(n1513) );
  or2s3 U773 ( .DIN1(n2841), .DIN2(n2795), .Q(n1512) );
  nnd2s3 U774 ( .DIN1(n1514), .DIN2(n1515), .Q(g7351) );
  nnd2s3 U775 ( .DIN1(n2841), .DIN2(n741), .Q(n1515) );
  nnd2s3 U776 ( .DIN1(n2845), .DIN2(n800), .Q(n1514) );
  nnd2s3 U777 ( .DIN1(n1516), .DIN2(n1517), .Q(g7350) );
  or2s3 U778 ( .DIN1(n2846), .DIN2(n1991), .Q(n1517) );
  nnd2s3 U779 ( .DIN1(n2845), .DIN2(n730), .Q(n1516) );
  nnd2s3 U780 ( .DIN1(n1518), .DIN2(n1519), .Q(g7349) );
  nnd2s3 U781 ( .DIN1(n2840), .DIN2(n694), .Q(n1519) );
  or2s3 U782 ( .DIN1(n2841), .DIN2(n2759), .Q(n1518) );
  nnd2s3 U783 ( .DIN1(n1520), .DIN2(n1521), .Q(g7348) );
  or2s3 U784 ( .DIN1(n2846), .DIN2(n2529), .Q(n1521) );
  or2s3 U785 ( .DIN1(n2841), .DIN2(n2772), .Q(n1520) );
  nnd2s3 U786 ( .DIN1(n1522), .DIN2(n1523), .Q(g7347) );
  nnd2s3 U787 ( .DIN1(n2841), .DIN2(n816), .Q(n1523) );
  or2s3 U788 ( .DIN1(n2842), .DIN2(n2783), .Q(n1522) );
  nnd2s3 U789 ( .DIN1(n1524), .DIN2(n1525), .Q(g7346) );
  nnd2s3 U790 ( .DIN1(n2841), .DIN2(n780), .Q(n1525) );
  or2s3 U791 ( .DIN1(n2841), .DIN2(n2797), .Q(n1524) );
  nnd2s3 U792 ( .DIN1(n1526), .DIN2(n1527), .Q(g7345) );
  nnd2s3 U793 ( .DIN1(n2841), .DIN2(n719), .Q(n1527) );
  or2s3 U794 ( .DIN1(n2842), .DIN2(n2805), .Q(n1526) );
  nnd2s3 U795 ( .DIN1(n1528), .DIN2(n1529), .Q(g7344) );
  or2s3 U796 ( .DIN1(n2846), .DIN2(n2533), .Q(n1529) );
  or2s3 U797 ( .DIN1(n2842), .DIN2(n2814), .Q(n1528) );
  nnd2s3 U798 ( .DIN1(n1530), .DIN2(n1531), .Q(g7343) );
  or2s3 U799 ( .DIN1(n2846), .DIN2(n2534), .Q(n1531) );
  nnd2s3 U800 ( .DIN1(n2845), .DIN2(n680), .Q(n1530) );
  nnd2s3 U801 ( .DIN1(n1532), .DIN2(n1533), .Q(g7342) );
  nnd2s3 U802 ( .DIN1(n2841), .DIN2(n603), .Q(n1533) );
  nnd2s3 U803 ( .DIN1(n2846), .DIN2(n611), .Q(n1532) );
  nnd2s3 U804 ( .DIN1(n1534), .DIN2(n1535), .Q(g7341) );
  nnd2s3 U805 ( .DIN1(n2841), .DIN2(n536), .Q(n1535) );
  or2s3 U806 ( .DIN1(n2842), .DIN2(n2758), .Q(n1534) );
  nnd2s3 U807 ( .DIN1(n1536), .DIN2(n1537), .Q(g7340) );
  nnd2s3 U808 ( .DIN1(n2841), .DIN2(n852), .Q(n1537) );
  or2s3 U809 ( .DIN1(n2842), .DIN2(n2771), .Q(n1536) );
  nnd2s3 U810 ( .DIN1(n1538), .DIN2(n1539), .Q(g7339) );
  or2s3 U811 ( .DIN1(n2847), .DIN2(n2541), .Q(n1539) );
  or2s3 U812 ( .DIN1(n2842), .DIN2(n2785), .Q(n1538) );
  nnd2s3 U813 ( .DIN1(n1540), .DIN2(n1541), .Q(g7338) );
  nnd2s3 U814 ( .DIN1(n2841), .DIN2(n763), .Q(n1541) );
  or2s3 U815 ( .DIN1(n2842), .DIN2(n2799), .Q(n1540) );
  nnd2s3 U816 ( .DIN1(g109), .DIN2(n1363), .Q(n1487) );
  nnd2s3 U817 ( .DIN1(n2776), .DIN2(n1353), .Q(n1363) );
  nnd2s3 U818 ( .DIN1(n1483), .DIN2(n1542), .Q(g7337) );
  nnd2s3 U819 ( .DIN1(g109), .DIN2(n524), .Q(n1542) );
  nnd2s3 U820 ( .DIN1(n1483), .DIN2(n1543), .Q(g7336) );
  nnd2s3 U821 ( .DIN1(g109), .DIN2(n775), .Q(n1543) );
  nnd2s3 U822 ( .DIN1(n1353), .DIN2(g109), .Q(n1483) );
  nor2s3 U823 ( .DIN1(n575), .DIN2(n2861), .Q(n1353) );
  nor2s3 U824 ( .DIN1(n2870), .DIN2(n2537), .Q(g7335) );
  nor2s3 U825 ( .DIN1(n2589), .DIN2(n2868), .Q(g7334) );
  nor2s3 U826 ( .DIN1(n2587), .DIN2(n2868), .Q(g7333) );
  nor2s3 U827 ( .DIN1(n2538), .DIN2(n2868), .Q(g7332) );
  nor2s3 U828 ( .DIN1(n2539), .DIN2(n2868), .Q(g7331) );
  nor2s3 U829 ( .DIN1(n2540), .DIN2(n2868), .Q(g7330) );
  nor2s3 U830 ( .DIN1(n2870), .DIN2(n2541), .Q(g7329) );
  nor2s3 U831 ( .DIN1(n2543), .DIN2(n2868), .Q(g7328) );
  nnd2s3 U832 ( .DIN1(n1544), .DIN2(n1545), .Q(g7326) );
  or3s3 U833 ( .DIN1(n1546), .DIN2(n2871), .DIN3(n741), .Q(n1545) );
  nnd2s3 U834 ( .DIN1(g7327), .DIN2(n1546), .Q(n1544) );
  xnr2s3 U835 ( .DIN1(n763), .DIN2(n1547), .Q(n1546) );
  xor2s3 U836 ( .DIN1(n2542), .DIN2(n2543), .Q(n1547) );
  nor2s3 U837 ( .DIN1(n2870), .DIN2(n2012), .Q(g7327) );
  and2s3 U838 ( .DIN1(g109), .DIN2(n2546), .Q(g7325) );
  nor2s3 U839 ( .DIN1(n1963), .DIN2(n2868), .Q(g7324) );
  nor2s3 U840 ( .DIN1(n2555), .DIN2(n2867), .Q(g7323) );
  nor2s3 U841 ( .DIN1(n1946), .DIN2(n2867), .Q(g7322) );
  nor2s3 U842 ( .DIN1(n906), .DIN2(n708), .Q(g7321) );
  nnd2s3 U843 ( .DIN1(g6825), .DIN2(n1548), .Q(n906) );
  nor2s3 U844 ( .DIN1(n2550), .DIN2(n2867), .Q(g7319) );
  nor2s3 U845 ( .DIN1(n2041), .DIN2(n2867), .Q(g7318) );
  and2s3 U846 ( .DIN1(g109), .DIN2(n2552), .Q(g7317) );
  nor2s3 U847 ( .DIN1(n2001), .DIN2(n2867), .Q(g7316) );
  and2s3 U848 ( .DIN1(g109), .DIN2(n2553), .Q(g7315) );
  nor2s3 U849 ( .DIN1(n1962), .DIN2(n2867), .Q(g7314) );
  and2s3 U850 ( .DIN1(g109), .DIN2(n2551), .Q(g7313) );
  nor2s3 U851 ( .DIN1(n1972), .DIN2(n2867), .Q(g7312) );
  nor2s3 U852 ( .DIN1(n2040), .DIN2(n2867), .Q(g7311) );
  and2s3 U853 ( .DIN1(g109), .DIN2(n2548), .Q(g7310) );
  and2s3 U854 ( .DIN1(g109), .DIN2(n2547), .Q(g7309) );
  nor2s3 U855 ( .DIN1(n1947), .DIN2(n2867), .Q(g7308) );
  nor2s3 U856 ( .DIN1(n1939), .DIN2(n2867), .Q(g7307) );
  nor2s3 U857 ( .DIN1(n2549), .DIN2(n2866), .Q(g7306) );
  nor2s3 U858 ( .DIN1(n2002), .DIN2(n2867), .Q(g7305) );
  nnd2s3 U859 ( .DIN1(n1549), .DIN2(n1550), .Q(g7304) );
  nnd2s3 U860 ( .DIN1(g6836), .DIN2(n1551), .Q(n1550) );
  xor2s3 U861 ( .DIN1(n1995), .DIN2(n564), .Q(n1551) );
  nnd2s3 U862 ( .DIN1(n1552), .DIN2(n613), .Q(n1549) );
  nnd2s3 U863 ( .DIN1(n1553), .DIN2(n1554), .Q(n1552) );
  nnd3s3 U864 ( .DIN1(g109), .DIN2(n564), .DIN3(n1995), .Q(n1554) );
  nnd2s3 U865 ( .DIN1(n1555), .DIN2(g6825), .Q(n1553) );
  xor2s3 U866 ( .DIN1(n1556), .DIN2(n2559), .Q(n1555) );
  nnd2s3 U867 ( .DIN1(n2554), .DIN2(n1557), .Q(n1556) );
  nnd2s3 U868 ( .DIN1(n1995), .DIN2(n1548), .Q(n1557) );
  and4s2 U869 ( .DIN1(n633), .DIN2(n1558), .DIN3(n1559), .DIN4(n1560), .Q(
        n1548) );
  nor6s3 U870 ( .DIN1(n2548), .DIN2(n2546), .DIN3(n2547), .DIN4(n2553), .DIN5(
        n2551), .DIN6(n2552), .Q(n1560) );
  nor6s3 U871 ( .DIN1(n697), .DIN2(n2560), .DIN3(n2561), .DIN4(n677), .DIN5(
        n712), .DIN6(n772), .Q(n1559) );
  nor6s3 U872 ( .DIN1(n868), .DIN2(n827), .DIN3(n803), .DIN4(n811), .DIN5(n853), .DIN6(n799), .Q(n1558) );
  nnd2s3 U873 ( .DIN1(n1562), .DIN2(n1563), .Q(g7303) );
  nnd2s3 U874 ( .DIN1(n1564), .DIN2(n685), .Q(n1563) );
  nnd2s3 U875 ( .DIN1(n649), .DIN2(n837), .Q(n1562) );
  nnd2s3 U876 ( .DIN1(n1565), .DIN2(n1566), .Q(g7302) );
  nnd2s3 U877 ( .DIN1(n1564), .DIN2(n837), .Q(n1566) );
  nnd2s3 U878 ( .DIN1(n649), .DIN2(n599), .Q(n1565) );
  nnd2s3 U879 ( .DIN1(n1567), .DIN2(n1568), .Q(g7301) );
  nnd2s3 U880 ( .DIN1(n1564), .DIN2(n599), .Q(n1568) );
  nnd2s3 U881 ( .DIN1(n649), .DIN2(n664), .Q(n1567) );
  nnd2s3 U882 ( .DIN1(n1569), .DIN2(n1570), .Q(g7300) );
  nnd2s3 U883 ( .DIN1(n1564), .DIN2(n664), .Q(n1570) );
  nnd2s3 U884 ( .DIN1(n649), .DIN2(n745), .Q(n1569) );
  nnd2s3 U885 ( .DIN1(n1571), .DIN2(n1572), .Q(g7299) );
  nnd2s3 U886 ( .DIN1(n1564), .DIN2(n745), .Q(n1572) );
  nnd2s3 U887 ( .DIN1(n649), .DIN2(n674), .Q(n1571) );
  nnd2s3 U888 ( .DIN1(n1573), .DIN2(n1574), .Q(g7298) );
  nnd2s3 U889 ( .DIN1(n1564), .DIN2(n674), .Q(n1574) );
  nnd2s3 U890 ( .DIN1(n649), .DIN2(n762), .Q(n1573) );
  nnd2s3 U891 ( .DIN1(n1575), .DIN2(n1576), .Q(g7297) );
  nnd2s3 U892 ( .DIN1(n1564), .DIN2(n762), .Q(n1576) );
  nnd2s3 U893 ( .DIN1(n649), .DIN2(n548), .Q(n1575) );
  nnd2s3 U894 ( .DIN1(n1577), .DIN2(n1578), .Q(g7296) );
  nnd2s3 U895 ( .DIN1(n1564), .DIN2(n548), .Q(n1578) );
  nnd2s3 U896 ( .DIN1(n649), .DIN2(n570), .Q(n1577) );
  nnd2s3 U897 ( .DIN1(n1579), .DIN2(n1580), .Q(g7295) );
  nnd2s3 U898 ( .DIN1(n1564), .DIN2(n631), .Q(n1580) );
  nnd2s3 U899 ( .DIN1(n649), .DIN2(n566), .Q(n1579) );
  nnd2s3 U900 ( .DIN1(n1581), .DIN2(n1582), .Q(g7294) );
  nnd2s3 U901 ( .DIN1(n1564), .DIN2(n566), .Q(n1582) );
  nnd2s3 U902 ( .DIN1(n649), .DIN2(n734), .Q(n1581) );
  nnd2s3 U903 ( .DIN1(n1583), .DIN2(n1584), .Q(g7293) );
  nnd2s3 U904 ( .DIN1(n1564), .DIN2(n734), .Q(n1584) );
  nnd2s3 U905 ( .DIN1(n649), .DIN2(n834), .Q(n1583) );
  nnd2s3 U906 ( .DIN1(n1585), .DIN2(n1586), .Q(g7292) );
  nnd2s3 U907 ( .DIN1(n1564), .DIN2(n834), .Q(n1586) );
  nnd2s3 U908 ( .DIN1(n649), .DIN2(n557), .Q(n1585) );
  nnd2s3 U909 ( .DIN1(n1587), .DIN2(n1588), .Q(g7291) );
  nnd2s3 U910 ( .DIN1(n1564), .DIN2(n557), .Q(n1588) );
  nnd2s3 U911 ( .DIN1(n649), .DIN2(n854), .Q(n1587) );
  nnd2s3 U912 ( .DIN1(n1589), .DIN2(n1590), .Q(g7290) );
  nnd2s3 U913 ( .DIN1(n1564), .DIN2(n854), .Q(n1590) );
  nnd2s3 U914 ( .DIN1(n649), .DIN2(n685), .Q(n1589) );
  nor2s3 U915 ( .DIN1(n1229), .DIN2(n1591), .Q(g7289) );
  xor2s3 U916 ( .DIN1(n2556), .DIN2(n1427), .Q(n1591) );
  nor2s3 U917 ( .DIN1(n1280), .DIN2(n1592), .Q(g7288) );
  xnr2s3 U918 ( .DIN1(n2557), .DIN2(n1430), .Q(n1592) );
  or2s3 U919 ( .DIN1(g4894), .DIN2(n2558), .Q(g7287) );
  nor2s3 U920 ( .DIN1(n706), .DIN2(n1593), .Q(g7285) );
  nor2s3 U921 ( .DIN1(n2870), .DIN2(n905), .Q(n1593) );
  nor2s3 U922 ( .DIN1(n2727), .DIN2(n646), .Q(g6845) );
  nnd2s3 U923 ( .DIN1(n1594), .DIN2(n1595), .Q(g6844) );
  nnd2s3 U925 ( .DIN1(g4907), .DIN2(n718), .Q(n1594) );
  nor3s3 U926 ( .DIN1(n2848), .DIN2(g4901), .DIN3(n1596), .Q(g6843) );
  nor2s3 U927 ( .DIN1(g1696), .DIN2(g4901), .Q(g6842) );
  nor2s3 U928 ( .DIN1(n2559), .DIN2(n2866), .Q(g6837) );
  nor2s3 U929 ( .DIN1(n613), .DIN2(n2866), .Q(g6836) );
  and2s3 U930 ( .DIN1(g109), .DIN2(n2561), .Q(g6835) );
  nor2s3 U931 ( .DIN1(n2870), .DIN2(n1995), .Q(g6825) );
  nor2s3 U932 ( .DIN1(n679), .DIN2(n1597), .Q(g6818) );
  nor2s3 U933 ( .DIN1(n2011), .DIN2(n2866), .Q(n1597) );
  nor2s3 U934 ( .DIN1(n1949), .DIN2(n1598), .Q(g6817) );
  nor2s3 U935 ( .DIN1(n1929), .DIN2(n1598), .Q(g6816) );
  nor2s3 U936 ( .DIN1(n1976), .DIN2(n1598), .Q(g6815) );
  nor2s3 U937 ( .DIN1(n1974), .DIN2(n1598), .Q(g6814) );
  nnd2s3 U938 ( .DIN1(g109), .DIN2(\DFF_126/net413 ), .Q(n1598) );
  nnd2s3 U939 ( .DIN1(n1599), .DIN2(n1600), .Q(g6813) );
  nnd2s3 U940 ( .DIN1(n1601), .DIN2(n746), .Q(n1600) );
  nnd2s3 U941 ( .DIN1(n650), .DIN2(n782), .Q(n1599) );
  nnd2s3 U942 ( .DIN1(n1602), .DIN2(n1603), .Q(g6812) );
  nnd2s3 U943 ( .DIN1(n1601), .DIN2(n693), .Q(n1603) );
  nnd2s3 U944 ( .DIN1(n650), .DIN2(n822), .Q(n1602) );
  nnd2s3 U945 ( .DIN1(n1604), .DIN2(n1605), .Q(g6811) );
  nnd2s3 U946 ( .DIN1(n1601), .DIN2(n740), .Q(n1605) );
  nnd2s3 U947 ( .DIN1(n650), .DIN2(n839), .Q(n1604) );
  nnd2s3 U948 ( .DIN1(n1606), .DIN2(n1607), .Q(g6810) );
  nnd2s3 U949 ( .DIN1(n1601), .DIN2(n713), .Q(n1607) );
  nnd2s3 U950 ( .DIN1(n650), .DIN2(n863), .Q(n1606) );
  nnd2s3 U951 ( .DIN1(n1608), .DIN2(n1609), .Q(g6809) );
  nnd2s3 U952 ( .DIN1(n1601), .DIN2(n751), .Q(n1609) );
  nnd2s3 U953 ( .DIN1(n650), .DIN2(n707), .Q(n1608) );
  nnd2s3 U954 ( .DIN1(n1610), .DIN2(n1611), .Q(g6808) );
  nnd2s3 U955 ( .DIN1(n1601), .DIN2(n831), .Q(n1611) );
  nnd2s3 U956 ( .DIN1(n650), .DIN2(n818), .Q(n1610) );
  nnd2s3 U957 ( .DIN1(n1612), .DIN2(n1613), .Q(g6807) );
  nnd2s3 U958 ( .DIN1(n1601), .DIN2(n824), .Q(n1613) );
  nnd2s3 U959 ( .DIN1(n650), .DIN2(n630), .Q(n1612) );
  nnd2s3 U960 ( .DIN1(n1614), .DIN2(n1615), .Q(g6806) );
  nnd2s3 U961 ( .DIN1(n1601), .DIN2(n601), .Q(n1615) );
  nnd2s3 U962 ( .DIN1(n650), .DIN2(n779), .Q(n1614) );
  nnd2s3 U963 ( .DIN1(n1616), .DIN2(n1617), .Q(g6805) );
  nnd2s3 U964 ( .DIN1(n1601), .DIN2(n723), .Q(n1617) );
  nnd2s3 U965 ( .DIN1(n650), .DIN2(n857), .Q(n1616) );
  nnd2s3 U966 ( .DIN1(n1618), .DIN2(n1619), .Q(g6804) );
  nnd2s3 U967 ( .DIN1(n1601), .DIN2(n556), .Q(n1619) );
  nnd2s3 U968 ( .DIN1(n650), .DIN2(n705), .Q(n1618) );
  nnd2s3 U969 ( .DIN1(n1620), .DIN2(n1621), .Q(g6803) );
  nnd2s3 U970 ( .DIN1(n1601), .DIN2(n727), .Q(n1621) );
  nnd2s3 U971 ( .DIN1(n650), .DIN2(n642), .Q(n1620) );
  nor2s3 U972 ( .DIN1(n1427), .DIN2(n1622), .Q(g6802) );
  nor2s3 U973 ( .DIN1(n1623), .DIN2(n1624), .Q(n1622) );
  nor2s3 U974 ( .DIN1(n1990), .DIN2(g6800), .Q(n1624) );
  nor2s3 U975 ( .DIN1(n1999), .DIN2(n1229), .Q(n1623) );
  nor2s3 U976 ( .DIN1(n1212), .DIN2(n1999), .Q(n1427) );
  nnd2s3 U977 ( .DIN1(n695), .DIN2(n1625), .Q(g6801) );
  nnd2s3 U978 ( .DIN1(n1626), .DIN2(n1212), .Q(n1625) );
  or2s3 U979 ( .DIN1(n2573), .DIN2(n1990), .Q(n1212) );
  nnd2s3 U980 ( .DIN1(n2573), .DIN2(n1990), .Q(n1626) );
  or2s3 U981 ( .DIN1(n1229), .DIN2(n2573), .Q(g6800) );
  nnd3s3 U982 ( .DIN1(n696), .DIN2(g745), .DIN3(g109), .Q(n1229) );
  and3s3 U983 ( .DIN1(n1627), .DIN2(n1430), .DIN3(n841), .Q(g6799) );
  or3s3 U984 ( .DIN1(n2058), .DIN2(n2574), .DIN3(n2051), .Q(n1430) );
  nnd2s3 U985 ( .DIN1(n2058), .DIN2(n1628), .Q(n1627) );
  nnd2s3 U986 ( .DIN1(n625), .DIN2(n808), .Q(n1628) );
  nnd2s3 U987 ( .DIN1(n1629), .DIN2(n1630), .Q(g6798) );
  nnd3s3 U988 ( .DIN1(n841), .DIN2(n808), .DIN3(n2051), .Q(n1630) );
  nnd2s3 U989 ( .DIN1(g6797), .DIN2(n625), .Q(n1629) );
  nor2s3 U990 ( .DIN1(n808), .DIN2(n1280), .Q(g6797) );
  nnd2s3 U991 ( .DIN1(n2575), .DIN2(g109), .Q(n1280) );
  or4s3 U993 ( .DIN1(n676), .DIN2(n1397), .DIN3(n1952), .DIN4(n2025), .Q(n1631) );
  nnd3s3 U994 ( .DIN1(n722), .DIN2(n813), .DIN3(n532), .Q(n1397) );
  nnd2s3 U995 ( .DIN1(n1632), .DIN2(n1633), .Q(g6337) );
  or2s3 U996 ( .DIN1(n2849), .DIN2(n1979), .Q(n1633) );
  nnd2s3 U997 ( .DIN1(n2848), .DIN2(n778), .Q(n1632) );
  nnd2s3 U998 ( .DIN1(n1634), .DIN2(n1635), .Q(g6336) );
  nnd2s3 U999 ( .DIN1(n2853), .DIN2(n778), .Q(n1635) );
  nnd2s3 U1000 ( .DIN1(n2848), .DIN2(g1710), .Q(n1634) );
  nor2s3 U1001 ( .DIN1(n2724), .DIN2(n2848), .Q(g6330) );
  and2s3 U1002 ( .DIN1(g109), .DIN2(n2585), .Q(g6313) );
  nor2s3 U1003 ( .DIN1(n1970), .DIN2(n2866), .Q(g6312) );
  nor2s3 U1004 ( .DIN1(n1944), .DIN2(n2866), .Q(g6311) );
  nor2s3 U1005 ( .DIN1(n2013), .DIN2(n2866), .Q(g6310) );
  nor2s3 U1006 ( .DIN1(n1971), .DIN2(n2866), .Q(g6309) );
  nor2s3 U1007 ( .DIN1(n1945), .DIN2(n2866), .Q(g6308) );
  nor2s3 U1008 ( .DIN1(n2014), .DIN2(n2866), .Q(g6307) );
  nor2s3 U1009 ( .DIN1(n2015), .DIN2(n2866), .Q(g6306) );
  nor2s3 U1010 ( .DIN1(n2016), .DIN2(n2866), .Q(g6305) );
  nor2s3 U1011 ( .DIN1(n1988), .DIN2(n2865), .Q(g6304) );
  nor2s3 U1012 ( .DIN1(n2870), .DIN2(n739), .Q(g6303) );
  nor2s3 U1013 ( .DIN1(n2871), .DIN2(n528), .Q(g6302) );
  nor2s3 U1014 ( .DIN1(n2871), .DIN2(n744), .Q(g6301) );
  nor2s3 U1015 ( .DIN1(n2871), .DIN2(n602), .Q(g6300) );
  nor2s3 U1016 ( .DIN1(n1969), .DIN2(n2865), .Q(g6299) );
  nor2s3 U1017 ( .DIN1(g4906), .DIN2(\DFF_489/net776 ), .Q(g5673) );
  nor2s3 U1018 ( .DIN1(g4906), .DIN2(\DFF_330/net617 ), .Q(g5671) );
  nor2s3 U1019 ( .DIN1(g4906), .DIN2(\DFF_385/net672 ), .Q(g5670) );
  nnd2s3 U1020 ( .DIN1(n1636), .DIN2(n1637), .Q(g5669) );
  nnd2s3 U1021 ( .DIN1(n683), .DIN2(n670), .Q(n1637) );
  nnd2s3 U1022 ( .DIN1(n1638), .DIN2(n714), .Q(n1636) );
  nnd2s3 U1023 ( .DIN1(n1639), .DIN2(n1640), .Q(g5668) );
  nnd2s3 U1024 ( .DIN1(n683), .DIN2(n812), .Q(n1640) );
  nnd2s3 U1025 ( .DIN1(n1638), .DIN2(n825), .Q(n1639) );
  nnd2s3 U1026 ( .DIN1(n1641), .DIN2(n1642), .Q(g5667) );
  nnd2s3 U1027 ( .DIN1(n683), .DIN2(n682), .Q(n1642) );
  nnd2s3 U1028 ( .DIN1(n1638), .DIN2(n623), .Q(n1641) );
  nnd2s3 U1029 ( .DIN1(n1643), .DIN2(n1644), .Q(g5666) );
  nnd2s3 U1030 ( .DIN1(n683), .DIN2(n828), .Q(n1644) );
  or2s3 U1031 ( .DIN1(n683), .DIN2(n2751), .Q(n1643) );
  nnd2s3 U1032 ( .DIN1(n1645), .DIN2(n1646), .Q(g5665) );
  nnd2s3 U1033 ( .DIN1(n683), .DIN2(n836), .Q(n1646) );
  or2s3 U1034 ( .DIN1(n683), .DIN2(n2765), .Q(n1645) );
  nnd2s3 U1035 ( .DIN1(n1647), .DIN2(n1648), .Q(g5664) );
  nnd2s3 U1036 ( .DIN1(n683), .DIN2(n676), .Q(n1648) );
  or2s3 U1037 ( .DIN1(n683), .DIN2(n2777), .Q(n1647) );
  nnd2s3 U1038 ( .DIN1(n1649), .DIN2(n1650), .Q(g5663) );
  nnd2s3 U1039 ( .DIN1(n683), .DIN2(n532), .Q(n1650) );
  or2s3 U1040 ( .DIN1(n683), .DIN2(n2791), .Q(n1649) );
  nnd2s3 U1041 ( .DIN1(n1651), .DIN2(n1652), .Q(g5662) );
  nnd2s3 U1042 ( .DIN1(n683), .DIN2(n722), .Q(n1652) );
  or2s3 U1043 ( .DIN1(n683), .DIN2(n2801), .Q(n1651) );
  nnd2s3 U1044 ( .DIN1(n1653), .DIN2(n1654), .Q(g5661) );
  nnd2s3 U1045 ( .DIN1(n683), .DIN2(n813), .Q(n1654) );
  nnd2s3 U1046 ( .DIN1(n1638), .DIN2(n720), .Q(n1653) );
  nnd2s3 U1047 ( .DIN1(n2617), .DIN2(n2578), .Q(g5660) );
  and3s3 U1048 ( .DIN1(g743), .DIN2(g109), .DIN3(g744), .Q(g5659) );
  and3s3 U1049 ( .DIN1(g741), .DIN2(g109), .DIN3(g742), .Q(g5658) );
  nor2s3 U1050 ( .DIN1(g4894), .DIN2(\DFF_157/net444 ), .Q(g5657) );
  nor2s3 U1051 ( .DIN1(g4894), .DIN2(n806), .Q(g5656) );
  nor2s3 U1052 ( .DIN1(g4894), .DIN2(\DFF_136/net423 ), .Q(g5655) );
  nor2s3 U1053 ( .DIN1(g4894), .DIN2(\DFF_336/net623 ), .Q(g5654) );
  nor2s3 U1054 ( .DIN1(n826), .DIN2(n873), .Q(g4907) );
  nnd2s3 U1055 ( .DIN1(g1700), .DIN2(\DFF_275/net562 ), .Q(g4901) );
  nor4s3 U1056 ( .DIN1(n2007), .DIN2(n2045), .DIN3(n2046), .DIN4(n2047), .Q(
        g4897) );
  nnd2s3 U1057 ( .DIN1(n1655), .DIN2(n1656), .Q(g4895) );
  nnd2s3 U1058 ( .DIN1(n608), .DIN2(n696), .Q(n1656) );
  nnd2s3 U1059 ( .DIN1(g4171), .DIN2(n607), .Q(n1655) );
  nnd2s3 U1060 ( .DIN1(n948), .DIN2(n1657), .Q(g4894) );
  nnd2s3 U1061 ( .DIN1(n1951), .DIN2(n797), .Q(n1657) );
  nnd3s3 U1062 ( .DIN1(n1975), .DIN2(n1951), .DIN3(n1126), .Q(n948) );
  nor2s3 U1063 ( .DIN1(n691), .DIN2(n660), .Q(n1126) );
  nor2s3 U1064 ( .DIN1(g750), .DIN2(n2577), .Q(g4171) );
  nor2s3 U1065 ( .DIN1(n684), .DIN2(g1737), .Q(g3329) );
  nor2s3 U1066 ( .DIN1(n1658), .DIN2(n1659), .Q(g11657) );
  and2s3 U1067 ( .DIN1(n1660), .DIN2(n1661), .Q(n1658) );
  nnd3s3 U1068 ( .DIN1(n552), .DIN2(n765), .DIN3(n1662), .Q(n1661) );
  nnd2s3 U1069 ( .DIN1(n1663), .DIN2(n551), .Q(n1660) );
  nnd2s3 U1070 ( .DIN1(g4898), .DIN2(n545), .Q(n1663) );
  nor4s3 U1071 ( .DIN1(n2000), .DIN2(n2796), .DIN3(n2782), .DIN4(n2757), .Q(
        g4898) );
  nor2s3 U1072 ( .DIN1(n1659), .DIN2(n1664), .Q(g11656) );
  xor2s3 U1073 ( .DIN1(n2000), .DIN2(n1662), .Q(n1664) );
  nor2s3 U1074 ( .DIN1(n1665), .DIN2(n2782), .Q(n1662) );
  nor2s3 U1075 ( .DIN1(n1659), .DIN2(n1666), .Q(g11655) );
  xnr2s3 U1076 ( .DIN1(n2782), .DIN2(n1665), .Q(n1666) );
  and3s3 U1077 ( .DIN1(n1667), .DIN2(n1665), .DIN3(n673), .Q(g11654) );
  nnd2s3 U1078 ( .DIN1(g109), .DIN2(n1668), .Q(n1659) );
  nnd3s3 U1079 ( .DIN1(n1669), .DIN2(n701), .DIN3(n2011), .Q(n1668) );
  or2s3 U1080 ( .DIN1(n1670), .DIN2(n2796), .Q(n1665) );
  nnd2s3 U1081 ( .DIN1(n2796), .DIN2(n1670), .Q(n1667) );
  nnd2s3 U1082 ( .DIN1(n1671), .DIN2(n1672), .Q(g11653) );
  nnd2s3 U1083 ( .DIN1(n608), .DIN2(n1673), .Q(n1672) );
  nnd2s3 U1084 ( .DIN1(n1674), .DIN2(n1675), .Q(n1673) );
  nnd2s3 U1085 ( .DIN1(n1676), .DIN2(n1677), .Q(n1675) );
  or2s3 U1086 ( .DIN1(n1678), .DIN2(n1677), .Q(n1674) );
  nnd2s3 U1087 ( .DIN1(n1432), .DIN2(n727), .Q(n1671) );
  nnd2s3 U1088 ( .DIN1(n1679), .DIN2(n1680), .Q(g11642) );
  nnd2s3 U1089 ( .DIN1(n1681), .DIN2(n608), .Q(n1680) );
  xnr2s3 U1090 ( .DIN1(n1678), .DIN2(n1676), .Q(n1681) );
  xor2s3 U1091 ( .DIN1(n1682), .DIN2(n1683), .Q(n1676) );
  xor2s3 U1092 ( .DIN1(n1684), .DIN2(n1685), .Q(n1683) );
  xor2s3 U1093 ( .DIN1(n1686), .DIN2(n1687), .Q(n1685) );
  xor2s3 U1094 ( .DIN1(n1688), .DIN2(n1689), .Q(n1687) );
  xor2s3 U1095 ( .DIN1(n1690), .DIN2(n1691), .Q(n1686) );
  xor2s3 U1096 ( .DIN1(n1692), .DIN2(n1693), .Q(n1684) );
  xor2s3 U1097 ( .DIN1(n1694), .DIN2(n1695), .Q(n1693) );
  xor2s3 U1098 ( .DIN1(n1696), .DIN2(n1697), .Q(n1692) );
  nnd2s3 U1099 ( .DIN1(n1698), .DIN2(n1699), .Q(n1678) );
  nnd2s3 U1100 ( .DIN1(n1700), .DIN2(n2830), .Q(n1699) );
  xor2s3 U1101 ( .DIN1(n1702), .DIN2(n1703), .Q(n1700) );
  nor2s3 U1102 ( .DIN1(n1704), .DIN2(n731), .Q(n1703) );
  nnd2s3 U1103 ( .DIN1(n2834), .DIN2(n724), .Q(n1698) );
  nnd2s3 U1104 ( .DIN1(n1432), .DIN2(n723), .Q(n1679) );
  nnd2s3 U1105 ( .DIN1(n1705), .DIN2(n1706), .Q(g11635) );
  nnd2s3 U1106 ( .DIN1(n544), .DIN2(n670), .Q(n1706) );
  nnd2s3 U1107 ( .DIN1(n1707), .DIN2(n793), .Q(n1705) );
  nnd2s3 U1108 ( .DIN1(n1708), .DIN2(n1709), .Q(g11634) );
  nnd2s3 U1109 ( .DIN1(n544), .DIN2(n812), .Q(n1709) );
  nnd2s3 U1110 ( .DIN1(n1707), .DIN2(n606), .Q(n1708) );
  nnd2s3 U1111 ( .DIN1(n1710), .DIN2(n1711), .Q(g11633) );
  nnd2s3 U1112 ( .DIN1(n544), .DIN2(n682), .Q(n1711) );
  nnd2s3 U1113 ( .DIN1(n1707), .DIN2(n767), .Q(n1710) );
  nnd2s3 U1114 ( .DIN1(n1712), .DIN2(n1713), .Q(g11632) );
  nnd2s3 U1115 ( .DIN1(n544), .DIN2(n828), .Q(n1713) );
  nnd2s3 U1116 ( .DIN1(n1707), .DIN2(n681), .Q(n1712) );
  nnd2s3 U1117 ( .DIN1(n1714), .DIN2(n1715), .Q(g11631) );
  nnd2s3 U1118 ( .DIN1(n544), .DIN2(n836), .Q(n1715) );
  nnd2s3 U1119 ( .DIN1(n1707), .DIN2(n584), .Q(n1714) );
  nnd2s3 U1120 ( .DIN1(n1716), .DIN2(n1717), .Q(g11630) );
  nnd2s3 U1121 ( .DIN1(n544), .DIN2(n676), .Q(n1717) );
  nnd2s3 U1122 ( .DIN1(n1707), .DIN2(n597), .Q(n1716) );
  nnd2s3 U1123 ( .DIN1(n1718), .DIN2(n1719), .Q(g11629) );
  nnd2s3 U1124 ( .DIN1(n544), .DIN2(n532), .Q(n1719) );
  or2s3 U1125 ( .DIN1(n544), .DIN2(n2786), .Q(n1718) );
  nnd2s3 U1126 ( .DIN1(n1720), .DIN2(n1721), .Q(g11628) );
  nnd2s3 U1127 ( .DIN1(n544), .DIN2(n722), .Q(n1721) );
  or2s3 U1128 ( .DIN1(n544), .DIN2(n2800), .Q(n1720) );
  nnd2s3 U1129 ( .DIN1(n1722), .DIN2(n1723), .Q(g11627) );
  nnd2s3 U1130 ( .DIN1(n544), .DIN2(n813), .Q(n1723) );
  nnd2s3 U1131 ( .DIN1(n1707), .DIN2(n798), .Q(n1722) );
  nnd2s3 U1132 ( .DIN1(n545), .DIN2(g1317), .Q(n1707) );
  or3s3 U1133 ( .DIN1(n1724), .DIN2(n1340), .DIN3(n1725), .Q(n1670) );
  nor6s3 U1134 ( .DIN1(n1726), .DIN2(n1727), .DIN3(n1728), .DIN4(n1729), 
        .DIN5(n1730), .DIN6(n1731), .Q(n1724) );
  xnr2s3 U1135 ( .DIN1(n1732), .DIN2(n1733), .Q(n1731) );
  xor2s3 U1136 ( .DIN1(n2605), .DIN2(n2654), .Q(n1730) );
  xor2s3 U1137 ( .DIN1(n2612), .DIN2(n2655), .Q(n1729) );
  xor2s3 U1138 ( .DIN1(n2611), .DIN2(n2648), .Q(n1728) );
  xor2s3 U1139 ( .DIN1(n2615), .DIN2(n2647), .Q(n1727) );
  or5s3 U1140 ( .DIN1(n1734), .DIN2(n1735), .DIN3(n1736), .DIN4(n1737), .DIN5(
        n1738), .Q(n1726) );
  xor2s3 U1141 ( .DIN1(n2604), .DIN2(n2652), .Q(n1738) );
  xor2s3 U1142 ( .DIN1(n2614), .DIN2(n2651), .Q(n1737) );
  xor2s3 U1143 ( .DIN1(n2616), .DIN2(n2650), .Q(n1736) );
  xor2s3 U1144 ( .DIN1(n2606), .DIN2(n2653), .Q(n1735) );
  xor2s3 U1145 ( .DIN1(n2613), .DIN2(n2649), .Q(n1734) );
  nnd2s3 U1146 ( .DIN1(n1739), .DIN2(n1740), .Q(g11611) );
  nnd2s3 U1147 ( .DIN1(n2848), .DIN2(n1741), .Q(n1740) );
  xor2s3 U1148 ( .DIN1(n1742), .DIN2(n1743), .Q(n1741) );
  xor2s3 U1149 ( .DIN1(n684), .DIN2(n1744), .Q(n1743) );
  nnd2s3 U1150 ( .DIN1(n1745), .DIN2(n1746), .Q(n1742) );
  nnd4s2 U1151 ( .DIN1(n1976), .DIN2(n1148), .DIN3(n1949), .DIN4(n1747), .Q(
        n1746) );
  nnd2s3 U1152 ( .DIN1(n527), .DIN2(n1748), .Q(n1745) );
  nnd3s3 U1153 ( .DIN1(n1148), .DIN2(n1949), .DIN3(n1976), .Q(n1748) );
  nor2s3 U1154 ( .DIN1(n620), .DIN2(n1974), .Q(n1148) );
  nnd2s3 U1155 ( .DIN1(n1749), .DIN2(n1750), .Q(n1747) );
  nnd2s3 U1156 ( .DIN1(n2016), .DIN2(n1751), .Q(n1750) );
  nnd2s3 U1157 ( .DIN1(n1988), .DIN2(n1752), .Q(n1751) );
  or5s3 U1158 ( .DIN1(n2585), .DIN2(n585), .DIN3(n632), .DIN4(n1753), .DIN5(
        n1754), .Q(n1752) );
  nnd4s2 U1159 ( .DIN1(n1970), .DIN2(n1944), .DIN3(n1969), .DIN4(n1755), .Q(
        n1754) );
  and3s3 U1160 ( .DIN1(n1971), .DIN2(n1945), .DIN3(n2013), .Q(n1755) );
  nnd4s2 U1161 ( .DIN1(n739), .DIN2(n528), .DIN3(n744), .DIN4(n602), .Q(n1753)
         );
  nnd2s3 U1162 ( .DIN1(n1988), .DIN2(n637), .Q(n1749) );
  nnd2s3 U1163 ( .DIN1(n2853), .DIN2(n549), .Q(n1739) );
  nor2s3 U1164 ( .DIN1(n2871), .DIN2(n1756), .Q(g11594) );
  xor2s3 U1165 ( .DIN1(n1757), .DIN2(n1758), .Q(n1756) );
  xor2s3 U1166 ( .DIN1(n2589), .DIN2(n1744), .Q(n1758) );
  and2s3 U1167 ( .DIN1(n1759), .DIN2(n1760), .Q(n1744) );
  nnd2s3 U1168 ( .DIN1(n2862), .DIN2(n1761), .Q(n1760) );
  nnd2s3 U1169 ( .DIN1(n1762), .DIN2(n1763), .Q(n1761) );
  nnd2s3 U1170 ( .DIN1(n1764), .DIN2(n1765), .Q(n1763) );
  nnd4s2 U1171 ( .DIN1(n550), .DIN2(n860), .DIN3(n615), .DIN4(n576), .Q(n1765)
         );
  nnd2s3 U1172 ( .DIN1(n1766), .DIN2(n571), .Q(n1764) );
  or5s3 U1173 ( .DIN1(n2643), .DIN2(n2644), .DIN3(n2645), .DIN4(n2646), .DIN5(
        n616), .Q(n1762) );
  or2s3 U1174 ( .DIN1(n2863), .DIN2(n1995), .Q(n1759) );
  xor2s3 U1175 ( .DIN1(n2588), .DIN2(n1767), .Q(n1757) );
  xor2s3 U1176 ( .DIN1(n2586), .DIN2(n2587), .Q(n1767) );
  nnd2s3 U1177 ( .DIN1(n1768), .DIN2(n1769), .Q(g11513) );
  nnd2s3 U1178 ( .DIN1(n608), .DIN2(n1695), .Q(n1769) );
  nnd2s3 U1179 ( .DIN1(n1770), .DIN2(n1771), .Q(n1695) );
  nnd2s3 U1180 ( .DIN1(n1772), .DIN2(n2831), .Q(n1771) );
  xor2s3 U1181 ( .DIN1(n1773), .DIN2(n2630), .Q(n1772) );
  nnd4s2 U1182 ( .DIN1(n1977), .DIN2(n1930), .DIN3(n789), .DIN4(n726), .Q(
        n1773) );
  or2s3 U1183 ( .DIN1(n2831), .DIN2(n2667), .Q(n1770) );
  nnd2s3 U1184 ( .DIN1(n1432), .DIN2(n746), .Q(n1768) );
  nnd2s3 U1185 ( .DIN1(n1774), .DIN2(n1775), .Q(g11512) );
  nnd2s3 U1186 ( .DIN1(n608), .DIN2(n1689), .Q(n1775) );
  nnd2s3 U1187 ( .DIN1(n1776), .DIN2(n1777), .Q(n1689) );
  nnd2s3 U1188 ( .DIN1(n1778), .DIN2(n2831), .Q(n1777) );
  xor2s3 U1189 ( .DIN1(n525), .DIN2(n1779), .Q(n1778) );
  nor2s3 U1190 ( .DIN1(n865), .DIN2(n1780), .Q(n1779) );
  or2s3 U1191 ( .DIN1(n2831), .DIN2(n2688), .Q(n1776) );
  nnd2s3 U1192 ( .DIN1(n1432), .DIN2(n693), .Q(n1774) );
  nnd2s3 U1193 ( .DIN1(n1781), .DIN2(n1782), .Q(g11511) );
  nnd2s3 U1194 ( .DIN1(n608), .DIN2(n1688), .Q(n1782) );
  nnd2s3 U1195 ( .DIN1(n1783), .DIN2(n1784), .Q(n1688) );
  nnd2s3 U1196 ( .DIN1(n1785), .DIN2(n2831), .Q(n1784) );
  xor2s3 U1197 ( .DIN1(n1786), .DIN2(n2629), .Q(n1785) );
  nnd2s3 U1198 ( .DIN1(n725), .DIN2(n1950), .Q(n1786) );
  or2s3 U1199 ( .DIN1(n2831), .DIN2(n2690), .Q(n1783) );
  nnd2s3 U1200 ( .DIN1(n1432), .DIN2(n740), .Q(n1781) );
  nnd2s3 U1201 ( .DIN1(n1787), .DIN2(n1788), .Q(g11510) );
  nnd2s3 U1202 ( .DIN1(n608), .DIN2(n1694), .Q(n1788) );
  nnd2s3 U1203 ( .DIN1(n1789), .DIN2(n1790), .Q(n1694) );
  nnd2s3 U1204 ( .DIN1(n1791), .DIN2(n2830), .Q(n1790) );
  xor2s3 U1205 ( .DIN1(n748), .DIN2(n1792), .Q(n1791) );
  nor2s3 U1206 ( .DIN1(n1930), .DIN2(n1793), .Q(n1792) );
  or2s3 U1207 ( .DIN1(n2831), .DIN2(n2684), .Q(n1789) );
  nnd2s3 U1208 ( .DIN1(n1432), .DIN2(n713), .Q(n1787) );
  nnd2s3 U1209 ( .DIN1(n1794), .DIN2(n1795), .Q(g11509) );
  nnd2s3 U1210 ( .DIN1(n608), .DIN2(n1682), .Q(n1795) );
  nnd2s3 U1211 ( .DIN1(n1796), .DIN2(n1797), .Q(n1682) );
  nnd2s3 U1212 ( .DIN1(n1798), .DIN2(n2830), .Q(n1797) );
  xor2s3 U1213 ( .DIN1(n843), .DIN2(n1799), .Q(n1798) );
  nor2s3 U1214 ( .DIN1(n1977), .DIN2(n1704), .Q(n1799) );
  nnd3s3 U1215 ( .DIN1(n1930), .DIN2(n726), .DIN3(n1950), .Q(n1704) );
  or2s3 U1216 ( .DIN1(n2831), .DIN2(n2682), .Q(n1796) );
  nnd2s3 U1217 ( .DIN1(n1432), .DIN2(n751), .Q(n1794) );
  nnd2s3 U1218 ( .DIN1(n1800), .DIN2(n1801), .Q(g11508) );
  nnd2s3 U1219 ( .DIN1(n608), .DIN2(n1697), .Q(n1801) );
  nnd2s3 U1220 ( .DIN1(n1802), .DIN2(n1803), .Q(n1697) );
  nnd2s3 U1221 ( .DIN1(n1804), .DIN2(n2830), .Q(n1803) );
  xor2s3 U1222 ( .DIN1(n678), .DIN2(n1805), .Q(n1804) );
  nor2s3 U1223 ( .DIN1(n865), .DIN2(n1793), .Q(n1805) );
  nnd3s3 U1224 ( .DIN1(n1950), .DIN2(n731), .DIN3(n2073), .Q(n1793) );
  or2s3 U1225 ( .DIN1(n2831), .DIN2(n2686), .Q(n1802) );
  nnd2s3 U1226 ( .DIN1(n1432), .DIN2(n831), .Q(n1800) );
  nnd2s3 U1227 ( .DIN1(n1806), .DIN2(n1807), .Q(g11507) );
  nnd2s3 U1228 ( .DIN1(n608), .DIN2(n1691), .Q(n1807) );
  nnd2s3 U1229 ( .DIN1(n1808), .DIN2(n1809), .Q(n1691) );
  nnd2s3 U1230 ( .DIN1(n1810), .DIN2(n2830), .Q(n1809) );
  xor2s3 U1231 ( .DIN1(n790), .DIN2(n1811), .Q(n1810) );
  nor2s3 U1232 ( .DIN1(n2073), .DIN2(n1812), .Q(n1811) );
  or2s3 U1233 ( .DIN1(n2831), .DIN2(n2665), .Q(n1808) );
  nnd2s3 U1234 ( .DIN1(n1432), .DIN2(n824), .Q(n1806) );
  nnd2s3 U1235 ( .DIN1(n1813), .DIN2(n1814), .Q(g11506) );
  nnd2s3 U1236 ( .DIN1(n608), .DIN2(n1690), .Q(n1814) );
  nnd2s3 U1237 ( .DIN1(n1815), .DIN2(n1816), .Q(n1690) );
  nnd2s3 U1238 ( .DIN1(n1817), .DIN2(n2830), .Q(n1816) );
  xor2s3 U1239 ( .DIN1(n609), .DIN2(n1818), .Q(n1817) );
  nor2s3 U1240 ( .DIN1(n726), .DIN2(n1812), .Q(n1818) );
  nnd3s3 U1241 ( .DIN1(n1950), .DIN2(n865), .DIN3(n1977), .Q(n1812) );
  or2s3 U1242 ( .DIN1(n2831), .DIN2(n2666), .Q(n1815) );
  nnd2s3 U1243 ( .DIN1(n1432), .DIN2(n601), .Q(n1813) );
  nnd2s3 U1244 ( .DIN1(n1819), .DIN2(n1820), .Q(g11505) );
  nnd2s3 U1245 ( .DIN1(n1432), .DIN2(n556), .Q(n1820) );
  nnd2s3 U1246 ( .DIN1(n608), .DIN2(n1696), .Q(n1819) );
  nnd2s3 U1247 ( .DIN1(n1821), .DIN2(n1822), .Q(n1696) );
  nnd2s3 U1248 ( .DIN1(n1823), .DIN2(n2830), .Q(n1822) );
  xor2s3 U1249 ( .DIN1(n640), .DIN2(n1824), .Q(n1823) );
  nor2s3 U1250 ( .DIN1(n1930), .DIN2(n1780), .Q(n1824) );
  nnd3s3 U1251 ( .DIN1(n1977), .DIN2(n789), .DIN3(n2073), .Q(n1780) );
  or2s3 U1252 ( .DIN1(n2831), .DIN2(n2668), .Q(n1821) );
  nnd2s3 U1253 ( .DIN1(n2599), .DIN2(g750), .Q(n1432) );
  nor2s3 U1254 ( .DIN1(n1825), .DIN2(n1826), .Q(g11473) );
  and2s3 U1255 ( .DIN1(n1827), .DIN2(n1828), .Q(n1825) );
  nnd3s3 U1256 ( .DIN1(n703), .DIN2(n842), .DIN3(n1829), .Q(n1828) );
  nnd2s3 U1257 ( .DIN1(n1830), .DIN2(n704), .Q(n1827) );
  nnd2s3 U1258 ( .DIN1(n2827), .DIN2(n518), .Q(n1830) );
  nor4s3 U1259 ( .DIN1(n2044), .DIN2(n2787), .DIN3(n2760), .DIN4(n2748), .Q(
        n2827) );
  nor2s3 U1260 ( .DIN1(n1826), .DIN2(n1831), .Q(g11472) );
  xor2s3 U1261 ( .DIN1(n2760), .DIN2(n1829), .Q(n1831) );
  nor2s3 U1262 ( .DIN1(n1832), .DIN2(n2044), .Q(n1829) );
  nor2s3 U1263 ( .DIN1(n1826), .DIN2(n1833), .Q(g11471) );
  xnr2s3 U1264 ( .DIN1(n2044), .DIN2(n1832), .Q(n1833) );
  and3s3 U1265 ( .DIN1(n1834), .DIN2(n1832), .DIN3(n768), .Q(g11470) );
  nnd2s3 U1266 ( .DIN1(g109), .DIN2(n1835), .Q(n1826) );
  nnd3s3 U1267 ( .DIN1(n1836), .DIN2(n769), .DIN3(n1837), .Q(n1835) );
  or2s3 U1268 ( .DIN1(n1838), .DIN2(n2787), .Q(n1832) );
  nnd2s3 U1269 ( .DIN1(n2787), .DIN2(n1838), .Q(n1834) );
  nor2s3 U1270 ( .DIN1(n1839), .DIN2(n1840), .Q(g11469) );
  nor2s3 U1271 ( .DIN1(n1841), .DIN2(n789), .Q(n1839) );
  nor2s3 U1272 ( .DIN1(n1842), .DIN2(n1840), .Q(g11468) );
  and2s3 U1273 ( .DIN1(n1843), .DIN2(n1844), .Q(n1842) );
  nnd3s3 U1274 ( .DIN1(n1845), .DIN2(n865), .DIN3(n1846), .Q(n1844) );
  or2s3 U1275 ( .DIN1(n1841), .DIN2(n1977), .Q(n1843) );
  nor2s3 U1276 ( .DIN1(n1847), .DIN2(n1845), .Q(n1841) );
  nor2s3 U1277 ( .DIN1(n1840), .DIN2(n1848), .Q(g11467) );
  xor2s3 U1278 ( .DIN1(n865), .DIN2(n521), .Q(n1848) );
  and3s3 U1279 ( .DIN1(n1849), .DIN2(n521), .DIN3(n600), .Q(g11466) );
  nnd2s3 U1280 ( .DIN1(g109), .DIN2(\DFF_441/net728 ), .Q(n1840) );
  nor2s3 U1281 ( .DIN1(n1847), .DIN2(n2073), .Q(n1846) );
  nnd2s3 U1282 ( .DIN1(n2073), .DIN2(n1847), .Q(n1849) );
  nnd2s3 U1283 ( .DIN1(n2828), .DIN2(n1850), .Q(n1847) );
  nnd2s3 U1284 ( .DIN1(n725), .DIN2(n789), .Q(n1850) );
  nnd3s3 U1285 ( .DIN1(n731), .DIN2(n726), .DIN3(n865), .Q(n1845) );
  nnd2s3 U1286 ( .DIN1(n1851), .DIN2(n1852), .Q(g11443) );
  nnd2s3 U1287 ( .DIN1(n1564), .DIN2(n570), .Q(n1852) );
  nor2s3 U1288 ( .DIN1(n2871), .DIN2(n649), .Q(n1564) );
  nnd2s3 U1289 ( .DIN1(n649), .DIN2(n1732), .Q(n1851) );
  nnd2s3 U1290 ( .DIN1(n1853), .DIN2(n1854), .Q(n1732) );
  nnd2s3 U1291 ( .DIN1(n618), .DIN2(n1855), .Q(n1854) );
  nnd2s3 U1292 ( .DIN1(n1856), .DIN2(n1857), .Q(n1855) );
  nnd2s3 U1293 ( .DIN1(n2052), .DIN2(n1858), .Q(n1857) );
  nnd2s3 U1294 ( .DIN1(n2031), .DIN2(n1859), .Q(n1858) );
  or5s3 U1295 ( .DIN1(n734), .DIN2(n834), .DIN3(n557), .DIN4(n1860), .DIN5(
        n1861), .Q(n1859) );
  nnd4s2 U1296 ( .DIN1(n2612), .DIN2(n2613), .DIN3(n2611), .DIN4(n1862), .Q(
        n1861) );
  and4s2 U1297 ( .DIN1(n2614), .DIN2(n2615), .DIN3(n2616), .DIN4(n2605), .Q(
        n1862) );
  nnd3s3 U1298 ( .DIN1(n2606), .DIN2(n2607), .DIN3(n2604), .Q(n1860) );
  nnd2s3 U1299 ( .DIN1(n2031), .DIN2(n631), .Q(n1856) );
  or2s3 U1300 ( .DIN1(n1733), .DIN2(n618), .Q(n1853) );
  nnd3s3 U1301 ( .DIN1(n856), .DIN2(n619), .DIN3(n1335), .Q(n1340) );
  nor2s3 U1302 ( .DIN1(n2601), .DIN2(n2602), .Q(n1335) );
  xnr2s3 U1303 ( .DIN1(n1863), .DIN2(n2816), .Q(n1733) );
  nnd2s3 U1304 ( .DIN1(n743), .DIN2(n1677), .Q(n1863) );
  or3s3 U1305 ( .DIN1(n778), .DIN2(n2617), .DIN3(n2857), .Q(n1725) );
  nor2s3 U1306 ( .DIN1(n1864), .DIN2(n1865), .Q(g11442) );
  nor2s3 U1307 ( .DIN1(n1866), .DIN2(n567), .Q(n1864) );
  nor2s3 U1308 ( .DIN1(n1867), .DIN2(n1868), .Q(n1866) );
  nor2s3 U1309 ( .DIN1(n1869), .DIN2(n1865), .Q(g11441) );
  and2s3 U1310 ( .DIN1(n1870), .DIN2(n1871), .Q(n1869) );
  nnd3s3 U1311 ( .DIN1(n1867), .DIN2(n757), .DIN3(n1872), .Q(n1871) );
  nnd2s3 U1312 ( .DIN1(n1873), .DIN2(n624), .Q(n1870) );
  or2s3 U1313 ( .DIN1(n1868), .DIN2(n1867), .Q(n1873) );
  nor2s3 U1314 ( .DIN1(n1865), .DIN2(n1874), .Q(g11440) );
  xor2s3 U1315 ( .DIN1(n757), .DIN2(n520), .Q(n1874) );
  and3s3 U1316 ( .DIN1(n1875), .DIN2(n520), .DIN3(n770), .Q(g11439) );
  nnd2s3 U1317 ( .DIN1(n2618), .DIN2(g109), .Q(n1865) );
  nor2s3 U1318 ( .DIN1(n1868), .DIN2(n2672), .Q(n1872) );
  nnd2s3 U1319 ( .DIN1(n2672), .DIN2(n1868), .Q(n1875) );
  nnd2s3 U1320 ( .DIN1(n568), .DIN2(n2830), .Q(n1868) );
  nnd3s3 U1321 ( .DIN1(n1876), .DIN2(n1877), .DIN3(n1878), .Q(g11409) );
  nnd2s3 U1322 ( .DIN1(n1384), .DIN2(n776), .Q(n1878) );
  nor2s3 U1323 ( .DIN1(n591), .DIN2(n920), .Q(n1384) );
  nnd3s3 U1324 ( .DIN1(n1879), .DIN2(n1880), .DIN3(n591), .Q(n1877) );
  nnd3s3 U1325 ( .DIN1(n1881), .DIN2(n718), .DIN3(n1882), .Q(n1880) );
  nnd2s3 U1326 ( .DIN1(n1883), .DIN2(n1884), .Q(n1882) );
  nnd2s3 U1327 ( .DIN1(n2825), .DIN2(n2822), .Q(n1884) );
  nnd2s3 U1328 ( .DIN1(g10774), .DIN2(n2824), .Q(n1883) );
  nnd2s3 U1329 ( .DIN1(n1885), .DIN2(n1886), .Q(n1881) );
  nnd2s3 U1330 ( .DIN1(n2823), .DIN2(n2820), .Q(n1886) );
  nnd2s3 U1331 ( .DIN1(n2818), .DIN2(n2821), .Q(n1885) );
  nnd2s3 U1333 ( .DIN1(n1889), .DIN2(n1890), .Q(n1888) );
  nnd2s3 U1334 ( .DIN1(n682), .DIN2(n812), .Q(n1890) );
  nnd2s3 U1335 ( .DIN1(n828), .DIN2(n836), .Q(n1889) );
  nnd2s3 U1336 ( .DIN1(n1891), .DIN2(n1892), .Q(n1887) );
  nnd2s3 U1337 ( .DIN1(n676), .DIN2(n532), .Q(n1892) );
  nnd2s3 U1338 ( .DIN1(n722), .DIN2(n813), .Q(n1891) );
  nnd3s3 U1339 ( .DIN1(n920), .DIN2(n1893), .DIN3(n1989), .Q(n1876) );
  nnd2s3 U1340 ( .DIN1(n935), .DIN2(n1980), .Q(n1893) );
  and2s3 U1341 ( .DIN1(n1894), .DIN2(n1895), .Q(n935) );
  nnd2s3 U1342 ( .DIN1(n1980), .DIN2(n698), .Q(n1895) );
  nor2s3 U1343 ( .DIN1(n809), .DIN2(n1386), .Q(n920) );
  nnd2s3 U1344 ( .DIN1(n1389), .DIN2(n862), .Q(n1386) );
  and2s3 U1345 ( .DIN1(n2626), .DIN2(n2627), .Q(n1389) );
  nnd2s3 U1346 ( .DIN1(n1896), .DIN2(n1897), .Q(g11408) );
  nnd2s3 U1347 ( .DIN1(n591), .DIN2(n1898), .Q(n1897) );
  nnd2s3 U1348 ( .DIN1(n1899), .DIN2(n1900), .Q(n1898) );
  nnd2s3 U1349 ( .DIN1(n535), .DIN2(n718), .Q(n1900) );
  nnd2s3 U1351 ( .DIN1(n1901), .DIN2(n927), .Q(n1896) );
  nnd2s3 U1352 ( .DIN1(n1894), .DIN2(n1902), .Q(n1901) );
  nnd2s3 U1353 ( .DIN1(n1903), .DIN2(g2731), .Q(n1902) );
  nnd3s3 U1354 ( .DIN1(n1904), .DIN2(n1905), .DIN3(g5672), .Q(n1903) );
  nor2s3 U1355 ( .DIN1(g4906), .DIN2(n733), .Q(g5672) );
  nnd2s3 U1356 ( .DIN1(n927), .DIN2(n1906), .Q(g4906) );
  nnd2s3 U1357 ( .DIN1(n1986), .DIN2(n589), .Q(n1906) );
  nnd3s3 U1358 ( .DIN1(n1986), .DIN2(n1948), .DIN3(n1043), .Q(n927) );
  nnd3s3 U1359 ( .DIN1(n1948), .DIN2(n747), .DIN3(n1043), .Q(n1905) );
  nor2s3 U1360 ( .DIN1(n652), .DIN2(n698), .Q(n1043) );
  xor2s3 U1361 ( .DIN1(n1907), .DIN2(n1908), .Q(n1904) );
  nnd2s3 U1362 ( .DIN1(n1909), .DIN2(n1910), .Q(n1908) );
  nnd2s3 U1363 ( .DIN1(n1989), .DIN2(n1911), .Q(n1910) );
  nnd2s3 U1364 ( .DIN1(n1948), .DIN2(n1912), .Q(n1911) );
  nnd2s3 U1365 ( .DIN1(n652), .DIN2(n702), .Q(n1912) );
  nnd2s3 U1366 ( .DIN1(n931), .DIN2(n776), .Q(n1909) );
  nor2s3 U1367 ( .DIN1(n702), .DIN2(n1953), .Q(n931) );
  or2s3 U1368 ( .DIN1(n936), .DIN2(n702), .Q(n1894) );
  nnd2s3 U1369 ( .DIN1(n1953), .DIN2(n652), .Q(n936) );
  nnd2s3 U1370 ( .DIN1(n1913), .DIN2(n1914), .Q(g11406) );
  nnd2s3 U1371 ( .DIN1(n517), .DIN2(n736), .Q(n1914) );
  nnd2s3 U1372 ( .DIN1(n1915), .DIN2(n667), .Q(n1913) );
  nnd2s3 U1373 ( .DIN1(n1916), .DIN2(n1917), .Q(g11405) );
  nnd2s3 U1374 ( .DIN1(n517), .DIN2(n654), .Q(n1917) );
  nnd2s3 U1375 ( .DIN1(n1915), .DIN2(n773), .Q(n1916) );
  nnd2s3 U1376 ( .DIN1(n1918), .DIN2(n1919), .Q(g11404) );
  nnd2s3 U1377 ( .DIN1(n517), .DIN2(n627), .Q(n1919) );
  nnd2s3 U1378 ( .DIN1(n1915), .DIN2(n791), .Q(n1918) );
  nnd2s3 U1379 ( .DIN1(n1920), .DIN2(n1921), .Q(g11403) );
  nnd2s3 U1380 ( .DIN1(n517), .DIN2(n671), .Q(n1921) );
  or2s3 U1381 ( .DIN1(n517), .DIN2(n2749), .Q(n1920) );
  nnd2s3 U1382 ( .DIN1(n1922), .DIN2(n1923), .Q(g11402) );
  nnd2s3 U1383 ( .DIN1(n517), .DIN2(n605), .Q(n1923) );
  or2s3 U1384 ( .DIN1(n517), .DIN2(n2761), .Q(n1922) );
  nnd2s3 U1385 ( .DIN1(n1924), .DIN2(n1927), .Q(g11401) );
  nnd2s3 U1386 ( .DIN1(n517), .DIN2(n622), .Q(n1927) );
  or2s3 U1387 ( .DIN1(n517), .DIN2(n2774), .Q(n1924) );
  nnd2s3 U1388 ( .DIN1(n1928), .DIN2(n1931), .Q(g11400) );
  nnd2s3 U1389 ( .DIN1(n517), .DIN2(n692), .Q(n1931) );
  or2s3 U1390 ( .DIN1(n517), .DIN2(n2788), .Q(n1928) );
  nnd2s3 U1391 ( .DIN1(n1934), .DIN2(n1940), .Q(g11399) );
  or2s3 U1392 ( .DIN1(n1915), .DIN2(n2664), .Q(n1940) );
  or2s3 U1393 ( .DIN1(n517), .DIN2(n2803), .Q(n1934) );
  nnd2s3 U1394 ( .DIN1(n1941), .DIN2(n1942), .Q(g11398) );
  nnd2s3 U1395 ( .DIN1(n517), .DIN2(n840), .Q(n1942) );
  nnd2s3 U1396 ( .DIN1(n1915), .DIN2(n690), .Q(n1941) );
  nnd3s3 U1397 ( .DIN1(n1943), .DIN2(n1836), .DIN3(n518), .Q(n1915) );
  or3s3 U1398 ( .DIN1(n2839), .DIN2(n1964), .DIN3(n568), .Q(n1838) );
  nor6s3 U1399 ( .DIN1(n1965), .DIN2(n1966), .DIN3(n1967), .DIN4(n1973), 
        .DIN5(n1997), .DIN6(n1998), .Q(n1964) );
  xor2s3 U1400 ( .DIN1(n724), .DIN2(n2003), .Q(n1998) );
  xor2s3 U1401 ( .DIN1(n2667), .DIN2(n2674), .Q(n1997) );
  xor2s3 U1402 ( .DIN1(n2668), .DIN2(n2676), .Q(n1973) );
  xor2s3 U1403 ( .DIN1(n2665), .DIN2(n2681), .Q(n1967) );
  xor2s3 U1404 ( .DIN1(n2666), .DIN2(n2675), .Q(n1966) );
  or5s3 U1405 ( .DIN1(n2004), .DIN2(n2005), .DIN3(n2006), .DIN4(n2024), .DIN5(
        n2026), .Q(n1965) );
  xor2s3 U1406 ( .DIN1(n2682), .DIN2(n2683), .Q(n2026) );
  xor2s3 U1407 ( .DIN1(n2684), .DIN2(n2685), .Q(n2024) );
  xor2s3 U1408 ( .DIN1(n2688), .DIN2(n2689), .Q(n2006) );
  xor2s3 U1409 ( .DIN1(n2690), .DIN2(n2691), .Q(n2005) );
  xor2s3 U1410 ( .DIN1(n2686), .DIN2(n2687), .Q(n2004) );
  or2s3 U1411 ( .DIN1(n1837), .DIN2(n2871), .Q(n1943) );
  nnd2s3 U1412 ( .DIN1(n2027), .DIN2(n2042), .Q(g11338) );
  nnd2s3 U1413 ( .DIN1(n2837), .DIN2(n640), .Q(n2042) );
  nnd2s3 U1414 ( .DIN1(n2828), .DIN2(n737), .Q(n2027) );
  nnd2s3 U1415 ( .DIN1(n2059), .DIN2(n2060), .Q(g11337) );
  nnd2s3 U1416 ( .DIN1(n2837), .DIN2(n737), .Q(n2060) );
  nnd2s3 U1417 ( .DIN1(n2828), .DIN2(n525), .Q(n2059) );
  nnd2s3 U1418 ( .DIN1(n2062), .DIN2(n2063), .Q(g11336) );
  nnd2s3 U1419 ( .DIN1(n2837), .DIN2(n525), .Q(n2063) );
  nnd2s3 U1420 ( .DIN1(n2828), .DIN2(n583), .Q(n2062) );
  nnd2s3 U1421 ( .DIN1(n2064), .DIN2(n2065), .Q(g11335) );
  nnd2s3 U1422 ( .DIN1(n2838), .DIN2(n583), .Q(n2065) );
  nnd2s3 U1423 ( .DIN1(n2828), .DIN2(n748), .Q(n2064) );
  nnd2s3 U1424 ( .DIN1(n2066), .DIN2(n2067), .Q(g11334) );
  nnd2s3 U1425 ( .DIN1(n2838), .DIN2(n748), .Q(n2067) );
  nnd2s3 U1426 ( .DIN1(n2828), .DIN2(n843), .Q(n2066) );
  nnd2s3 U1427 ( .DIN1(n2068), .DIN2(n2069), .Q(g11333) );
  nnd2s3 U1428 ( .DIN1(n2838), .DIN2(n843), .Q(n2069) );
  nnd2s3 U1429 ( .DIN1(n2828), .DIN2(n678), .Q(n2068) );
  nnd2s3 U1430 ( .DIN1(n2070), .DIN2(n2071), .Q(g11332) );
  nnd2s3 U1431 ( .DIN1(n2838), .DIN2(n678), .Q(n2071) );
  nnd2s3 U1432 ( .DIN1(n2828), .DIN2(n790), .Q(n2070) );
  nnd2s3 U1433 ( .DIN1(n2072), .DIN2(n2075), .Q(g11331) );
  nnd2s3 U1434 ( .DIN1(n2838), .DIN2(n790), .Q(n2075) );
  nnd2s3 U1435 ( .DIN1(n2828), .DIN2(n609), .Q(n2072) );
  nnd2s3 U1436 ( .DIN1(n2076), .DIN2(n2077), .Q(g11330) );
  nnd2s3 U1437 ( .DIN1(n2839), .DIN2(n598), .Q(n2077) );
  nnd2s3 U1438 ( .DIN1(n2828), .DIN2(n573), .Q(n2076) );
  nnd2s3 U1439 ( .DIN1(n2078), .DIN2(n2079), .Q(g11329) );
  nnd2s3 U1440 ( .DIN1(n2839), .DIN2(n573), .Q(n2079) );
  nnd2s3 U1441 ( .DIN1(n2828), .DIN2(n754), .Q(n2078) );
  nnd2s3 U1442 ( .DIN1(n2080), .DIN2(n2081), .Q(g11328) );
  nnd2s3 U1443 ( .DIN1(n2839), .DIN2(n754), .Q(n2081) );
  nnd2s3 U1444 ( .DIN1(n2828), .DIN2(n533), .Q(n2080) );
  nnd2s3 U1445 ( .DIN1(n2082), .DIN2(n2083), .Q(g11327) );
  nnd2s3 U1446 ( .DIN1(n2833), .DIN2(n533), .Q(n2083) );
  nnd2s3 U1447 ( .DIN1(n2828), .DIN2(n761), .Q(n2082) );
  nnd2s3 U1448 ( .DIN1(n2084), .DIN2(n2085), .Q(g11326) );
  nnd2s3 U1449 ( .DIN1(n2834), .DIN2(n761), .Q(n2085) );
  nnd2s3 U1450 ( .DIN1(n2829), .DIN2(n759), .Q(n2084) );
  nnd2s3 U1451 ( .DIN1(n2086), .DIN2(n2087), .Q(g11325) );
  nnd2s3 U1452 ( .DIN1(n2834), .DIN2(n759), .Q(n2087) );
  nnd2s3 U1453 ( .DIN1(n2829), .DIN2(n640), .Q(n2086) );
  nnd2s3 U1454 ( .DIN1(n2088), .DIN2(n2089), .Q(g11324) );
  nnd2s3 U1455 ( .DIN1(n1702), .DIN2(n2830), .Q(n2089) );
  nnd2s3 U1456 ( .DIN1(n2090), .DIN2(n2091), .Q(n1702) );
  nnd2s3 U1457 ( .DIN1(n2053), .DIN2(n2092), .Q(n2091) );
  nnd2s3 U1458 ( .DIN1(n2032), .DIN2(n2093), .Q(n2092) );
  or5s3 U1459 ( .DIN1(n533), .DIN2(n761), .DIN3(n759), .DIN4(n2094), .DIN5(
        n2095), .Q(n2093) );
  nnd4s2 U1460 ( .DIN1(n2641), .DIN2(n2630), .DIN3(n2637), .DIN4(n2096), .Q(
        n2095) );
  and4s2 U1461 ( .DIN1(n2639), .DIN2(n2638), .DIN3(n2636), .DIN4(n2640), .Q(
        n2096) );
  nnd3s3 U1462 ( .DIN1(n2631), .DIN2(n2629), .DIN3(n2635), .Q(n2094) );
  nnd2s3 U1463 ( .DIN1(n2032), .DIN2(n598), .Q(n2090) );
  nnd2s3 U1464 ( .DIN1(n2835), .DIN2(n609), .Q(n2088) );
  nnd2s3 U1465 ( .DIN1(n2097), .DIN2(n2098), .Q(g11270) );
  nnd2s3 U1466 ( .DIN1(n2835), .DIN2(n626), .Q(n2098) );
  nnd2s3 U1467 ( .DIN1(n2829), .DIN2(n760), .Q(n2097) );
  nnd2s3 U1468 ( .DIN1(n2099), .DIN2(n2100), .Q(g11269) );
  nnd2s3 U1469 ( .DIN1(n2835), .DIN2(n760), .Q(n2100) );
  nnd2s3 U1470 ( .DIN1(n2829), .DIN2(n562), .Q(n2099) );
  nnd2s3 U1471 ( .DIN1(n2101), .DIN2(n2102), .Q(g11268) );
  nnd2s3 U1472 ( .DIN1(n2835), .DIN2(n562), .Q(n2102) );
  nnd2s3 U1473 ( .DIN1(n2829), .DIN2(n617), .Q(n2101) );
  nnd2s3 U1474 ( .DIN1(n2103), .DIN2(n2104), .Q(g11267) );
  nnd2s3 U1475 ( .DIN1(n2835), .DIN2(n617), .Q(n2104) );
  nnd2s3 U1476 ( .DIN1(n2829), .DIN2(n777), .Q(n2103) );
  nnd2s3 U1477 ( .DIN1(n2105), .DIN2(n2106), .Q(g11266) );
  nnd2s3 U1478 ( .DIN1(n2836), .DIN2(n777), .Q(n2106) );
  nnd2s3 U1479 ( .DIN1(n2829), .DIN2(n807), .Q(n2105) );
  nnd2s3 U1480 ( .DIN1(n2107), .DIN2(n2108), .Q(g11265) );
  nnd2s3 U1481 ( .DIN1(n2836), .DIN2(n807), .Q(n2108) );
  nnd2s3 U1482 ( .DIN1(n2829), .DIN2(n634), .Q(n2107) );
  nnd2s3 U1483 ( .DIN1(n2109), .DIN2(n2110), .Q(g11264) );
  nnd2s3 U1484 ( .DIN1(n2836), .DIN2(n634), .Q(n2110) );
  nnd2s3 U1485 ( .DIN1(n2829), .DIN2(n750), .Q(n2109) );
  nnd2s3 U1486 ( .DIN1(n2111), .DIN2(n2112), .Q(g11263) );
  nnd2s3 U1487 ( .DIN1(n2836), .DIN2(n750), .Q(n2112) );
  nnd2s3 U1488 ( .DIN1(n2829), .DIN2(n804), .Q(n2111) );
  nnd2s3 U1489 ( .DIN1(n2113), .DIN2(n2114), .Q(g11262) );
  nnd2s3 U1490 ( .DIN1(n2837), .DIN2(n561), .Q(n2114) );
  nnd2s3 U1491 ( .DIN1(n2829), .DIN2(n546), .Q(n2113) );
  nnd2s3 U1492 ( .DIN1(n2115), .DIN2(n2116), .Q(g11261) );
  nnd2s3 U1493 ( .DIN1(n2836), .DIN2(n546), .Q(n2116) );
  nnd2s3 U1494 ( .DIN1(n2829), .DIN2(n641), .Q(n2115) );
  nnd2s3 U1495 ( .DIN1(n2117), .DIN2(n2118), .Q(g11260) );
  nnd2s3 U1496 ( .DIN1(n2833), .DIN2(n641), .Q(n2118) );
  nnd2s3 U1497 ( .DIN1(n2830), .DIN2(n781), .Q(n2117) );
  nnd2s3 U1498 ( .DIN1(n2119), .DIN2(n2120), .Q(g11259) );
  nnd2s3 U1499 ( .DIN1(n2833), .DIN2(n781), .Q(n2120) );
  nnd2s3 U1500 ( .DIN1(n2829), .DIN2(n653), .Q(n2119) );
  nnd2s3 U1501 ( .DIN1(n2121), .DIN2(n2122), .Q(g11258) );
  nnd2s3 U1502 ( .DIN1(n2834), .DIN2(n653), .Q(n2122) );
  nnd2s3 U1503 ( .DIN1(n2830), .DIN2(n870), .Q(n2121) );
  nnd2s3 U1504 ( .DIN1(n2123), .DIN2(n2124), .Q(g11257) );
  nnd2s3 U1505 ( .DIN1(n2834), .DIN2(n870), .Q(n2124) );
  nnd2s3 U1506 ( .DIN1(n2830), .DIN2(n626), .Q(n2123) );
  nnd2s3 U1507 ( .DIN1(n2125), .DIN2(n2126), .Q(g11256) );
  nnd2s3 U1508 ( .DIN1(n2003), .DIN2(n2830), .Q(n2126) );
  nnd2s3 U1509 ( .DIN1(n2127), .DIN2(n2128), .Q(n2003) );
  nnd2s3 U1510 ( .DIN1(n2129), .DIN2(n2130), .Q(n2128) );
  nnd2s3 U1511 ( .DIN1(n2131), .DIN2(n2132), .Q(n2130) );
  nnd2s3 U1512 ( .DIN1(n2054), .DIN2(n2133), .Q(n2132) );
  nnd2s3 U1513 ( .DIN1(n2033), .DIN2(n2134), .Q(n2133) );
  or5s3 U1514 ( .DIN1(n641), .DIN2(n781), .DIN3(n653), .DIN4(n2135), .DIN5(
        n2136), .Q(n2134) );
  nnd4s2 U1515 ( .DIN1(n2674), .DIN2(n2683), .DIN3(n2681), .DIN4(n2137), .Q(
        n2136) );
  and4s2 U1516 ( .DIN1(n2685), .DIN2(n2689), .DIN3(n2691), .DIN4(n2687), .Q(
        n2137) );
  nnd3s3 U1517 ( .DIN1(n2676), .DIN2(n2677), .DIN3(n2675), .Q(n2135) );
  nnd2s3 U1518 ( .DIN1(n2033), .DIN2(n561), .Q(n2131) );
  nnd2s3 U1519 ( .DIN1(n568), .DIN2(n724), .Q(n2127) );
  nor2s3 U1520 ( .DIN1(n1867), .DIN2(n2670), .Q(n2129) );
  or3s3 U1521 ( .DIN1(n2672), .DIN2(n2671), .DIN3(n2673), .Q(n1867) );
  nnd2s3 U1522 ( .DIN1(n2837), .DIN2(n804), .Q(n2125) );
  or5s3 U1523 ( .DIN1(n692), .DIN2(n840), .DIN3(n654), .DIN4(n2138), .DIN5(
        n2139), .Q(n1701) );
  or5s3 U1524 ( .DIN1(n736), .DIN2(n627), .DIN3(n605), .DIN4(n671), .DIN5(n622), .Q(n2139) );
  nnd3s3 U1525 ( .DIN1(g109), .DIN2(n2140), .DIN3(n2664), .Q(n2138) );
  or5s3 U1526 ( .DIN1(n2821), .DIN2(n2822), .DIN3(n2818), .DIN4(n2820), .DIN5(
        n2141), .Q(n2140) );
  nnd4s2 U1527 ( .DIN1(n577), .DIN2(n571), .DIN3(n569), .DIN4(n553), .Q(n2141)
         );
  and2s3 U1528 ( .DIN1(g10628), .DIN2(n2142), .Q(g11206) );
  nnd2s3 U1529 ( .DIN1(n2143), .DIN2(n2144), .Q(g11185) );
  or2s3 U1530 ( .DIN1(n2145), .DIN2(n1398), .Q(n2144) );
  nor6s3 U1531 ( .DIN1(n2821), .DIN2(n2818), .DIN3(n2820), .DIN4(n1907), 
        .DIN5(n553), .DIN6(n2146), .Q(n2145) );
  nor2s3 U1532 ( .DIN1(g6262), .DIN2(n2147), .Q(n2146) );
  nnd2s3 U1533 ( .DIN1(n1398), .DIN2(n616), .Q(n2143) );
  nor2s3 U1534 ( .DIN1(n646), .DIN2(n576), .Q(g11184) );
  nor2s3 U1535 ( .DIN1(n646), .DIN2(n615), .Q(g11183) );
  nor2s3 U1536 ( .DIN1(n646), .DIN2(n860), .Q(g11182) );
  nor2s3 U1537 ( .DIN1(n646), .DIN2(n550), .Q(g11181) );
  nnd2s3 U1538 ( .DIN1(g1696), .DIN2(n2725), .Q(n1398) );
  nnd2s3 U1539 ( .DIN1(n2148), .DIN2(n2149), .Q(g11180) );
  nnd2s3 U1540 ( .DIN1(n2848), .DIN2(n2150), .Q(n2149) );
  nnd2s3 U1541 ( .DIN1(n2151), .DIN2(n1677), .Q(n2150) );
  nnd2s3 U1542 ( .DIN1(n1766), .DIN2(n577), .Q(n1677) );
  nnd2s3 U1543 ( .DIN1(n895), .DIN2(n902), .Q(n1766) );
  nnd3s3 U1544 ( .DIN1(g6257), .DIN2(n901), .DIN3(n943), .Q(n2147) );
  nor5s3 U1545 ( .DIN1(g6263), .DIN2(g6260), .DIN3(g6259), .DIN4(g6258), 
        .DIN5(n908), .Q(n943) );
  xor2s3 U1546 ( .DIN1(n2152), .DIN2(n2153), .Q(n2151) );
  xor2s3 U1547 ( .DIN1(n2154), .DIN2(n2155), .Q(n2153) );
  xor2s3 U1548 ( .DIN1(n2156), .DIN2(n2157), .Q(n2155) );
  xor2s3 U1549 ( .DIN1(n2655), .DIN2(n2816), .Q(n2157) );
  xor2s3 U1550 ( .DIN1(n2653), .DIN2(n2654), .Q(n2156) );
  xor2s3 U1551 ( .DIN1(n2158), .DIN2(n2159), .Q(n2154) );
  xor2s3 U1552 ( .DIN1(n2651), .DIN2(n2652), .Q(n2159) );
  xor2s3 U1553 ( .DIN1(n2649), .DIN2(n2650), .Q(n2158) );
  xnr2s3 U1554 ( .DIN1(n2648), .DIN2(n2647), .Q(n2152) );
  or2s3 U1555 ( .DIN1(n2850), .DIN2(n2726), .Q(n2148) );
  xor2s3 U1556 ( .DIN1(n2819), .DIN2(n2142), .Q(g11163) );
  and2s3 U1557 ( .DIN1(n2160), .DIN2(n2161), .Q(n2142) );
  nnd2s3 U1558 ( .DIN1(g109), .DIN2(n2162), .Q(n2161) );
  nnd4s2 U1559 ( .DIN1(n2163), .DIN2(n2164), .DIN3(n2165), .DIN4(n2166), .Q(
        n2162) );
  nnd2s3 U1560 ( .DIN1(n679), .DIN2(n2822), .Q(n2166) );
  nnd3s3 U1561 ( .DIN1(\DFF_194/net481 ), .DIN2(g3069), .DIN3(g109), .Q(n1669)
         );
  nnd2s3 U1562 ( .DIN1(n2726), .DIN2(n2825), .Q(n2165) );
  or2s3 U1563 ( .DIN1(n553), .DIN2(n2011), .Q(n2164) );
  nnd2s3 U1564 ( .DIN1(n2824), .DIN2(g2648), .Q(n2163) );
  nnd2s3 U1565 ( .DIN1(g6846), .DIN2(g10774), .Q(n2160) );
  nor2s3 U1566 ( .DIN1(n1638), .DIN2(n2865), .Q(g6846) );
  nnd2s3 U1567 ( .DIN1(n684), .DIN2(g1765), .Q(n1638) );
  nnd2s3 U1568 ( .DIN1(n2167), .DIN2(n2168), .Q(g11052) );
  nnd2s3 U1569 ( .DIN1(n2848), .DIN2(n2169), .Q(n2168) );
  nnd2s3 U1570 ( .DIN1(n2854), .DIN2(n753), .Q(n2167) );
  nnd2s3 U1571 ( .DIN1(n2170), .DIN2(n2171), .Q(g11051) );
  nnd2s3 U1572 ( .DIN1(n2854), .DIN2(n709), .Q(n2171) );
  nnd2s3 U1573 ( .DIN1(n2172), .DIN2(n2173), .Q(g11050) );
  nnd2s3 U1574 ( .DIN1(n2854), .DIN2(n756), .Q(n2172) );
  nnd2s3 U1575 ( .DIN1(n2174), .DIN2(n2175), .Q(g11049) );
  nnd2s3 U1576 ( .DIN1(n2854), .DIN2(n729), .Q(n2175) );
  nnd2s3 U1577 ( .DIN1(n2176), .DIN2(n2177), .Q(g11048) );
  nnd2s3 U1578 ( .DIN1(n2855), .DIN2(n771), .Q(n2177) );
  nnd2s3 U1579 ( .DIN1(n2178), .DIN2(n2179), .Q(g11047) );
  nnd2s3 U1580 ( .DIN1(n2855), .DIN2(n844), .Q(n2179) );
  nnd2s3 U1581 ( .DIN1(n2180), .DIN2(n2181), .Q(g11044) );
  nnd2s3 U1582 ( .DIN1(n2848), .DIN2(n2182), .Q(n2181) );
  nnd2s3 U1583 ( .DIN1(n2855), .DIN2(n786), .Q(n2180) );
  nnd2s3 U1584 ( .DIN1(n2183), .DIN2(n2184), .Q(g11043) );
  nnd2s3 U1585 ( .DIN1(n2855), .DIN2(n582), .Q(n2183) );
  nnd2s3 U1586 ( .DIN1(n2170), .DIN2(n2185), .Q(g11042) );
  nnd2s3 U1587 ( .DIN1(n2856), .DIN2(n579), .Q(n2185) );
  nnd2s3 U1588 ( .DIN1(n2848), .DIN2(n2186), .Q(n2170) );
  nnd2s3 U1589 ( .DIN1(n2187), .DIN2(n2188), .Q(n2186) );
  nnd2s3 U1590 ( .DIN1(n738), .DIN2(n1269), .Q(n2188) );
  nnd2s3 U1591 ( .DIN1(n1152), .DIN2(n2189), .Q(n1269) );
  nnd2s3 U1592 ( .DIN1(n2862), .DIN2(n735), .Q(n2189) );
  nnd2s3 U1593 ( .DIN1(g2355), .DIN2(n772), .Q(n1152) );
  nnd2s3 U1594 ( .DIN1(n2190), .DIN2(n2191), .Q(n2187) );
  nnd2s3 U1595 ( .DIN1(g109), .DIN2(n571), .Q(n2191) );
  nnd2s3 U1596 ( .DIN1(n2192), .DIN2(n2173), .Q(g11041) );
  nnd2s3 U1597 ( .DIN1(n2848), .DIN2(n2193), .Q(n2173) );
  nnd2s3 U1598 ( .DIN1(n2194), .DIN2(n2195), .Q(n2193) );
  nnd2s3 U1599 ( .DIN1(n738), .DIN2(n1267), .Q(n2195) );
  nnd2s3 U1600 ( .DIN1(n1160), .DIN2(n2196), .Q(n1267) );
  nnd2s3 U1601 ( .DIN1(n2862), .DIN2(n643), .Q(n2196) );
  nnd2s3 U1602 ( .DIN1(g2355), .DIN2(n799), .Q(n1160) );
  nnd2s3 U1603 ( .DIN1(n2190), .DIN2(n1907), .Q(n2194) );
  nnd2s3 U1604 ( .DIN1(n2855), .DIN2(n829), .Q(n2192) );
  nnd2s3 U1605 ( .DIN1(n2174), .DIN2(n2197), .Q(g11040) );
  nnd2s3 U1606 ( .DIN1(n2856), .DIN2(n758), .Q(n2197) );
  nnd4s2 U1607 ( .DIN1(n2850), .DIN2(n2198), .DIN3(n2199), .DIN4(n2200), .Q(
        n2174) );
  nnd2s3 U1608 ( .DIN1(n738), .DIN2(n1265), .Q(n2199) );
  nnd2s3 U1609 ( .DIN1(n2201), .DIN2(n2202), .Q(n1265) );
  nnd2s3 U1610 ( .DIN1(n2705), .DIN2(n2863), .Q(n2202) );
  nnd2s3 U1611 ( .DIN1(g2355), .DIN2(n1972), .Q(n2201) );
  nnd2s3 U1612 ( .DIN1(n2203), .DIN2(n553), .Q(n2198) );
  nnd2s3 U1613 ( .DIN1(n2176), .DIN2(n2204), .Q(g11039) );
  nnd2s3 U1614 ( .DIN1(n2856), .DIN2(n815), .Q(n2204) );
  nnd4s2 U1615 ( .DIN1(n2850), .DIN2(n2205), .DIN3(n2206), .DIN4(n2200), .Q(
        n2176) );
  nnd2s3 U1616 ( .DIN1(n738), .DIN2(n1263), .Q(n2206) );
  nnd2s3 U1617 ( .DIN1(n2207), .DIN2(n2208), .Q(n1263) );
  nnd2s3 U1618 ( .DIN1(n2707), .DIN2(n2862), .Q(n2208) );
  nnd2s3 U1619 ( .DIN1(g2355), .DIN2(n1962), .Q(n2207) );
  nnd2s3 U1620 ( .DIN1(n2203), .DIN2(n526), .Q(n2205) );
  nnd2s3 U1621 ( .DIN1(n2178), .DIN2(n2209), .Q(g11038) );
  nnd2s3 U1622 ( .DIN1(n2856), .DIN2(n832), .Q(n2209) );
  nnd3s3 U1623 ( .DIN1(n2210), .DIN2(n2211), .DIN3(n2848), .Q(n2178) );
  nnd3s3 U1624 ( .DIN1(g109), .DIN2(n523), .DIN3(n2190), .Q(n2211) );
  nnd2s3 U1625 ( .DIN1(n738), .DIN2(n1261), .Q(n2210) );
  nnd2s3 U1626 ( .DIN1(n2212), .DIN2(n2213), .Q(n1261) );
  nnd2s3 U1627 ( .DIN1(n2709), .DIN2(n2863), .Q(n2213) );
  nnd2s3 U1628 ( .DIN1(g2355), .DIN2(n2001), .Q(n2212) );
  nnd2s3 U1629 ( .DIN1(n2214), .DIN2(n2184), .Q(g11037) );
  nnd2s3 U1630 ( .DIN1(n2848), .DIN2(n2215), .Q(n2184) );
  nnd2s3 U1631 ( .DIN1(n2216), .DIN2(n2217), .Q(n2215) );
  nnd3s3 U1632 ( .DIN1(g109), .DIN2(n2821), .DIN3(n2190), .Q(n2217) );
  nnd2s3 U1633 ( .DIN1(n738), .DIN2(n1259), .Q(n2216) );
  nnd2s3 U1634 ( .DIN1(n1187), .DIN2(n2218), .Q(n1259) );
  nnd2s3 U1635 ( .DIN1(n2862), .DIN2(n549), .Q(n2218) );
  nnd2s3 U1636 ( .DIN1(g2355), .DIN2(n811), .Q(n1187) );
  nnd2s3 U1637 ( .DIN1(n2857), .DIN2(n858), .Q(n2214) );
  nnd2s3 U1638 ( .DIN1(n2219), .DIN2(n2220), .Q(g11036) );
  nnd3s3 U1639 ( .DIN1(n1601), .DIN2(n2221), .DIN3(n2190), .Q(n2220) );
  nnd2s3 U1640 ( .DIN1(g109), .DIN2(n553), .Q(n2221) );
  nnd2s3 U1641 ( .DIN1(n650), .DIN2(n785), .Q(n2219) );
  nnd2s3 U1642 ( .DIN1(n2222), .DIN2(n2223), .Q(g11035) );
  nnd2s3 U1643 ( .DIN1(n1601), .DIN2(n2224), .Q(n2223) );
  nnd2s3 U1644 ( .DIN1(n1979), .DIN2(n2225), .Q(n2224) );
  nnd2s3 U1645 ( .DIN1(n2226), .DIN2(n2820), .Q(n2225) );
  nnd2s3 U1646 ( .DIN1(n650), .DIN2(n554), .Q(n2222) );
  nnd2s3 U1647 ( .DIN1(n2227), .DIN2(n2228), .Q(g11034) );
  nnd2s3 U1648 ( .DIN1(n1601), .DIN2(n2182), .Q(n2228) );
  nnd3s3 U1649 ( .DIN1(n2229), .DIN2(n2230), .DIN3(n1979), .Q(n2182) );
  nnd2s3 U1650 ( .DIN1(n2226), .DIN2(n2818), .Q(n2230) );
  nnd2s3 U1651 ( .DIN1(n738), .DIN2(n1277), .Q(n2229) );
  nnd2s3 U1652 ( .DIN1(n1473), .DIN2(n2231), .Q(n1277) );
  nnd2s3 U1653 ( .DIN1(n2862), .DIN2(n604), .Q(n2231) );
  nnd2s3 U1654 ( .DIN1(g2355), .DIN2(n712), .Q(n1473) );
  nnd2s3 U1655 ( .DIN1(n650), .DIN2(n716), .Q(n2227) );
  nnd2s3 U1656 ( .DIN1(n2232), .DIN2(n2233), .Q(g11033) );
  nnd2s3 U1657 ( .DIN1(n1601), .DIN2(n2169), .Q(n2233) );
  nnd3s3 U1658 ( .DIN1(n2234), .DIN2(n2200), .DIN3(n2235), .Q(n2169) );
  nnd2s3 U1659 ( .DIN1(n2203), .DIN2(n2821), .Q(n2235) );
  nnd2s3 U1660 ( .DIN1(n2203), .DIN2(n2236), .Q(n2200) );
  nnd2s3 U1661 ( .DIN1(n1979), .DIN2(g109), .Q(n2236) );
  nnd2s3 U1662 ( .DIN1(n738), .DIN2(n1275), .Q(n2234) );
  nnd2s3 U1663 ( .DIN1(n1463), .DIN2(n2237), .Q(n1275) );
  nnd2s3 U1664 ( .DIN1(n2862), .DIN2(n628), .Q(n2237) );
  nnd2s3 U1665 ( .DIN1(g2355), .DIN2(n827), .Q(n1463) );
  nnd2s3 U1666 ( .DIN1(n650), .DIN2(n848), .Q(n2232) );
  nnd2s3 U1667 ( .DIN1(n2238), .DIN2(n2239), .Q(g10882) );
  nnd2s3 U1668 ( .DIN1(n1596), .DIN2(n1907), .Q(n2239) );
  nnd2s3 U1669 ( .DIN1(g109), .DIN2(n547), .Q(n1907) );
  nnd2s3 U1670 ( .DIN1(n647), .DIN2(n686), .Q(n2238) );
  nnd2s3 U1671 ( .DIN1(n2240), .DIN2(n2241), .Q(g10881) );
  nnd2s3 U1672 ( .DIN1(n2242), .DIN2(n2823), .Q(n2241) );
  or2s3 U1673 ( .DIN1(n1596), .DIN2(n2752), .Q(n2240) );
  nnd2s3 U1674 ( .DIN1(n2243), .DIN2(n2244), .Q(g10880) );
  nnd2s3 U1675 ( .DIN1(n2242), .DIN2(n2820), .Q(n2244) );
  or2s3 U1676 ( .DIN1(n1596), .DIN2(n2766), .Q(n2243) );
  nnd2s3 U1677 ( .DIN1(n2245), .DIN2(n2246), .Q(g10879) );
  nnd2s3 U1678 ( .DIN1(n2242), .DIN2(n2818), .Q(n2246) );
  or2s3 U1679 ( .DIN1(n1596), .DIN2(n2778), .Q(n2245) );
  nnd2s3 U1680 ( .DIN1(n2247), .DIN2(n2248), .Q(g10878) );
  nnd2s3 U1681 ( .DIN1(n2242), .DIN2(n2821), .Q(n2248) );
  nor2s3 U1682 ( .DIN1(n647), .DIN2(n2865), .Q(n2242) );
  or2s3 U1683 ( .DIN1(n1596), .DIN2(n2792), .Q(n2247) );
  nor2s3 U1684 ( .DIN1(n872), .DIN2(n2725), .Q(n1596) );
  nnd2s3 U1685 ( .DIN1(n2249), .DIN2(n2250), .Q(g10877) );
  nnd2s3 U1686 ( .DIN1(n2856), .DIN2(n784), .Q(n2250) );
  nnd2s3 U1687 ( .DIN1(n2848), .DIN2(n2251), .Q(n2249) );
  nnd2s3 U1688 ( .DIN1(n2252), .DIN2(n2253), .Q(g10876) );
  nnd2s3 U1689 ( .DIN1(n2852), .DIN2(n529), .Q(n2253) );
  nnd2s3 U1690 ( .DIN1(n2848), .DIN2(n2254), .Q(n2252) );
  nnd2s3 U1691 ( .DIN1(n2725), .DIN2(n872), .Q(n1149) );
  nnd2s3 U1692 ( .DIN1(n2255), .DIN2(n2256), .Q(g10875) );
  nnd2s3 U1693 ( .DIN1(n1601), .DIN2(n2251), .Q(n2256) );
  nnd3s3 U1694 ( .DIN1(n2257), .DIN2(n2258), .DIN3(n1979), .Q(n2251) );
  nnd2s3 U1695 ( .DIN1(n2226), .DIN2(n2824), .Q(n2258) );
  nor2s3 U1696 ( .DIN1(n2870), .DIN2(n738), .Q(n2226) );
  nnd2s3 U1697 ( .DIN1(n738), .DIN2(n1273), .Q(n2257) );
  nnd2s3 U1698 ( .DIN1(n1465), .DIN2(n2259), .Q(n1273) );
  nnd2s3 U1699 ( .DIN1(n2861), .DIN2(n764), .Q(n2259) );
  nnd2s3 U1700 ( .DIN1(g2355), .DIN2(n853), .Q(n1465) );
  nnd2s3 U1701 ( .DIN1(n650), .DIN2(n711), .Q(n2255) );
  nnd2s3 U1702 ( .DIN1(n2260), .DIN2(n2261), .Q(g10874) );
  nnd2s3 U1703 ( .DIN1(n1601), .DIN2(n2254), .Q(n2261) );
  nnd2s3 U1704 ( .DIN1(n2262), .DIN2(n2263), .Q(n2254) );
  nnd2s3 U1705 ( .DIN1(n2190), .DIN2(n2264), .Q(n2263) );
  nnd2s3 U1706 ( .DIN1(g109), .DIN2(n577), .Q(n2264) );
  and2s3 U1707 ( .DIN1(n1979), .DIN2(n2203), .Q(n2190) );
  nnd2s3 U1708 ( .DIN1(n738), .DIN2(n1271), .Q(n2262) );
  nnd2s3 U1709 ( .DIN1(n1144), .DIN2(n2265), .Q(n1271) );
  nnd2s3 U1710 ( .DIN1(n2862), .DIN2(n558), .Q(n2265) );
  nnd2s3 U1711 ( .DIN1(g2355), .DIN2(n697), .Q(n1144) );
  nnd2s3 U1712 ( .DIN1(n2724), .DIN2(n1979), .Q(n2203) );
  nnd2s3 U1713 ( .DIN1(n650), .DIN2(n614), .Q(n2260) );
  nor2s3 U1714 ( .DIN1(n2725), .DIN2(g1696), .Q(n1601) );
  nnd2s3 U1715 ( .DIN1(n2266), .DIN2(n522), .Q(g10801) );
  xor2s3 U1716 ( .DIN1(n2267), .DIN2(n2268), .Q(n2819) );
  xor2s3 U1717 ( .DIN1(n2269), .DIN2(n2270), .Q(n2268) );
  xor2s3 U1718 ( .DIN1(n2271), .DIN2(n2272), .Q(n2270) );
  xor2s3 U1719 ( .DIN1(n553), .DIN2(n547), .Q(n2272) );
  xor2s3 U1720 ( .DIN1(n2825), .DIN2(n577), .Q(n2271) );
  xor2s3 U1721 ( .DIN1(n2273), .DIN2(n2274), .Q(n2269) );
  xor2s3 U1722 ( .DIN1(n2824), .DIN2(n2821), .Q(n2274) );
  xor2s3 U1723 ( .DIN1(n2818), .DIN2(n526), .Q(n2273) );
  nnd2s3 U1724 ( .DIN1(n2030), .DIN2(n896), .Q(n2267) );
  nnd2s3 U1725 ( .DIN1(g109), .DIN2(n2275), .Q(g10628) );
  or5s3 U1726 ( .DIN1(n2276), .DIN2(n2277), .DIN3(n2278), .DIN4(n2279), .DIN5(
        n2280), .Q(n2275) );
  and2s3 U1727 ( .DIN1(g877), .DIN2(n2821), .Q(n2280) );
  nor2s3 U1728 ( .DIN1(n523), .DIN2(n905), .Q(n2279) );
  nor2s3 U1729 ( .DIN1(n526), .DIN2(n1228), .Q(n2278) );
  nnd3s3 U1730 ( .DIN1(\DFF_121/net408 ), .DIN2(g2986), .DIN3(g109), .Q(n1228)
         );
  nor2s3 U1731 ( .DIN1(n553), .DIN2(n1836), .Q(n2277) );
  nnd2s3 U1732 ( .DIN1(g109), .DIN2(g757), .Q(n1836) );
  nor2s3 U1733 ( .DIN1(n547), .DIN2(n1837), .Q(n2276) );
  nnd2s3 U1734 ( .DIN1(g3007), .DIN2(\DFF_93/net380 ), .Q(n1837) );
  nnd2s3 U1735 ( .DIN1(n2266), .DIN2(n571), .Q(g10465) );
  or5s3 U1736 ( .DIN1(n2281), .DIN2(n2282), .DIN3(n2283), .DIN4(n2284), .DIN5(
        n2285), .Q(n2825) );
  nnd4s2 U1737 ( .DIN1(n2286), .DIN2(n2287), .DIN3(n2288), .DIN4(n2289), .Q(
        n2285) );
  and3s3 U1738 ( .DIN1(n2290), .DIN2(n2291), .DIN3(n2292), .Q(n2289) );
  nnd2s3 U1739 ( .DIN1(g4201), .DIN2(n2293), .Q(n2292) );
  nnd2s3 U1740 ( .DIN1(n881), .DIN2(n732), .Q(n2291) );
  nnd2s3 U1741 ( .DIN1(n882), .DIN2(n572), .Q(n2290) );
  nnd2s3 U1742 ( .DIN1(n892), .DIN2(n773), .Q(n2288) );
  nnd2s3 U1743 ( .DIN1(g4213), .DIN2(n2294), .Q(n2287) );
  nnd2s3 U1744 ( .DIN1(n888), .DIN2(n606), .Q(n2286) );
  nnd4s2 U1745 ( .DIN1(n2295), .DIN2(n2296), .DIN3(n2297), .DIN4(n2298), .Q(
        n2284) );
  nnd2s3 U1746 ( .DIN1(n2299), .DIN2(n680), .Q(n2298) );
  nnd2s3 U1747 ( .DIN1(n879), .DIN2(n800), .Q(n2297) );
  nnd2s3 U1748 ( .DIN1(n880), .DIN2(n847), .Q(n2296) );
  nnd2s3 U1749 ( .DIN1(n885), .DIN2(n825), .Q(n2295) );
  nor2s3 U1750 ( .DIN1(n894), .DIN2(n2300), .Q(n2283) );
  nor2s3 U1751 ( .DIN1(n2732), .DIN2(n2301), .Q(n2282) );
  nor2s3 U1752 ( .DIN1(n2733), .DIN2(n2302), .Q(n2281) );
  nnd2s3 U1753 ( .DIN1(n2266), .DIN2(n547), .Q(g10463) );
  or4s3 U1754 ( .DIN1(n2303), .DIN2(n2304), .DIN3(n2305), .DIN4(n2306), .Q(
        n2822) );
  nnd4s2 U1755 ( .DIN1(n2307), .DIN2(n2308), .DIN3(n2309), .DIN4(n2310), .Q(
        n2306) );
  nnd4s2 U1756 ( .DIN1(n878), .DIN2(n2311), .DIN3(n2312), .DIN4(n2313), .Q(
        n2310) );
  nnd2s3 U1757 ( .DIN1(n883), .DIN2(g16), .Q(n2309) );
  nnd2s3 U1758 ( .DIN1(n884), .DIN2(g7), .Q(n2308) );
  nnd2s3 U1759 ( .DIN1(n896), .DIN2(g37), .Q(n2307) );
  nnd4s2 U1760 ( .DIN1(n2314), .DIN2(n2315), .DIN3(n2316), .DIN4(n2317), .Q(
        n2305) );
  nnd2s3 U1761 ( .DIN1(n885), .DIN2(n623), .Q(n2317) );
  nnd2s3 U1762 ( .DIN1(n887), .DIN2(n686), .Q(n2316) );
  nnd2s3 U1763 ( .DIN1(n880), .DIN2(n636), .Q(n2315) );
  or2s3 U1764 ( .DIN1(n2302), .DIN2(n2745), .Q(n2314) );
  nnd4s2 U1765 ( .DIN1(n2319), .DIN2(n2320), .DIN3(n2321), .DIN4(n2322), .Q(
        n2304) );
  nnd2s3 U1766 ( .DIN1(n881), .DIN2(n861), .Q(n2322) );
  nnd2s3 U1767 ( .DIN1(n882), .DIN2(n823), .Q(n2321) );
  nnd2s3 U1768 ( .DIN1(n2299), .DIN2(n611), .Q(n2320) );
  nnd2s3 U1769 ( .DIN1(n879), .DIN2(n730), .Q(n2319) );
  nnd4s2 U1770 ( .DIN1(n2323), .DIN2(n2324), .DIN3(n2325), .DIN4(n2326), .Q(
        n2303) );
  nnd2s3 U1771 ( .DIN1(g4212), .DIN2(n2294), .Q(n2326) );
  nnd2s3 U1772 ( .DIN1(n888), .DIN2(n767), .Q(n2325) );
  nnd2s3 U1773 ( .DIN1(g4200), .DIN2(n2293), .Q(n2324) );
  nnd2s3 U1774 ( .DIN1(n892), .DIN2(n791), .Q(n2323) );
  nnd2s3 U1775 ( .DIN1(n2266), .DIN2(n553), .Q(g10461) );
  nnd3s3 U1776 ( .DIN1(n2327), .DIN2(n2328), .DIN3(n2329), .Q(n2823) );
  nor6s3 U1777 ( .DIN1(n2330), .DIN2(n2331), .DIN3(n2332), .DIN4(n2333), 
        .DIN5(n2334), .DIN6(n2335), .Q(n2329) );
  nor2s3 U1778 ( .DIN1(n2749), .DIN2(n2336), .Q(n2335) );
  and2s3 U1779 ( .DIN1(g4199), .DIN2(n2293), .Q(n2334) );
  nnd3s3 U1780 ( .DIN1(n2337), .DIN2(n2338), .DIN3(n2339), .Q(n2333) );
  nnd2s3 U1781 ( .DIN1(n891), .DIN2(n704), .Q(n2339) );
  nnd2s3 U1782 ( .DIN1(g4211), .DIN2(n2294), .Q(n2338) );
  nnd2s3 U1783 ( .DIN1(n888), .DIN2(n681), .Q(n2337) );
  and2s3 U1784 ( .DIN1(g4194), .DIN2(n2340), .Q(n2332) );
  nor2s3 U1785 ( .DIN1(n2045), .DIN2(n2341), .Q(n2331) );
  nnd3s3 U1786 ( .DIN1(n2342), .DIN2(n2343), .DIN3(n2344), .Q(n2330) );
  nnd2s3 U1787 ( .DIN1(g4208), .DIN2(n889), .Q(n2344) );
  nnd2s3 U1788 ( .DIN1(n883), .DIN2(g17), .Q(n2343) );
  nnd2s3 U1789 ( .DIN1(n884), .DIN2(g8), .Q(n2342) );
  nor6s3 U1790 ( .DIN1(n2345), .DIN2(n877), .DIN3(n2346), .DIN4(n2347), .DIN5(
        n2348), .DIN6(n2349), .Q(n2328) );
  nor2s3 U1791 ( .DIN1(n2758), .DIN2(n876), .Q(n2349) );
  nor2s3 U1792 ( .DIN1(n2757), .DIN2(n2350), .Q(n2348) );
  nor2s3 U1793 ( .DIN1(n2759), .DIN2(n2351), .Q(n2347) );
  nor2s3 U1794 ( .DIN1(n2756), .DIN2(n2352), .Q(n2346) );
  nor2s3 U1795 ( .DIN1(n2755), .DIN2(n2353), .Q(n2345) );
  nor5s3 U1796 ( .DIN1(n2354), .DIN2(n2355), .DIN3(n2356), .DIN4(n2357), 
        .DIN5(n2358), .Q(n2327) );
  nor2s3 U1797 ( .DIN1(n2752), .DIN2(n2359), .Q(n2358) );
  nor2s3 U1798 ( .DIN1(n2751), .DIN2(n2360), .Q(n2357) );
  nor2s3 U1799 ( .DIN1(n2753), .DIN2(n2318), .Q(n2356) );
  nor2s3 U1800 ( .DIN1(n2301), .DIN2(\DFF_228/net515 ), .Q(n2355) );
  nor2s3 U1801 ( .DIN1(n2754), .DIN2(n2302), .Q(n2354) );
  nnd2s3 U1802 ( .DIN1(n2266), .DIN2(n526), .Q(g10459) );
  nnd3s3 U1803 ( .DIN1(n2361), .DIN2(n2362), .DIN3(n2363), .Q(n2820) );
  nor6s3 U1804 ( .DIN1(n2364), .DIN2(n2365), .DIN3(n2366), .DIN4(n2367), 
        .DIN5(n2368), .DIN6(n2369), .Q(n2363) );
  nor2s3 U1805 ( .DIN1(n2761), .DIN2(n2336), .Q(n2369) );
  and2s3 U1806 ( .DIN1(g4198), .DIN2(n2293), .Q(n2368) );
  nnd3s3 U1807 ( .DIN1(n2370), .DIN2(n2371), .DIN3(n2372), .Q(n2367) );
  nnd2s3 U1808 ( .DIN1(n891), .DIN2(n842), .Q(n2372) );
  nnd2s3 U1809 ( .DIN1(g4210), .DIN2(n2294), .Q(n2371) );
  nnd2s3 U1810 ( .DIN1(n888), .DIN2(n584), .Q(n2370) );
  and2s3 U1811 ( .DIN1(g4193), .DIN2(n2340), .Q(n2366) );
  nor2s3 U1812 ( .DIN1(n2046), .DIN2(n2341), .Q(n2365) );
  nnd3s3 U1813 ( .DIN1(n2373), .DIN2(n2374), .DIN3(n2375), .Q(n2364) );
  nnd2s3 U1814 ( .DIN1(g4207), .DIN2(n889), .Q(n2375) );
  nnd2s3 U1815 ( .DIN1(n883), .DIN2(n775), .Q(n2374) );
  or2s3 U1816 ( .DIN1(n2313), .DIN2(n2764), .Q(n2373) );
  nor6s3 U1817 ( .DIN1(n2376), .DIN2(n877), .DIN3(n2377), .DIN4(n2378), .DIN5(
        n2379), .DIN6(n2380), .Q(n2362) );
  nor2s3 U1818 ( .DIN1(n2771), .DIN2(n876), .Q(n2380) );
  nor2s3 U1819 ( .DIN1(n2000), .DIN2(n2350), .Q(n2379) );
  nor2s3 U1820 ( .DIN1(n2772), .DIN2(n2351), .Q(n2378) );
  nor2s3 U1821 ( .DIN1(n2770), .DIN2(n2352), .Q(n2377) );
  nor2s3 U1822 ( .DIN1(n2769), .DIN2(n2353), .Q(n2376) );
  nor5s3 U1823 ( .DIN1(n2381), .DIN2(n2382), .DIN3(n2383), .DIN4(n2384), 
        .DIN5(n2385), .Q(n2361) );
  nor2s3 U1824 ( .DIN1(n2766), .DIN2(n2359), .Q(n2385) );
  nor2s3 U1825 ( .DIN1(n2765), .DIN2(n2360), .Q(n2384) );
  nor2s3 U1826 ( .DIN1(n2767), .DIN2(n2318), .Q(n2383) );
  nor2s3 U1827 ( .DIN1(n2301), .DIN2(\DFF_242/net529 ), .Q(n2382) );
  nor2s3 U1828 ( .DIN1(n2768), .DIN2(n2302), .Q(n2381) );
  nnd2s3 U1829 ( .DIN1(n2266), .DIN2(n523), .Q(g10457) );
  or5s3 U1830 ( .DIN1(n2386), .DIN2(n2387), .DIN3(n2388), .DIN4(n2389), .DIN5(
        n2390), .Q(n2818) );
  or5s3 U1831 ( .DIN1(n2391), .DIN2(n2392), .DIN3(n2393), .DIN4(n2394), .DIN5(
        n2395), .Q(n2390) );
  or5s3 U1832 ( .DIN1(n2396), .DIN2(n2397), .DIN3(n2398), .DIN4(n2399), .DIN5(
        n2400), .Q(n2395) );
  nor2s3 U1833 ( .DIN1(n2301), .DIN2(\DFF_384/net671 ), .Q(n2400) );
  nor2s3 U1834 ( .DIN1(n2780), .DIN2(n2302), .Q(n2399) );
  nor2s3 U1835 ( .DIN1(n2779), .DIN2(n2318), .Q(n2398) );
  nor2s3 U1836 ( .DIN1(n2778), .DIN2(n2359), .Q(n2397) );
  nor2s3 U1837 ( .DIN1(n2777), .DIN2(n2360), .Q(n2396) );
  nnd3s3 U1838 ( .DIN1(n2401), .DIN2(n2402), .DIN3(n2403), .Q(n2394) );
  nnd2s3 U1839 ( .DIN1(g4197), .DIN2(n2293), .Q(n2403) );
  nnd2s3 U1840 ( .DIN1(n881), .DIN2(n796), .Q(n2402) );
  nnd2s3 U1841 ( .DIN1(n882), .DIN2(n612), .Q(n2401) );
  nor2s3 U1842 ( .DIN1(n2783), .DIN2(n2351), .Q(n2393) );
  nor2s3 U1843 ( .DIN1(n2785), .DIN2(n876), .Q(n2392) );
  nor2s3 U1844 ( .DIN1(n2782), .DIN2(n2350), .Q(n2391) );
  nnd4s2 U1845 ( .DIN1(n2404), .DIN2(n2405), .DIN3(n2406), .DIN4(n2407), .Q(
        n2389) );
  and3s3 U1846 ( .DIN1(n2408), .DIN2(n2409), .DIN3(n2410), .Q(n2407) );
  nnd2s3 U1847 ( .DIN1(g4192), .DIN2(n2340), .Q(n2410) );
  or2s3 U1848 ( .DIN1(n2313), .DIN2(n2775), .Q(n2409) );
  nnd2s3 U1849 ( .DIN1(g4206), .DIN2(n889), .Q(n2408) );
  nnd2s3 U1850 ( .DIN1(n883), .DIN2(n524), .Q(n2406) );
  nnd2s3 U1851 ( .DIN1(g4196), .DIN2(n2411), .Q(n2404) );
  nnd3s3 U1852 ( .DIN1(n2412), .DIN2(n2413), .DIN3(n2414), .Q(n2388) );
  or2s3 U1853 ( .DIN1(n2341), .DIN2(n2007), .Q(n2414) );
  nnd2s3 U1854 ( .DIN1(g4209), .DIN2(n2294), .Q(n2413) );
  nnd2s3 U1855 ( .DIN1(n888), .DIN2(n597), .Q(n2412) );
  nor2s3 U1856 ( .DIN1(n2774), .DIN2(n2336), .Q(n2387) );
  nor2s3 U1857 ( .DIN1(n2044), .DIN2(n2415), .Q(n2386) );
  nnd2s3 U1858 ( .DIN1(n2266), .DIN2(n535), .Q(g10455) );
  nnd3s3 U1859 ( .DIN1(n2416), .DIN2(n2417), .DIN3(n2418), .Q(n2821) );
  nor6s3 U1860 ( .DIN1(n2419), .DIN2(n2420), .DIN3(n2421), .DIN4(n2422), 
        .DIN5(n2423), .DIN6(n2424), .Q(n2418) );
  nor2s3 U1861 ( .DIN1(n2047), .DIN2(n2341), .Q(n2424) );
  nor2s3 U1862 ( .DIN1(n2786), .DIN2(n2425), .Q(n2423) );
  and2s3 U1863 ( .DIN1(g4191), .DIN2(n2340), .Q(n2422) );
  nor2s3 U1864 ( .DIN1(n2788), .DIN2(n2336), .Q(n2421) );
  nor2s3 U1865 ( .DIN1(n2787), .DIN2(n2415), .Q(n2420) );
  nnd4s2 U1866 ( .DIN1(n2426), .DIN2(n2427), .DIN3(n2428), .DIN4(n2429), .Q(
        n2419) );
  and3s3 U1867 ( .DIN1(n2430), .DIN2(n2431), .DIN3(n2432), .Q(n2429) );
  nnd2s3 U1868 ( .DIN1(g4205), .DIN2(n2294), .Q(n2432) );
  nnd2s3 U1869 ( .DIN1(n884), .DIN2(n869), .Q(n2431) );
  nnd2s3 U1870 ( .DIN1(g4216), .DIN2(n889), .Q(n2430) );
  nnd2s3 U1871 ( .DIN1(n883), .DIN2(n639), .Q(n2428) );
  nnd2s3 U1872 ( .DIN1(n2790), .DIN2(n896), .Q(n2427) );
  nnd2s3 U1873 ( .DIN1(g4204), .DIN2(n2411), .Q(n2426) );
  nor6s3 U1874 ( .DIN1(n2434), .DIN2(n894), .DIN3(n877), .DIN4(n2435), .DIN5(
        n2436), .DIN6(n2437), .Q(n2417) );
  and2s3 U1875 ( .DIN1(g4195), .DIN2(n2293), .Q(n2437) );
  nor2s3 U1876 ( .DIN1(n2798), .DIN2(n2353), .Q(n2436) );
  nor2s3 U1877 ( .DIN1(n2796), .DIN2(n2350), .Q(n2435) );
  nnd4s2 U1878 ( .DIN1(n2311), .DIN2(n2312), .DIN3(n878), .DIN4(n2438), .Q(
        n2405) );
  and3s3 U1879 ( .DIN1(n2433), .DIN2(n2350), .DIN3(n2313), .Q(n2438) );
  nnd2s3 U1880 ( .DIN1(n2439), .DIN2(g6257), .Q(n2313) );
  nnd2s3 U1881 ( .DIN1(n2440), .DIN2(n890), .Q(n2433) );
  nnd2s3 U1882 ( .DIN1(n2439), .DIN2(n897), .Q(n2312) );
  and4s2 U1883 ( .DIN1(g6258), .DIN2(n2441), .DIN3(n899), .DIN4(n900), .Q(
        n2439) );
  nor2s3 U1884 ( .DIN1(n2795), .DIN2(n2352), .Q(n2434) );
  nor6s3 U1885 ( .DIN1(n2442), .DIN2(n2443), .DIN3(n2444), .DIN4(n2445), 
        .DIN5(n2446), .DIN6(n2447), .Q(n2416) );
  nor2s3 U1886 ( .DIN1(n2793), .DIN2(n2318), .Q(n2447) );
  nor2s3 U1887 ( .DIN1(n2792), .DIN2(n2359), .Q(n2446) );
  nor2s3 U1888 ( .DIN1(n2794), .DIN2(n2302), .Q(n2445) );
  nor2s3 U1889 ( .DIN1(n2797), .DIN2(n2351), .Q(n2444) );
  nor2s3 U1890 ( .DIN1(n2799), .DIN2(n876), .Q(n2443) );
  nor2s3 U1891 ( .DIN1(n2791), .DIN2(n2360), .Q(n2442) );
  nnd2s3 U1892 ( .DIN1(n2266), .DIN2(n569), .Q(g10379) );
  or5s3 U1893 ( .DIN1(n2448), .DIN2(n2449), .DIN3(n2450), .DIN4(n2451), .DIN5(
        n2452), .Q(n2824) );
  or5s3 U1894 ( .DIN1(n2453), .DIN2(n2454), .DIN3(n2455), .DIN4(n2456), .DIN5(
        n2457), .Q(n2452) );
  nor2s3 U1895 ( .DIN1(n2805), .DIN2(n876), .Q(n2457) );
  nor2s3 U1896 ( .DIN1(n2301), .DIN2(\DFF_319/net606 ), .Q(n2456) );
  nor2s3 U1897 ( .DIN1(n2801), .DIN2(n2359), .Q(n2455) );
  nor2s3 U1898 ( .DIN1(n2800), .DIN2(n2350), .Q(n2454) );
  and2s3 U1899 ( .DIN1(g4215), .DIN2(n2294), .Q(n2453) );
  nnd2s3 U1900 ( .DIN1(n2458), .DIN2(n2459), .Q(n2451) );
  nnd2s3 U1901 ( .DIN1(g4203), .DIN2(n2293), .Q(n2459) );
  or5s3 U1902 ( .DIN1(n886), .DIN2(n887), .DIN3(n2294), .DIN4(n894), .DIN5(
        n2460), .Q(n2458) );
  nnd4s2 U1903 ( .DIN1(n2440), .DIN2(g6262), .DIN3(g6261), .DIN4(n2461), .Q(
        n2311) );
  nor2s3 U1904 ( .DIN1(n2803), .DIN2(n2415), .Q(n2450) );
  nor2s3 U1905 ( .DIN1(n2802), .DIN2(n2352), .Q(n2449) );
  nor2s3 U1906 ( .DIN1(n2804), .DIN2(n2318), .Q(n2448) );
  nnd2s3 U1907 ( .DIN1(n2266), .DIN2(n577), .Q(g10377) );
  or5s3 U1908 ( .DIN1(n2462), .DIN2(n2463), .DIN3(n2464), .DIN4(n2465), .DIN5(
        n2466), .Q(g10774) );
  nnd4s2 U1909 ( .DIN1(n2467), .DIN2(n2468), .DIN3(n2469), .DIN4(n2470), .Q(
        n2466) );
  and4s2 U1910 ( .DIN1(n2471), .DIN2(n2472), .DIN3(n2473), .DIN4(n2474), .Q(
        n2470) );
  nnd2s3 U1911 ( .DIN1(n881), .DIN2(n578), .Q(n2474) );
  nnd2s3 U1912 ( .DIN1(n878), .DIN2(n2350), .Q(n2473) );
  or5s3 U1913 ( .DIN1(n885), .DIN2(n887), .DIN3(n888), .DIN4(n2294), .DIN5(
        n2460), .Q(n2300) );
  nnd4s2 U1914 ( .DIN1(n2301), .DIN2(n2475), .DIN3(n2476), .DIN4(n2477), .Q(
        n2460) );
  nor6s3 U1915 ( .DIN1(n2293), .DIN2(n881), .DIN3(n2411), .DIN4(n2340), .DIN5(
        n882), .DIN6(n2478), .Q(n2477) );
  nnd2s3 U1916 ( .DIN1(n2479), .DIN2(n2441), .Q(n2353) );
  nor5s3 U1917 ( .DIN1(g6259), .DIN2(n897), .DIN3(n900), .DIN4(n898), .DIN5(
        n2480), .Q(n2340) );
  and2s3 U1918 ( .DIN1(n2440), .DIN2(n893), .Q(n2411) );
  nnd2s3 U1919 ( .DIN1(n2441), .DIN2(n2481), .Q(n2352) );
  and3s3 U1920 ( .DIN1(n2415), .DIN2(n2336), .DIN3(n2341), .Q(n2476) );
  nnd3s3 U1921 ( .DIN1(n893), .DIN2(n898), .DIN3(n2482), .Q(n2341) );
  nnd2s3 U1922 ( .DIN1(g4214), .DIN2(n2294), .Q(n2472) );
  and2s3 U1923 ( .DIN1(n890), .DIN2(n2483), .Q(n2294) );
  nnd2s3 U1924 ( .DIN1(n888), .DIN2(n793), .Q(n2471) );
  nnd2s3 U1925 ( .DIN1(n890), .DIN2(n2479), .Q(n2425) );
  nnd2s3 U1926 ( .DIN1(n892), .DIN2(n667), .Q(n2469) );
  nnd2s3 U1927 ( .DIN1(n893), .DIN2(n2479), .Q(n2336) );
  and4s2 U1928 ( .DIN1(g6260), .DIN2(n897), .DIN3(n898), .DIN4(n899), .Q(n2479) );
  nnd2s3 U1929 ( .DIN1(n891), .DIN2(n690), .Q(n2468) );
  nnd2s3 U1930 ( .DIN1(n893), .DIN2(n2481), .Q(n2415) );
  nnd2s3 U1931 ( .DIN1(g4202), .DIN2(n2293), .Q(n2467) );
  and2s3 U1932 ( .DIN1(n2483), .DIN2(n893), .Q(n2293) );
  nnd3s3 U1933 ( .DIN1(n2461), .DIN2(n902), .DIN3(g6261), .Q(n2480) );
  nnd3s3 U1934 ( .DIN1(n2484), .DIN2(n2485), .DIN3(n2486), .Q(n2465) );
  nnd2s3 U1935 ( .DIN1(n887), .DIN2(n720), .Q(n2486) );
  nnd3s3 U1936 ( .DIN1(n890), .DIN2(g6258), .DIN3(n2482), .Q(n2359) );
  and3s3 U1937 ( .DIN1(g6260), .DIN2(g6257), .DIN3(g6259), .Q(n2482) );
  nnd2s3 U1938 ( .DIN1(n886), .DIN2(n798), .Q(n2485) );
  nnd2s3 U1939 ( .DIN1(n890), .DIN2(n2481), .Q(n2350) );
  and4s2 U1940 ( .DIN1(g6260), .DIN2(g6257), .DIN3(n898), .DIN4(n899), .Q(
        n2481) );
  nnd2s3 U1941 ( .DIN1(n885), .DIN2(n714), .Q(n2484) );
  or5s3 U1942 ( .DIN1(g6257), .DIN2(n900), .DIN3(n899), .DIN4(n898), .DIN5(
        n2487), .Q(n2360) );
  nnd3s3 U1943 ( .DIN1(n2461), .DIN2(n901), .DIN3(g6262), .Q(n2487) );
  nor2s3 U1944 ( .DIN1(n2812), .DIN2(n2301), .Q(n2464) );
  nor2s3 U1945 ( .DIN1(n2815), .DIN2(n2318), .Q(n2463) );
  nnd2s3 U1946 ( .DIN1(n2478), .DIN2(n2302), .Q(n2318) );
  nnd4s2 U1947 ( .DIN1(n2488), .DIN2(n2441), .DIN3(n897), .DIN4(n898), .Q(
        n2302) );
  and3s3 U1948 ( .DIN1(n2441), .DIN2(n898), .DIN3(n2488), .Q(n2478) );
  nor2s3 U1949 ( .DIN1(n2814), .DIN2(n876), .Q(n2462) );
  nor2s3 U1950 ( .DIN1(n2475), .DIN2(n879), .Q(n2299) );
  and2s3 U1951 ( .DIN1(n2351), .DIN2(n2489), .Q(n2475) );
  nnd2s3 U1952 ( .DIN1(n2483), .DIN2(n2441), .Q(n2489) );
  and3s3 U1953 ( .DIN1(n2488), .DIN2(g6257), .DIN3(g6258), .Q(n2483) );
  nnd2s3 U1954 ( .DIN1(n2440), .DIN2(n2441), .Q(n2351) );
  and3s3 U1955 ( .DIN1(n901), .DIN2(n902), .DIN3(n2461), .Q(n2441) );
  nor2s3 U1956 ( .DIN1(n908), .DIN2(n903), .Q(n2461) );
  or2s3 U1957 ( .DIN1(g6256), .DIN2(n2490), .Q(n908) );
  nor2s3 U1958 ( .DIN1(n2301), .DIN2(n2491), .Q(n2490) );
  nor2s3 U1959 ( .DIN1(g6263), .DIN2(g6254), .Q(n2491) );
  and3s3 U1960 ( .DIN1(n2488), .DIN2(n897), .DIN3(g6258), .Q(n2440) );
  nor2s3 U1961 ( .DIN1(n899), .DIN2(g6260), .Q(n2488) );
  nor2s3 U1962 ( .DIN1(n896), .DIN2(g6254), .Q(n2266) );
  nor2s3 U1963 ( .DIN1(n903), .DIN2(g6255), .Q(n2301) );
  i1s3 U1964 ( .DIN(n2510), .Q(n514) );
  i1s3 U1966 ( .DIN(n1363), .Q(n516) );
  i1s3 U1968 ( .DIN(n1838), .Q(n518) );
  i1s3 U1970 ( .DIN(n1872), .Q(n520) );
  i1s3 U1971 ( .DIN(n1846), .Q(n521) );
  i1s3 U1972 ( .DIN(n2819), .Q(n522) );
  i1s3 U1973 ( .DIN(n2818), .Q(n523) );
  i1s3 U1974 ( .DIN(n2776), .Q(n524) );
  i1s3 U1975 ( .DIN(n2631), .Q(n525) );
  i1s3 U1976 ( .DIN(n2820), .Q(n526) );
  i1s3 U1977 ( .DIN(n1747), .Q(n527) );
  i1s3 U1978 ( .DIN(n2583), .Q(n528) );
  i1s3 U1979 ( .DIN(n2719), .Q(n529) );
  i1s3 U1980 ( .DIN(n1357), .Q(n530) );
  i1s3 U1981 ( .DIN(n1248), .Q(n531) );
  i1s3 U1982 ( .DIN(n2621), .Q(n532) );
  i1s3 U1983 ( .DIN(n2634), .Q(n533) );
  i1s3 U1984 ( .DIN(n2498), .Q(n534) );
  i1s3 U1985 ( .DIN(n2821), .Q(n535) );
  i1s3 U1986 ( .DIN(n2542), .Q(n536) );
  i1s3 U1989 ( .DIN(n915), .Q(n539) );
  i1s3 U1991 ( .DIN(n1115), .Q(n541) );
  i1s3 U1992 ( .DIN(n1371), .Q(n542) );
  i1s3 U1993 ( .DIN(n1376), .Q(n543) );
  i1s3 U1995 ( .DIN(n1670), .Q(n545) );
  i1s3 U1996 ( .DIN(n2033), .Q(n546) );
  i1s3 U1997 ( .DIN(n2822), .Q(n547) );
  i1s3 U1998 ( .DIN(n2611), .Q(n548) );
  i1s3 U1999 ( .DIN(n2711), .Q(n549) );
  i1s3 U2000 ( .DIN(n2646), .Q(n550) );
  i1s3 U2001 ( .DIN(n2757), .Q(n551) );
  i1s3 U2002 ( .DIN(g4898), .Q(n552) );
  i1s3 U2003 ( .DIN(n2823), .Q(n553) );
  i1s3 U2004 ( .DIN(n2713), .Q(n554) );
  i1s3 U2005 ( .DIN(n2523), .Q(n555) );
  i1s3 U2006 ( .DIN(n2598), .Q(n556) );
  i1s3 U2007 ( .DIN(n2608), .Q(n557) );
  i1s3 U2008 ( .DIN(n2723), .Q(n558) );
  i1s3 U2009 ( .DIN(n2589), .Q(n559) );
  i1s3 U2010 ( .DIN(n2507), .Q(n560) );
  i1s3 U2011 ( .DIN(n2054), .Q(n561) );
  i1s3 U2012 ( .DIN(n2689), .Q(n562) );
  i1s3 U2013 ( .DIN(n2500), .Q(n563) );
  i1s3 U2014 ( .DIN(n1555), .Q(n564) );
  i1s3 U2015 ( .DIN(n906), .Q(n565) );
  i1s3 U2016 ( .DIN(n2031), .Q(n566) );
  i1s3 U2017 ( .DIN(n2670), .Q(n567) );
  i1s3 U2018 ( .DIN(n2129), .Q(n568) );
  i1s3 U2019 ( .DIN(n2824), .Q(n569) );
  i1s3 U2020 ( .DIN(n2605), .Q(n570) );
  i1s3 U2021 ( .DIN(n2825), .Q(n571) );
  i1s3 U2022 ( .DIN(n2728), .Q(n572) );
  i1s3 U2023 ( .DIN(n2032), .Q(n573) );
  i1s3 U2025 ( .DIN(n2536), .Q(n575) );
  i1s3 U2026 ( .DIN(n2643), .Q(n576) );
  i1s3 U2027 ( .DIN(g10774), .Q(n577) );
  i1s3 U2028 ( .DIN(n2806), .Q(n578) );
  i1s3 U2029 ( .DIN(n2700), .Q(n579) );
  i1s3 U2030 ( .DIN(n970), .Q(n580) );
  i1s3 U2031 ( .DIN(n1957), .Q(n581) );
  i1s3 U2032 ( .DIN(n2699), .Q(n582) );
  i1s3 U2033 ( .DIN(n2629), .Q(n583) );
  i1s3 U2034 ( .DIN(n2762), .Q(n584) );
  i1s3 U2035 ( .DIN(n2015), .Q(n585) );
  i1s3 U2038 ( .DIN(n1037), .Q(n588) );
  i1s3 U2039 ( .DIN(n1948), .Q(n589) );
  i1s3 U2040 ( .DIN(n1384), .Q(n590) );
  i1s3 U2041 ( .DIN(n927), .Q(n591) );
  i1s3 U2042 ( .DIN(n1062), .Q(n592) );
  i1s3 U2043 ( .DIN(n1063), .Q(n593) );
  i1s3 U2044 ( .DIN(n1956), .Q(n594) );
  i1s3 U2045 ( .DIN(n985), .Q(n595) );
  i1s3 U2046 ( .DIN(n986), .Q(n596) );
  i1s3 U2047 ( .DIN(n2773), .Q(n597) );
  i1s3 U2048 ( .DIN(n2053), .Q(n598) );
  i1s3 U2049 ( .DIN(n2615), .Q(n599) );
  i1s3 U2050 ( .DIN(n1840), .Q(n600) );
  i1s3 U2051 ( .DIN(n2597), .Q(n601) );
  i1s3 U2052 ( .DIN(n2581), .Q(n602) );
  i1s3 U2053 ( .DIN(n2535), .Q(n603) );
  i1s3 U2054 ( .DIN(n2715), .Q(n604) );
  i1s3 U2055 ( .DIN(n2658), .Q(n605) );
  i1s3 U2056 ( .DIN(n2730), .Q(n606) );
  i1s3 U2057 ( .DIN(n2599), .Q(n607) );
  i1s3 U2059 ( .DIN(n2641), .Q(n609) );
  i1s3 U2060 ( .DIN(n2494), .Q(n610) );
  i1s3 U2061 ( .DIN(n2740), .Q(n611) );
  i1s3 U2062 ( .DIN(n2784), .Q(n612) );
  i1s3 U2063 ( .DIN(n2560), .Q(n613) );
  i1s3 U2064 ( .DIN(n2722), .Q(n614) );
  i1s3 U2065 ( .DIN(n2644), .Q(n615) );
  i1s3 U2066 ( .DIN(n2642), .Q(n616) );
  i1s3 U2067 ( .DIN(n2691), .Q(n617) );
  i1s3 U2068 ( .DIN(n1340), .Q(n618) );
  i1s3 U2069 ( .DIN(n2603), .Q(n619) );
  i1s3 U2070 ( .DIN(n1929), .Q(n620) );
  i1s3 U2071 ( .DIN(n2816), .Q(n621) );
  i1s3 U2072 ( .DIN(n2656), .Q(n622) );
  i1s3 U2073 ( .DIN(n2747), .Q(n623) );
  i1s3 U2074 ( .DIN(n2671), .Q(n624) );
  i1s3 U2075 ( .DIN(n2051), .Q(n625) );
  i1s3 U2076 ( .DIN(n2676), .Q(n626) );
  i1s3 U2077 ( .DIN(n2659), .Q(n627) );
  i1s3 U2078 ( .DIN(n2717), .Q(n628) );
  i1s3 U2079 ( .DIN(n2515), .Q(n629) );
  i1s3 U2080 ( .DIN(n2568), .Q(n630) );
  i1s3 U2081 ( .DIN(n2052), .Q(n631) );
  i1s3 U2082 ( .DIN(n2014), .Q(n632) );
  i1s3 U2083 ( .DIN(n1561), .Q(n633) );
  i1s3 U2084 ( .DIN(n2687), .Q(n634) );
  i1s3 U2085 ( .DIN(n2050), .Q(n635) );
  i1s3 U2086 ( .DIN(n2744), .Q(n636) );
  i1s3 U2087 ( .DIN(n2016), .Q(n637) );
  i1s3 U2088 ( .DIN(n1936), .Q(n638) );
  i1s3 U2089 ( .DIN(n2017), .Q(n639) );
  i1s3 U2090 ( .DIN(n2636), .Q(n640) );
  i1s3 U2091 ( .DIN(n2680), .Q(n641) );
  i1s3 U2092 ( .DIN(n2572), .Q(n642) );
  i1s3 U2093 ( .DIN(n2703), .Q(n643) );
  i1s3 U2094 ( .DIN(n2504), .Q(n644) );
  i1s3 U2095 ( .DIN(n1400), .Q(n645) );
  i1s3 U2096 ( .DIN(n1398), .Q(n646) );
  i1s3 U2097 ( .DIN(n1596), .Q(n647) );
  i1s3 U2101 ( .DIN(n1026), .Q(n651) );
  i1s3 U2102 ( .DIN(n1980), .Q(n652) );
  i1s3 U2103 ( .DIN(n2678), .Q(n653) );
  i1s3 U2104 ( .DIN(n2661), .Q(n654) );
  i1s3 U2105 ( .DIN(n1479), .Q(n655) );
  i1s3 U2106 ( .DIN(n2817), .Q(n656) );
  i1s3 U2107 ( .DIN(n948), .Q(n657) );
  i1s3 U2108 ( .DIN(n960), .Q(n658) );
  i1s3 U2109 ( .DIN(n1103), .Q(n659) );
  i1s3 U2110 ( .DIN(n1978), .Q(n660) );
  i1s3 U2111 ( .DIN(n2009), .Q(n661) );
  i1s3 U2112 ( .DIN(n964), .Q(n662) );
  i1s3 U2113 ( .DIN(n1951), .Q(n663) );
  i1s3 U2114 ( .DIN(n2616), .Q(n664) );
  i1s3 U2115 ( .DIN(n2013), .Q(n665) );
  i1s3 U2116 ( .DIN(n1386), .Q(n666) );
  i1s3 U2117 ( .DIN(n2808), .Q(n667) );
  i1s3 U2118 ( .DIN(n2509), .Q(n668) );
  i1s3 U2119 ( .DIN(n2492), .Q(n669) );
  i1s3 U2120 ( .DIN(n2628), .Q(n670) );
  i1s3 U2121 ( .DIN(n2657), .Q(n671) );
  i1s3 U2122 ( .DIN(n2505), .Q(n672) );
  i1s3 U2123 ( .DIN(n1659), .Q(n673) );
  i1s3 U2124 ( .DIN(n2612), .Q(n674) );
  i1s3 U2125 ( .DIN(n1932), .Q(n675) );
  i1s3 U2126 ( .DIN(n1984), .Q(n676) );
  i1s3 U2127 ( .DIN(n1962), .Q(n677) );
  i1s3 U2128 ( .DIN(n2638), .Q(n678) );
  i1s3 U2129 ( .DIN(n1669), .Q(n679) );
  i1s3 U2130 ( .DIN(n2736), .Q(n680) );
  i1s3 U2131 ( .DIN(n2750), .Q(n681) );
  i1s3 U2132 ( .DIN(n1952), .Q(n682) );
  i1s3 U2134 ( .DIN(n2727), .Q(n684) );
  i1s3 U2135 ( .DIN(n2606), .Q(n685) );
  i1s3 U2136 ( .DIN(n2746), .Q(n686) );
  i1s3 U2137 ( .DIN(n1933), .Q(n687) );
  i1s3 U2138 ( .DIN(n2519), .Q(n688) );
  i1s3 U2139 ( .DIN(n2503), .Q(n689) );
  i1s3 U2140 ( .DIN(n2807), .Q(n690) );
  i1s3 U2141 ( .DIN(n1985), .Q(n691) );
  i1s3 U2142 ( .DIN(n2663), .Q(n692) );
  i1s3 U2143 ( .DIN(n2591), .Q(n693) );
  i1s3 U2144 ( .DIN(n2528), .Q(n694) );
  i1s3 U2145 ( .DIN(n1229), .Q(n695) );
  i1s3 U2146 ( .DIN(n2577), .Q(n696) );
  i1s3 U2147 ( .DIN(n1939), .Q(n697) );
  i1s3 U2148 ( .DIN(n1953), .Q(n698) );
  i1s3 U2149 ( .DIN(n2028), .Q(n699) );
  i1s3 U2150 ( .DIN(n1329), .Q(n700) );
  i1s3 U2151 ( .DIN(n2578), .Q(n701) );
  i1s3 U2152 ( .DIN(n1986), .Q(n702) );
  i1s3 U2153 ( .DIN(n2827), .Q(n703) );
  i1s3 U2154 ( .DIN(n2748), .Q(n704) );
  i1s3 U2155 ( .DIN(n2571), .Q(n705) );
  i1s3 U2156 ( .DIN(n1228), .Q(n706) );
  i1s3 U2157 ( .DIN(n2566), .Q(n707) );
  i1s3 U2158 ( .DIN(n2545), .Q(n708) );
  i1s3 U2159 ( .DIN(n2693), .Q(n709) );
  i1s3 U2160 ( .DIN(n1994), .Q(n710) );
  i1s3 U2161 ( .DIN(n2720), .Q(n711) );
  i1s3 U2162 ( .DIN(n1946), .Q(n712) );
  i1s3 U2163 ( .DIN(n2593), .Q(n713) );
  i1s3 U2164 ( .DIN(n2811), .Q(n714) );
  i1s3 U2165 ( .DIN(n2497), .Q(n715) );
  i1s3 U2166 ( .DIN(n2714), .Q(n716) );
  i1s3 U2167 ( .DIN(n1949), .Q(n717) );
  i1s3 U2169 ( .DIN(n2532), .Q(n719) );
  i1s3 U2170 ( .DIN(n2813), .Q(n720) );
  i1s3 U2171 ( .DIN(n2008), .Q(n721) );
  i1s3 U2172 ( .DIN(n2620), .Q(n722) );
  i1s3 U2173 ( .DIN(n2580), .Q(n723) );
  i1s3 U2174 ( .DIN(n2669), .Q(n724) );
  i1s3 U2175 ( .DIN(n1845), .Q(n725) );
  i1s3 U2176 ( .DIN(n2073), .Q(n726) );
  i1s3 U2177 ( .DIN(n2579), .Q(n727) );
  i1s3 U2178 ( .DIN(n1982), .Q(n728) );
  i1s3 U2179 ( .DIN(n2695), .Q(n729) );
  i1s3 U2180 ( .DIN(n2741), .Q(n730) );
  i1s3 U2181 ( .DIN(n1977), .Q(n731) );
  i1s3 U2182 ( .DIN(n2729), .Q(n732) );
  i1s3 U2183 ( .DIN(g1850), .Q(n733) );
  i1s3 U2184 ( .DIN(n2610), .Q(n734) );
  i1s3 U2185 ( .DIN(n2701), .Q(n735) );
  i1s3 U2186 ( .DIN(n2660), .Q(n736) );
  i1s3 U2187 ( .DIN(n2630), .Q(n737) );
  i1s3 U2189 ( .DIN(n2584), .Q(n739) );
  i1s3 U2190 ( .DIN(n2592), .Q(n740) );
  i1s3 U2191 ( .DIN(n2012), .Q(n741) );
  i1s3 U2192 ( .DIN(n2525), .Q(n742) );
  i1s3 U2193 ( .DIN(n2600), .Q(n743) );
  i1s3 U2194 ( .DIN(n2582), .Q(n744) );
  i1s3 U2195 ( .DIN(n2614), .Q(n745) );
  i1s3 U2196 ( .DIN(n2590), .Q(n746) );
  i1s3 U2197 ( .DIN(n1983), .Q(n747) );
  i1s3 U2198 ( .DIN(n2639), .Q(n748) );
  i1s3 U2199 ( .DIN(n2518), .Q(n749) );
  i1s3 U2200 ( .DIN(n2681), .Q(n750) );
  i1s3 U2201 ( .DIN(n2594), .Q(n751) );
  i1s3 U2202 ( .DIN(n1993), .Q(n752) );
  i1s3 U2203 ( .DIN(n2692), .Q(n753) );
  i1s3 U2204 ( .DIN(n2635), .Q(n754) );
  i1s3 U2205 ( .DIN(n2506), .Q(n755) );
  i1s3 U2206 ( .DIN(n2694), .Q(n756) );
  i1s3 U2207 ( .DIN(n2673), .Q(n757) );
  i1s3 U2208 ( .DIN(n2704), .Q(n758) );
  i1s3 U2209 ( .DIN(n2632), .Q(n759) );
  i1s3 U2210 ( .DIN(n2674), .Q(n760) );
  i1s3 U2211 ( .DIN(n2633), .Q(n761) );
  i1s3 U2212 ( .DIN(n2613), .Q(n762) );
  i1s3 U2213 ( .DIN(n2544), .Q(n763) );
  i1s3 U2214 ( .DIN(n2721), .Q(n764) );
  i1s3 U2215 ( .DIN(n2000), .Q(n765) );
  i1s3 U2216 ( .DIN(n2514), .Q(n766) );
  i1s3 U2217 ( .DIN(n2742), .Q(n767) );
  i1s3 U2218 ( .DIN(n1826), .Q(n768) );
  i1s3 U2219 ( .DIN(n2618), .Q(n769) );
  i1s3 U2220 ( .DIN(n1865), .Q(n770) );
  i1s3 U2221 ( .DIN(n2696), .Q(n771) );
  i1s3 U2222 ( .DIN(n1947), .Q(n772) );
  i1s3 U2223 ( .DIN(n2731), .Q(n773) );
  i1s3 U2224 ( .DIN(n2501), .Q(n774) );
  i1s3 U2225 ( .DIN(n2763), .Q(n775) );
  i1s3 U2226 ( .DIN(n1989), .Q(n776) );
  i1s3 U2227 ( .DIN(n2685), .Q(n777) );
  i1s3 U2228 ( .DIN(n2061), .Q(n778) );
  i1s3 U2229 ( .DIN(n2569), .Q(n779) );
  i1s3 U2230 ( .DIN(n2531), .Q(n780) );
  i1s3 U2231 ( .DIN(n2679), .Q(n781) );
  i1s3 U2232 ( .DIN(n2562), .Q(n782) );
  i1s3 U2233 ( .DIN(n2538), .Q(n783) );
  i1s3 U2234 ( .DIN(n2718), .Q(n784) );
  i1s3 U2235 ( .DIN(n2712), .Q(n785) );
  i1s3 U2236 ( .DIN(n2698), .Q(n786) );
  i1s3 U2237 ( .DIN(n1974), .Q(n787) );
  i1s3 U2238 ( .DIN(n2502), .Q(n788) );
  i1s3 U2239 ( .DIN(n1950), .Q(n789) );
  i1s3 U2240 ( .DIN(n2637), .Q(n790) );
  i1s3 U2241 ( .DIN(n2743), .Q(n791) );
  i1s3 U2242 ( .DIN(n1937), .Q(n792) );
  i1s3 U2243 ( .DIN(n2809), .Q(n793) );
  i1s3 U2244 ( .DIN(n1971), .Q(n794) );
  i1s3 U2245 ( .DIN(n2588), .Q(n795) );
  i1s3 U2246 ( .DIN(n2781), .Q(n796) );
  i1s3 U2247 ( .DIN(n1975), .Q(n797) );
  i1s3 U2248 ( .DIN(n2810), .Q(n798) );
  i1s3 U2249 ( .DIN(n2040), .Q(n799) );
  i1s3 U2250 ( .DIN(n2737), .Q(n800) );
  i1s3 U2251 ( .DIN(n2527), .Q(n801) );
  i1s3 U2252 ( .DIN(n2556), .Q(n802) );
  i1s3 U2253 ( .DIN(n1972), .Q(n803) );
  i1s3 U2254 ( .DIN(n2675), .Q(n804) );
  i1s3 U2255 ( .DIN(n2586), .Q(n805) );
  i1s3 U2256 ( .DIN(g632), .Q(n806) );
  i1s3 U2257 ( .DIN(n2683), .Q(n807) );
  i1s3 U2258 ( .DIN(n2574), .Q(n808) );
  i1s3 U2259 ( .DIN(n2624), .Q(n809) );
  i1s3 U2260 ( .DIN(n2540), .Q(n810) );
  i1s3 U2261 ( .DIN(n2041), .Q(n811) );
  i1s3 U2262 ( .DIN(n2623), .Q(n812) );
  i1s3 U2263 ( .DIN(n2619), .Q(n813) );
  i1s3 U2264 ( .DIN(n2520), .Q(n814) );
  i1s3 U2265 ( .DIN(n2706), .Q(n815) );
  i1s3 U2266 ( .DIN(n2530), .Q(n816) );
  i1s3 U2267 ( .DIN(g7329), .Q(n817) );
  i1s3 U2268 ( .DIN(n2567), .Q(n818) );
  i1s3 U2269 ( .DIN(n2587), .Q(n819) );
  i1s3 U2270 ( .DIN(n2493), .Q(n820) );
  i1s3 U2271 ( .DIN(n2508), .Q(n821) );
  i1s3 U2272 ( .DIN(n2563), .Q(n822) );
  i1s3 U2273 ( .DIN(n2739), .Q(n823) );
  i1s3 U2274 ( .DIN(n2596), .Q(n824) );
  i1s3 U2275 ( .DIN(n2734), .Q(n825) );
  i1s3 U2276 ( .DIN(n2576), .Q(n826) );
  i1s3 U2277 ( .DIN(n1963), .Q(n827) );
  i1s3 U2278 ( .DIN(n2025), .Q(n828) );
  i1s3 U2279 ( .DIN(n2702), .Q(n829) );
  i1s3 U2280 ( .DIN(n1981), .Q(n830) );
  i1s3 U2281 ( .DIN(n2595), .Q(n831) );
  i1s3 U2282 ( .DIN(n2708), .Q(n832) );
  i1s3 U2283 ( .DIN(n2516), .Q(n833) );
  i1s3 U2284 ( .DIN(n2609), .Q(n834) );
  i1s3 U2285 ( .DIN(n2499), .Q(n835) );
  i1s3 U2286 ( .DIN(n2622), .Q(n836) );
  i1s3 U2287 ( .DIN(n2604), .Q(n837) );
  i1s3 U2288 ( .DIN(n2029), .Q(n838) );
  i1s3 U2289 ( .DIN(n2564), .Q(n839) );
  i1s3 U2290 ( .DIN(n2662), .Q(n840) );
  i1s3 U2291 ( .DIN(n1280), .Q(n841) );
  i1s3 U2292 ( .DIN(n2760), .Q(n842) );
  i1s3 U2293 ( .DIN(n2640), .Q(n843) );
  i1s3 U2294 ( .DIN(n2697), .Q(n844) );
  i1s3 U2295 ( .DIN(n2495), .Q(n845) );
  i1s3 U2296 ( .DIN(n2524), .Q(n846) );
  i1s3 U2297 ( .DIN(n2735), .Q(n847) );
  i1s3 U2298 ( .DIN(n2716), .Q(n848) );
  i1s3 U2299 ( .DIN(n1954), .Q(n849) );
  i1s3 U2300 ( .DIN(n1987), .Q(n850) );
  i1s3 U2301 ( .DIN(n2522), .Q(n851) );
  i1s3 U2302 ( .DIN(n2543), .Q(n852) );
  i1s3 U2303 ( .DIN(n2002), .Q(n853) );
  i1s3 U2304 ( .DIN(n2607), .Q(n854) );
  i1s3 U2305 ( .DIN(n1976), .Q(n855) );
  i1s3 U2306 ( .DIN(n2048), .Q(n856) );
  i1s3 U2307 ( .DIN(n2570), .Q(n857) );
  i1s3 U2308 ( .DIN(n2710), .Q(n858) );
  i1s3 U2309 ( .DIN(n2539), .Q(n859) );
  i1s3 U2310 ( .DIN(n2645), .Q(n860) );
  i1s3 U2311 ( .DIN(n2738), .Q(n861) );
  i1s3 U2312 ( .DIN(n2625), .Q(n862) );
  i1s3 U2313 ( .DIN(n2565), .Q(n863) );
  i1s3 U2314 ( .DIN(n2496), .Q(n864) );
  i1s3 U2315 ( .DIN(n1930), .Q(n865) );
  i1s3 U2316 ( .DIN(n1958), .Q(n866) );
  i1s3 U2317 ( .DIN(n1955), .Q(n867) );
  i1s3 U2318 ( .DIN(n2001), .Q(n868) );
  i1s3 U2319 ( .DIN(n2789), .Q(n869) );
  i1s3 U2320 ( .DIN(n2677), .Q(n870) );
  i1s3 U2322 ( .DIN(g1696), .Q(n872) );
  i1s3 U2323 ( .DIN(g1700), .Q(n873) );
  i1s3 U2324 ( .DIN(g2355), .Q(n874) );
  i1s3 U2325 ( .DIN(g23), .Q(g3327) );
  i1s3 U2326 ( .DIN(n2299), .Q(n876) );
  i1s3 U2327 ( .DIN(n2405), .Q(n877) );
  i1s3 U2328 ( .DIN(n2300), .Q(n878) );
  i1s3 U2329 ( .DIN(n2351), .Q(n879) );
  i1s3 U2330 ( .DIN(n2318), .Q(n880) );
  i1s3 U2331 ( .DIN(n2352), .Q(n881) );
  i1s3 U2332 ( .DIN(n2353), .Q(n882) );
  i1s3 U2333 ( .DIN(n2312), .Q(n883) );
  i1s3 U2334 ( .DIN(n2313), .Q(n884) );
  i1s3 U2335 ( .DIN(n2360), .Q(n885) );
  i1s3 U2336 ( .DIN(n2350), .Q(n886) );
  i1s3 U2337 ( .DIN(n2359), .Q(n887) );
  i1s3 U2338 ( .DIN(n2425), .Q(n888) );
  i1s3 U2339 ( .DIN(n2433), .Q(n889) );
  i1s3 U2340 ( .DIN(n2487), .Q(n890) );
  i1s3 U2341 ( .DIN(n2415), .Q(n891) );
  i1s3 U2342 ( .DIN(n2336), .Q(n892) );
  i1s3 U2343 ( .DIN(n2480), .Q(n893) );
  i1s3 U2344 ( .DIN(n2311), .Q(n894) );
  i1s3 U2345 ( .DIN(n2147), .Q(n895) );
  i1s3 U2346 ( .DIN(n2301), .Q(n896) );
  i1s3 U2347 ( .DIN(g6257), .Q(n897) );
  i1s3 U2348 ( .DIN(g6258), .Q(n898) );
  i1s3 U2349 ( .DIN(g6259), .Q(n899) );
  i1s3 U2350 ( .DIN(g6260), .Q(n900) );
  i1s3 U2351 ( .DIN(g6261), .Q(n901) );
  i1s3 U2352 ( .DIN(g6262), .Q(n902) );
  i1s3 U2353 ( .DIN(g6263), .Q(n903) );
  i1s3 U2355 ( .DIN(g881), .Q(n905) );
  nnd5s3 U2356 ( .DIN1(n2550), .DIN2(n2549), .DIN3(n2554), .DIN4(n2559), 
        .DIN5(n2555), .Q(n1561) );
  nnd2s1 U2357 ( .DIN1(n2074), .DIN2(n785), .Q(n1235) );
  nnd2s1 U2358 ( .DIN1(n2074), .DIN2(n554), .Q(n1237) );
  nnd2s1 U2359 ( .DIN1(n2074), .DIN2(n716), .Q(n1239) );
  nnd2s2 U2360 ( .DIN1(n2074), .DIN2(n848), .Q(n1241) );
  nnd2s2 U2361 ( .DIN1(n2074), .DIN2(n711), .Q(n1243) );
  nnd2s2 U2362 ( .DIN1(n2074), .DIN2(n614), .Q(n1245) );
  nor6s1 U2363 ( .DIN1(n1631), .DIN2(n2628), .DIN3(n2074), .DIN4(n2623), 
        .DIN5(n2576), .DIN6(n2622), .Q(g6339) );
  nnd3s2 U2364 ( .DIN1(g1700), .DIN2(n826), .DIN3(n2074), .Q(n1595) );
  nnd2s2 U2365 ( .DIN1(n2074), .DIN2(n2628), .Q(n1899) );
  nnd3s2 U2366 ( .DIN1(n1887), .DIN2(n1888), .DIN3(n2074), .Q(n1879) );
  ib1s1 U2367 ( .DIN(n2074), .Q(n718) );
  ib1s9 U2368 ( .DIN(n2833), .Q(n2828) );
  ib1s9 U2369 ( .DIN(n2832), .Q(n2829) );
  ib1s9 U2370 ( .DIN(n2832), .Q(n2830) );
  ib1s9 U2371 ( .DIN(n2832), .Q(n2831) );
  ib1s9 U2372 ( .DIN(n2843), .Q(n2840) );
  ib1s9 U2373 ( .DIN(n2843), .Q(n2841) );
  ib1s9 U2374 ( .DIN(n2843), .Q(n2842) );
  ib1s9 U2375 ( .DIN(n2851), .Q(n2848) );
  ib1s9 U2376 ( .DIN(n2851), .Q(n2849) );
  ib1s9 U2377 ( .DIN(n2864), .Q(n2861) );
  ib1s9 U2378 ( .DIN(n2864), .Q(n2862) );
  ib1s9 U2379 ( .DIN(g109), .Q(n2865) );
  ib1s9 U2380 ( .DIN(g109), .Q(n2866) );
  ib1s9 U2381 ( .DIN(g109), .Q(n2867) );
  ib1s9 U2382 ( .DIN(g109), .Q(n2868) );
  ib1s9 U2383 ( .DIN(g109), .Q(n2869) );
  ib1s9 U2384 ( .DIN(g109), .Q(n2870) );
  ib1s9 U2385 ( .DIN(g6264), .Q(n904) );
  ib1s5 U2386 ( .DIN(n2203), .Q(n738) );
  ib1s5 U2387 ( .DIN(n1638), .Q(n683) );
  ib1s5 U2388 ( .DIN(n1601), .Q(n650) );
  ib1s5 U2389 ( .DIN(n1725), .Q(n649) );
  ib1s5 U2390 ( .DIN(n1432), .Q(n608) );
  ib1s5 U2391 ( .DIN(n1220), .Q(n587) );
  ib1s5 U2392 ( .DIN(n975), .Q(n586) );
  ib1s5 U2393 ( .DIN(n1435), .Q(n574) );
  ib1s5 U2394 ( .DIN(n1707), .Q(n544) );
  ib1s5 U2395 ( .DIN(n1112), .Q(n540) );
  ib1s5 U2396 ( .DIN(n1052), .Q(n538) );
  ib1s5 U2397 ( .DIN(n1192), .Q(n537) );
  ib1s5 U2398 ( .DIN(n1915), .Q(n517) );
  nnd4s3 U2399 ( .DIN1(n935), .DIN2(n927), .DIN3(n922), .DIN4(n580), .Q(n967)
         );
  i1s12 U2400 ( .DIN(n1701), .Q(n2832) );
  i1s12 U2401 ( .DIN(n1701), .Q(n2833) );
  i1s12 U2402 ( .DIN(n1701), .Q(n2834) );
  i1s12 U2403 ( .DIN(n1701), .Q(n2835) );
  i1s12 U2404 ( .DIN(n1701), .Q(n2836) );
  i1s12 U2405 ( .DIN(n1701), .Q(n2837) );
  i1s12 U2406 ( .DIN(n1701), .Q(n2838) );
  i1s12 U2407 ( .DIN(n1701), .Q(n2839) );
  i1s12 U2408 ( .DIN(n1487), .Q(n2843) );
  i1s12 U2409 ( .DIN(n1487), .Q(n2844) );
  i1s12 U2410 ( .DIN(n1487), .Q(n2845) );
  i1s12 U2411 ( .DIN(n1487), .Q(n2846) );
  i1s12 U2412 ( .DIN(n1487), .Q(n2847) );
  i1s12 U2413 ( .DIN(n2851), .Q(n2850) );
  i1s12 U2414 ( .DIN(n2860), .Q(n2851) );
  i1s12 U2415 ( .DIN(n2859), .Q(n2852) );
  i1s12 U2416 ( .DIN(n2859), .Q(n2853) );
  i1s12 U2417 ( .DIN(n2859), .Q(n2854) );
  i1s12 U2418 ( .DIN(n2858), .Q(n2855) );
  i1s12 U2419 ( .DIN(n2858), .Q(n2856) );
  i1s12 U2420 ( .DIN(n2858), .Q(n2857) );
  i1s12 U2421 ( .DIN(n1149), .Q(n2858) );
  i1s12 U2422 ( .DIN(n1149), .Q(n2859) );
  i1s12 U2423 ( .DIN(n1149), .Q(n2860) );
  i1s12 U2424 ( .DIN(n2864), .Q(n2863) );
  i1s12 U2425 ( .DIN(n874), .Q(n2864) );
  i1s12 U2426 ( .DIN(g109), .Q(n2871) );
  sdffs1 \DFF_533/Q_reg  ( .DIN(g7784), .SDIN(n3277), .SSEL(test_se), .CLK(CK), 
        .Q(g8984), .QN(n2034) );
  sdffs1 \DFF_532/Q_reg  ( .DIN(g8695), .SDIN(n3276), .SSEL(test_se), .CLK(CK), 
        .Q(n3277), .QN(n2510) );
  sdffs1 \DFF_531/Q_reg  ( .DIN(g7337), .SDIN(n3275), .SSEL(test_se), .CLK(CK), 
        .Q(n3276), .QN(n2776) );
  sdffs1 \DFF_530/Q_reg  ( .DIN(g10879), .SDIN(n3274), .SSEL(test_se), .CLK(CK), .Q(n3275), .QN(n2778) );
  sdffs1 \DFF_529/Q_reg  ( .DIN(g11336), .SDIN(n3273), .SSEL(test_se), .CLK(CK), .Q(n3274), .QN(n2631) );
  sdffs1 \DFF_528/Q_reg  ( .DIN(g8078), .SDIN(g1360), .SSEL(test_se), .CLK(CK), 
        .Q(n3273), .QN(n2764) );
  sdffs1 \DFF_526/Q_reg  ( .DIN(g9824), .SDIN(n2583), .SSEL(test_se), .CLK(CK), 
        .Q(g1360) );
  sdffs1 \DFF_525/Q_reg  ( .DIN(g6302), .SDIN(n3272), .SSEL(test_se), .CLK(CK), 
        .Q(n2583) );
  sdffs1 \DFF_524/Q_reg  ( .DIN(g10876), .SDIN(n3271), .SSEL(test_se), .CLK(CK), .Q(n3272), .QN(n2719) );
  sdffs1 \DFF_523/Q_reg  ( .DIN(g7812), .SDIN(n3270), .SSEL(test_se), .CLK(CK), 
        .Q(n3271), .QN(n2621) );
  sdffs1 \DFF_522/Q_reg  ( .DIN(g11327), .SDIN(n3269), .SSEL(test_se), .CLK(CK), .Q(n3270), .QN(n2634) );
  sdffs1 \DFF_521/Q_reg  ( .DIN(g8430), .SDIN(n3268), .SSEL(test_se), .CLK(CK), 
        .Q(n3269), .QN(n2498) );
  sdffs1 \DFF_520/Q_reg  ( .DIN(g7352), .SDIN(n3267), .SSEL(test_se), .CLK(CK), 
        .Q(n3268), .QN(n2795) );
  sdffs1 \DFF_519/Q_reg  ( .DIN(g8446), .SDIN(n3266), .SSEL(test_se), .CLK(CK), 
        .Q(n3267), .QN(n2542) );
  sdffs1 \DFF_518/Q_reg  ( .DIN(g8064), .SDIN(n2585), .SSEL(test_se), .CLK(CK), 
        .Q(n3266), .QN(n2517) );
  sdffs1 \DFF_517/Q_reg  ( .DIN(g6313), .SDIN(n3265), .SSEL(test_se), .CLK(CK), 
        .Q(n2585) );
  sdffs1 \DFF_516/Q_reg  ( .DIN(g8869), .SDIN(n3264), .SSEL(test_se), .CLK(CK), 
        .Q(n3265), .QN(n2705) );
  sdffs1 \DFF_515/Q_reg  ( .DIN(g7801), .SDIN(n3263), .SSEL(test_se), .CLK(CK), 
        .Q(n3264), .QN(n2654) );
  sdffs1 \DFF_514/Q_reg  ( .DIN(g7348), .SDIN(g8981), .SSEL(test_se), .CLK(CK), 
        .Q(n3263), .QN(n2772) );
  sdffs1 \DFF_513/Q_reg  ( .DIN(g7781), .SDIN(n3262), .SSEL(test_se), .CLK(CK), 
        .Q(g8981), .QN(n2019) );
  sdffs1 \DFF_512/Q_reg  ( .DIN(g11261), .SDIN(n3261), .SSEL(test_se), .CLK(CK), .Q(n3262), .QN(n2033) );
  sdffs1 \DFF_511/Q_reg  ( .DIN(g7772), .SDIN(n3260), .SSEL(test_se), .CLK(CK), 
        .Q(n3261), .QN(n2745) );
  sdffs1 \DFF_510/Q_reg  ( .DIN(g7296), .SDIN(n3259), .SSEL(test_se), .CLK(CK), 
        .Q(n3260), .QN(n2611) );
  sdffs1 \DFF_509/Q_reg  ( .DIN(g11611), .SDIN(n3258), .SSEL(test_se), .CLK(CK), .Q(n3259), .QN(n2711) );
  sdffs1 \DFF_508/Q_reg  ( .DIN(g8421), .SDIN(n2646), .SSEL(test_se), .CLK(CK), 
        .Q(n3258), .QN(n1960) );
  sdffs1 \DFF_507/Q_reg  ( .DIN(g11181), .SDIN(n3257), .SSEL(test_se), .CLK(CK), .Q(n2646) );
  sdffs1 \DFF_506/Q_reg  ( .DIN(g11657), .SDIN(n3256), .SSEL(test_se), .CLK(CK), .Q(n3257), .QN(n2757) );
  sdffs1 \DFF_505/Q_reg  ( .DIN(g7339), .SDIN(n3255), .SSEL(test_se), .CLK(CK), 
        .Q(n3256), .QN(n2785) );
  sdffs1 \DFF_504/Q_reg  ( .DIN(g11035), .SDIN(n3254), .SSEL(test_se), .CLK(CK), .Q(n3255), .QN(n2713) );
  sdffs1 \DFF_503/Q_reg  ( .DIN(g8988), .SDIN(g2611), .SSEL(test_se), .CLK(CK), 
        .Q(n3254), .QN(n2523) );
  sdffs1 \DFF_502/Q_reg  ( .DIN(g6282), .SDIN(n3253), .SSEL(test_se), .CLK(CK), 
        .Q(g2611) );
  sdffs1 \DFF_501/Q_reg  ( .DIN(g5665), .SDIN(g5645), .SSEL(test_se), .CLK(CK), 
        .Q(n3253), .QN(n2765) );
  sdffs1 \DFF_500/Q_reg  ( .DIN(g7752), .SDIN(n3252), .SSEL(test_se), .CLK(CK), 
        .Q(g5645) );
  sdffs1 \DFF_499/Q_reg  ( .DIN(g11505), .SDIN(n3251), .SSEL(test_se), .CLK(CK), .Q(n3252), .QN(n2598) );
  sdffs1 \DFF_498/Q_reg  ( .DIN(g7291), .SDIN(n3250), .SSEL(test_se), .CLK(CK), 
        .Q(n3251), .QN(n2608) );
  sdffs1 \DFF_497/Q_reg  ( .DIN(g7802), .SDIN(g8976), .SSEL(test_se), .CLK(CK), 
        .Q(n3250), .QN(n2648) );
  sdffs1 \DFF_496/Q_reg  ( .DIN(g7774), .SDIN(n3249), .SSEL(test_se), .CLK(CK), 
        .Q(g8976), .QN(n2038) );
  sdffs1 \DFF_495/Q_reg  ( .DIN(g8872), .SDIN(n3248), .SSEL(test_se), .CLK(CK), 
        .Q(n3249), .QN(n2723) );
  sdffs1 \DFF_494/Q_reg  ( .DIN(g7333), .SDIN(n3247), .SSEL(test_se), .CLK(CK), 
        .Q(n3248), .QN(n2589) );
  sdffs1 \DFF_493/Q_reg  ( .DIN(g8283), .SDIN(n3246), .SSEL(test_se), .CLK(CK), 
        .Q(n3247), .QN(n2507) );
  sdffs1 \DFF_492/Q_reg  ( .DIN(g11262), .SDIN(n3245), .SSEL(test_se), .CLK(CK), .Q(n3246), .QN(n2054) );
  sdffs1 \DFF_491/Q_reg  ( .DIN(g11268), .SDIN(n3244), .SSEL(test_se), .CLK(CK), .Q(n3245), .QN(n2689) );
  sdffs1 \DFF_490/Q_reg  ( .DIN(g8424), .SDIN(n3243), .SSEL(test_se), .CLK(CK), 
        .Q(n3244), .QN(n1959) );
  sdffs1 \DFF_489/Q_reg  ( .DIN(g5672), .SDIN(n3242), .SSEL(test_se), .CLK(CK), 
        .Q(n3243), .QN(\DFF_489/net776 ) );
  sdffs1 \DFF_488/Q_reg  ( .DIN(g8428), .SDIN(n2553), .SSEL(test_se), .CLK(CK), 
        .Q(n3242), .QN(n2500) );
  sdffs1 \DFF_487/Q_reg  ( .DIN(g7314), .SDIN(n3241), .SSEL(test_se), .CLK(CK), 
        .Q(n2553) );
  sdffs1 \DFF_486/Q_reg  ( .DIN(g7294), .SDIN(n3240), .SSEL(test_se), .CLK(CK), 
        .Q(n3241), .QN(n2031) );
  sdffs1 \DFF_485/Q_reg  ( .DIN(g7761), .SDIN(n2561), .SSEL(test_se), .CLK(CK), 
        .Q(n3240), .QN(n2779) );
  sdffs1 \DFF_484/Q_reg  ( .DIN(g6825), .SDIN(n3239), .SSEL(test_se), .CLK(CK), 
        .Q(n2561) );
  sdffs1 \DFF_483/Q_reg  ( .DIN(g11442), .SDIN(n3238), .SSEL(test_se), .CLK(CK), .Q(n3239), .QN(n2670) );
  sdffs1 \DFF_482/Q_reg  ( .DIN(g8868), .SDIN(n3237), .SSEL(test_se), .CLK(CK), 
        .Q(n3238), .QN(n2707) );
  sdffs1 \DFF_481/Q_reg  ( .DIN(g11628), .SDIN(n3236), .SSEL(test_se), .CLK(CK), .Q(n3237), .QN(n2800) );
  sdffs1 \DFF_480/Q_reg  ( .DIN(g11443), .SDIN(g8982), .SSEL(test_se), .CLK(CK), .Q(n3236), .QN(n2605) );
  sdffs1 \DFF_479/Q_reg  ( .DIN(g7782), .SDIN(n3235), .SSEL(test_se), .CLK(CK), 
        .Q(g8982), .QN(n2035) );
  sdffs1 \DFF_478/Q_reg  ( .DIN(g5647), .SDIN(n3234), .SSEL(test_se), .CLK(CK), 
        .Q(n3235), .QN(n2686) );
  sdffs1 \DFF_477/Q_reg  ( .DIN(g7365), .SDIN(g2607), .SSEL(test_se), .CLK(CK), 
        .Q(n3234), .QN(n2728) );
  sdffs1 \DFF_476/Q_reg  ( .DIN(g6284), .SDIN(n3233), .SSEL(test_se), .CLK(CK), 
        .Q(g2607) );
  sdffs1 \DFF_475/Q_reg  ( .DIN(g11329), .SDIN(n3232), .SSEL(test_se), .CLK(CK), .Q(n3233), .QN(n2032) );
  sdffs1 \DFF_474/Q_reg  ( .DIN(g8419), .SDIN(n2536), .SSEL(test_se), .CLK(CK), 
        .Q(n3232), .QN(n1961) );
  sdffs1 \DFF_473/Q_reg  ( .DIN(g7321), .SDIN(n2643), .SSEL(test_se), .CLK(CK), 
        .Q(n2536) );
  sdffs1 \DFF_472/Q_reg  ( .DIN(g11184), .SDIN(g1710), .SSEL(test_se), .CLK(CK), .Q(n2643) );
  sdffs1 \DFF_471/Q_reg  ( .DIN(g4901), .SDIN(n3231), .SSEL(test_se), .CLK(CK), 
        .Q(g1710) );
  sdffs1 \DFF_470/Q_reg  ( .DIN(g11655), .SDIN(n3230), .SSEL(test_se), .CLK(CK), .Q(n3231), .QN(n2782) );
  sdffs1 \DFF_468/Q_reg  ( .DIN(g6311), .SDIN(n3229), .SSEL(test_se), .CLK(CK), 
        .Q(n3230), .QN(n1944) );
  sdffs1 \DFF_467/Q_reg  ( .DIN(g5648), .SDIN(n3228), .SSEL(test_se), .CLK(CK), 
        .Q(n3229), .QN(n2682) );
  sdffs1 \DFF_466/Q_reg  ( .DIN(g7358), .SDIN(n3227), .SSEL(test_se), .CLK(CK), 
        .Q(n3228), .QN(n2806) );
  sdffs1 \DFF_465/Q_reg  ( .DIN(g11042), .SDIN(g2610), .SSEL(test_se), .CLK(CK), .Q(n3227), .QN(n2700) );
  sdffs1 \DFF_464/Q_reg  ( .DIN(g6281), .SDIN(n3226), .SSEL(test_se), .CLK(CK), 
        .Q(g2610) );
  sdffs1 \DFF_463/Q_reg  ( .DIN(g7347), .SDIN(g755), .SSEL(test_se), .CLK(CK), 
        .Q(n3226), .QN(n2783) );
  sdffs1 \DFF_462/Q_reg  ( .DIN(g6265), .SDIN(n3225), .SSEL(test_se), .CLK(CK), 
        .Q(g755) );
  sdffs1 \DFF_461/Q_reg  ( .DIN(g9352), .SDIN(n3224), .SSEL(test_se), .CLK(CK), 
        .Q(n3225), .QN(n1957) );
  sdffs1 \DFF_460/Q_reg  ( .DIN(g11043), .SDIN(n3223), .SSEL(test_se), .CLK(CK), .Q(n3224), .QN(n2699) );
  sdffs1 \DFF_459/Q_reg  ( .DIN(g11335), .SDIN(n3222), .SSEL(test_se), .CLK(CK), .Q(n3223), .QN(n2629) );
  sdffs1 \DFF_458/Q_reg  ( .DIN(g11631), .SDIN(n3221), .SSEL(test_se), .CLK(CK), .Q(n3222), .QN(n2762) );
  sdffs1 \DFF_457/Q_reg  ( .DIN(g6306), .SDIN(n3220), .SSEL(test_se), .CLK(CK), 
        .Q(n3221), .QN(n2015) );
  sdffs1 \DFF_456/Q_reg  ( .DIN(g7362), .SDIN(n3219), .SSEL(test_se), .CLK(CK), 
        .Q(n3220), .QN(n2769) );
  sdffs1 \DFF_455/Q_reg  ( .DIN(g9895), .SDIN(n3218), .SSEL(test_se), .CLK(CK), 
        .Q(n3219), .QN(n1948) );
  sdffs1 \DFF_454/Q_reg  ( .DIN(g11399), .SDIN(n3217), .SSEL(test_se), .CLK(CK), .Q(n3218), .QN(n2803) );
  sdffs1 \DFF_453/Q_reg  ( .DIN(g7346), .SDIN(n3216), .SSEL(test_se), .CLK(CK), 
        .Q(n3217), .QN(n2797) );
  sdffs1 \DFF_452/Q_reg  ( .DIN(n565), .SDIN(g2608), .SSEL(test_se), .CLK(CK), 
        .Q(n3216), .QN(\DFF_452/net739 ) );
  sdffs1 \DFF_451/Q_reg  ( .DIN(g6285), .SDIN(n3215), .SSEL(test_se), .CLK(CK), 
        .Q(g2608) );
  sdffs1 \DFF_450/Q_reg  ( .DIN(g9341), .SDIN(n3214), .SSEL(test_se), .CLK(CK), 
        .Q(n3215), .QN(n1968) );
  sdffs1 \DFF_449/Q_reg  ( .DIN(g9348), .SDIN(n3213), .SSEL(test_se), .CLK(CK), 
        .Q(n3214), .QN(n1956) );
  sdffs1 \DFF_448/Q_reg  ( .DIN(g11630), .SDIN(n3212), .SSEL(test_se), .CLK(CK), .Q(n3213), .QN(n2773) );
  sdffs1 \DFF_447/Q_reg  ( .DIN(g11330), .SDIN(g5647), .SSEL(test_se), .CLK(CK), .Q(n3212), .QN(n2053) );
  sdffs1 \DFF_446/Q_reg  ( .DIN(g7754), .SDIN(g7), .SSEL(test_se), .CLK(CK), 
        .Q(g5647) );
  sdffs1 \DFF_445/Q_reg  ( .DIN(g2731), .SDIN(n3211), .SSEL(test_se), .CLK(CK), 
        .Q(g7) );
  sdffs1 \DFF_444/Q_reg  ( .DIN(g8420), .SDIN(g5649), .SSEL(test_se), .CLK(CK), 
        .Q(n3211), .QN(n1996) );
  sdffs1 \DFF_443/Q_reg  ( .DIN(g7756), .SDIN(n3210), .SSEL(test_se), .CLK(CK), 
        .Q(g5649) );
  sdffs1 \DFF_442/Q_reg  ( .DIN(g7301), .SDIN(n3209), .SSEL(test_se), .CLK(CK), 
        .Q(n3210), .QN(n2615) );
  sdffs1 \DFF_441/Q_reg  ( .DIN(g874), .SDIN(n3208), .SSEL(test_se), .CLK(CK), 
        .Q(n3209), .QN(\DFF_441/net728 ) );
  sdffs1 \DFF_440/Q_reg  ( .DIN(g11506), .SDIN(n2581), .SSEL(test_se), .CLK(CK), .Q(n3208), .QN(n2597) );
  sdffs1 \DFF_438/Q_reg  ( .DIN(g6300), .SDIN(n3207), .SSEL(test_se), .CLK(CK), 
        .Q(n2581) );
  sdffs1 \DFF_437/Q_reg  ( .DIN(g8445), .SDIN(n3206), .SSEL(test_se), .CLK(CK), 
        .Q(n3207), .QN(n2535) );
  sdffs1 \DFF_436/Q_reg  ( .DIN(g113), .SDIN(n3205), .SSEL(test_se), .CLK(CK), 
        .Q(n3206), .QN(\DFF_436/net723 ) );
  sdffs1 \DFF_435/Q_reg  ( .DIN(g8449), .SDIN(g4181), .SSEL(test_se), .CLK(CK), 
        .Q(n3205), .QN(n2715) );
  sdffs1 \DFF_434/Q_reg  ( .DIN(g8567), .SDIN(n3204), .SSEL(test_se), .CLK(CK), 
        .Q(g4181), .QN(n2055) );
  sdffs1 \DFF_433/Q_reg  ( .DIN(g4186), .SDIN(n3203), .SSEL(test_se), .CLK(CK), 
        .Q(n3204), .QN(n2658) );
  sdffs1 \DFF_432/Q_reg  ( .DIN(g11634), .SDIN(g4172), .SSEL(test_se), .CLK(CK), .Q(n3203), .QN(n2730) );
  sdffs1 \DFF_431/Q_reg  ( .DIN(g4895), .SDIN(n3202), .SSEL(test_se), .CLK(CK), 
        .Q(g4172), .QN(n2599) );
  sdffs1 \DFF_430/Q_reg  ( .DIN(g11324), .SDIN(g4183), .SSEL(test_se), .CLK(CK), .Q(n3202), .QN(n2641) );
  sdffs1 \DFF_429/Q_reg  ( .DIN(g6801), .SDIN(n3201), .SSEL(test_se), .CLK(CK), 
        .Q(g4183), .QN(n1990) );
  sdffs1 \DFF_428/Q_reg  ( .DIN(g7804), .SDIN(n3200), .SSEL(test_se), .CLK(CK), 
        .Q(n3201), .QN(n2655) );
  sdffs1 \DFF_427/Q_reg  ( .DIN(g8434), .SDIN(n3199), .SSEL(test_se), .CLK(CK), 
        .Q(n3200), .QN(n2494) );
  sdffs1 \DFF_426/Q_reg  ( .DIN(g7342), .SDIN(n3198), .SSEL(test_se), .CLK(CK), 
        .Q(n3199), .QN(n2740) );
  sdffs1 \DFF_425/Q_reg  ( .DIN(g7361), .SDIN(n2560), .SSEL(test_se), .CLK(CK), 
        .Q(n3198), .QN(n2784) );
  sdffs1 \DFF_424/Q_reg  ( .DIN(g6835), .SDIN(n3197), .SSEL(test_se), .CLK(CK), 
        .Q(n2560) );
  sdffs1 \DFF_423/Q_reg  ( .DIN(g10874), .SDIN(n2644), .SSEL(test_se), .CLK(CK), .Q(n3197), .QN(n2722) );
  sdffs1 \DFF_421/Q_reg  ( .DIN(g11183), .SDIN(n3196), .SSEL(test_se), .CLK(CK), .Q(n2644) );
  sdffs1 \DFF_420/Q_reg  ( .DIN(g11185), .SDIN(n3195), .SSEL(test_se), .CLK(CK), .Q(n3196), .QN(n2642) );
  sdffs1 \DFF_419/Q_reg  ( .DIN(g11267), .SDIN(n3194), .SSEL(test_se), .CLK(CK), .Q(n3195), .QN(n2691) );
  sdffs1 \DFF_418/Q_reg  ( .DIN(g8277), .SDIN(n3193), .SSEL(test_se), .CLK(CK), 
        .Q(n3194), .QN(n2603) );
  sdffs1 \DFF_417/Q_reg  ( .DIN(g6816), .SDIN(n3192), .SSEL(test_se), .CLK(CK), 
        .Q(n3193), .QN(n1929) );
  sdffs1 \DFF_416/Q_reg  ( .DIN(g6312), .SDIN(n3191), .SSEL(test_se), .CLK(CK), 
        .Q(n3192), .QN(n1970) );
  sdffs1 \DFF_415/Q_reg  ( .DIN(g8991), .SDIN(n3190), .SSEL(test_se), .CLK(CK), 
        .Q(n3191), .QN(n2526) );
  sdffs1 \DFF_414/Q_reg  ( .DIN(g7803), .SDIN(n3189), .SSEL(test_se), .CLK(CK), 
        .Q(n3190), .QN(n2649) );
  sdffs1 \DFF_413/Q_reg  ( .DIN(g7798), .SDIN(n3188), .SSEL(test_se), .CLK(CK), 
        .Q(n3189), .QN(n2816) );
  sdffs1 \DFF_412/Q_reg  ( .DIN(g4185), .SDIN(g2604), .SSEL(test_se), .CLK(CK), 
        .Q(n3188), .QN(n2656) );
  sdffs1 \DFF_411/Q_reg  ( .DIN(g6253), .SDIN(n3187), .SSEL(test_se), .CLK(CK), 
        .Q(g2604) );
  sdffs1 \DFF_410/Q_reg  ( .DIN(g5667), .SDIN(n3186), .SSEL(test_se), .CLK(CK), 
        .Q(n3187), .QN(n2747) );
  sdffs1 \DFF_409/Q_reg  ( .DIN(g11441), .SDIN(n3185), .SSEL(test_se), .CLK(CK), .Q(n3186), .QN(n2671) );
  sdffs1 \DFF_408/Q_reg  ( .DIN(g11402), .SDIN(g4174), .SSEL(test_se), .CLK(CK), .Q(n3185), .QN(n2761) );
  sdffs1 \DFF_407/Q_reg  ( .DIN(g6798), .SDIN(n3184), .SSEL(test_se), .CLK(CK), 
        .Q(g4174), .QN(n2051) );
  sdffs1 \DFF_406/Q_reg  ( .DIN(g11270), .SDIN(n3183), .SSEL(test_se), .CLK(CK), .Q(n3184), .QN(n2676) );
  sdffs1 \DFF_405/Q_reg  ( .DIN(g4188), .SDIN(n3182), .SSEL(test_se), .CLK(CK), 
        .Q(n3183), .QN(n2659) );
  sdffs1 \DFF_404/Q_reg  ( .DIN(g8874), .SDIN(n2515), .SSEL(test_se), .CLK(CK), 
        .Q(n3182), .QN(n2717) );
  sdffs1 \DFF_403/Q_reg  ( .DIN(g8066), .SDIN(n3181), .SSEL(test_se), .CLK(CK), 
        .Q(n2515) );
  sdffs1 \DFF_402/Q_reg  ( .DIN(g6807), .SDIN(n3180), .SSEL(test_se), .CLK(CK), 
        .Q(n3181), .QN(n2568) );
  sdffs1 \DFF_401/Q_reg  ( .DIN(g7295), .SDIN(n3179), .SSEL(test_se), .CLK(CK), 
        .Q(n3180), .QN(n2052) );
  sdffs1 \DFF_400/Q_reg  ( .DIN(g7304), .SDIN(n3178), .SSEL(test_se), .CLK(CK), 
        .Q(n3179), .QN(n1995) );
  sdffs1 \DFF_399/Q_reg  ( .DIN(g6307), .SDIN(g875), .SSEL(test_se), .CLK(CK), 
        .Q(n3178), .QN(n2014) );
  sdffs1 \DFF_398/Q_reg  ( .DIN(g9822), .SDIN(g5643), .SSEL(test_se), .CLK(CK), 
        .Q(g875) );
  sdffs1 \DFF_397/Q_reg  ( .DIN(g7750), .SDIN(n3177), .SSEL(test_se), .CLK(CK), 
        .Q(g5643) );
  sdffs1 \DFF_396/Q_reg  ( .DIN(g7318), .SDIN(n3176), .SSEL(test_se), .CLK(CK), 
        .Q(n3177), .QN(n2554) );
  sdffs1 \DFF_395/Q_reg  ( .DIN(g9339), .SDIN(n3175), .SSEL(test_se), .CLK(CK), 
        .Q(n3176), .QN(n2039) );
  sdffs1 \DFF_394/Q_reg  ( .DIN(g11264), .SDIN(g4186), .SSEL(test_se), .CLK(CK), .Q(n3175), .QN(n2687) );
  sdffs1 \DFF_393/Q_reg  ( .DIN(g7786), .SDIN(n3174), .SSEL(test_se), .CLK(CK), 
        .Q(g4186), .QN(n2050) );
  sdffs1 \DFF_392/Q_reg  ( .DIN(g7355), .SDIN(n3173), .SSEL(test_se), .CLK(CK), 
        .Q(n3174), .QN(n2756) );
  sdffs1 \DFF_391/Q_reg  ( .DIN(g7338), .SDIN(n3172), .SSEL(test_se), .CLK(CK), 
        .Q(n3173), .QN(n2799) );
  sdffs1 \DFF_390/Q_reg  ( .DIN(g7764), .SDIN(g4184), .SSEL(test_se), .CLK(CK), 
        .Q(n3172), .QN(n2744) );
  sdffs1 \DFF_389/Q_reg  ( .DIN(g6802), .SDIN(n3171), .SSEL(test_se), .CLK(CK), 
        .Q(g4184), .QN(n1999) );
  sdffs1 \DFF_388/Q_reg  ( .DIN(g5664), .SDIN(g4188), .SSEL(test_se), .CLK(CK), 
        .Q(n3171), .QN(n2777) );
  sdffs1 \DFF_387/Q_reg  ( .DIN(g8274), .SDIN(n3170), .SSEL(test_se), .CLK(CK), 
        .Q(g4188), .QN(n2049) );
  sdffs1 \DFF_386/Q_reg  ( .DIN(g7760), .SDIN(n3169), .SSEL(test_se), .CLK(CK), 
        .Q(n3170), .QN(n2793) );
  sdffs1 \DFF_385/Q_reg  ( .DIN(g7366), .SDIN(n3168), .SSEL(test_se), .CLK(CK), 
        .Q(n3169), .QN(\DFF_385/net672 ) );
  sdffs1 \DFF_384/Q_reg  ( .DIN(n2818), .SDIN(n3167), .SSEL(test_se), .CLK(CK), 
        .Q(n3168), .QN(\DFF_384/net671 ) );
  sdffs1 \DFF_383/Q_reg  ( .DIN(g6305), .SDIN(n3166), .SSEL(test_se), .CLK(CK), 
        .Q(n3167), .QN(n2016) );
  sdffs1 \DFF_382/Q_reg  ( .DIN(g8418), .SDIN(n3165), .SSEL(test_se), .CLK(CK), 
        .Q(n3166), .QN(n1938) );
  sdffs1 \DFF_381/Q_reg  ( .DIN(g9340), .SDIN(n3164), .SSEL(test_se), .CLK(CK), 
        .Q(n3165), .QN(n1936) );
  sdffs1 \DFF_380/Q_reg  ( .DIN(g7745), .SDIN(n3163), .SSEL(test_se), .CLK(CK), 
        .Q(n3164), .QN(n2017) );
  sdffs1 \DFF_379/Q_reg  ( .DIN(g11338), .SDIN(n3162), .SSEL(test_se), .CLK(CK), .Q(n3163), .QN(n2636) );
  sdffs1 \DFF_378/Q_reg  ( .DIN(g11260), .SDIN(g2601), .SSEL(test_se), .CLK(CK), .Q(n3162), .QN(n2680) );
  sdffs1 \DFF_377/Q_reg  ( .DIN(g6281), .SDIN(n3161), .SSEL(test_se), .CLK(CK), 
        .Q(g2601) );
  sdffs1 \DFF_376/Q_reg  ( .DIN(g6803), .SDIN(n3160), .SSEL(test_se), .CLK(CK), 
        .Q(n3161), .QN(n2572) );
  sdffs1 \DFF_374/Q_reg  ( .DIN(g8870), .SDIN(n3159), .SSEL(test_se), .CLK(CK), 
        .Q(n3160), .QN(n2703) );
  sdffs1 \DFF_373/Q_reg  ( .DIN(g8286), .SDIN(n3158), .SSEL(test_se), .CLK(CK), 
        .Q(n3159), .QN(n2504) );
  sdffs1 \DFF_372/Q_reg  ( .DIN(g6843), .SDIN(n3157), .SSEL(test_se), .CLK(CK), 
        .Q(n3158), .QN(n2725) );
  sdffs1 \DFF_371/Q_reg  ( .DIN(g7360), .SDIN(n3156), .SSEL(test_se), .CLK(CK), 
        .Q(n3157), .QN(n2798) );
  sdffs1 \DFF_370/Q_reg  ( .DIN(g10880), .SDIN(n3155), .SSEL(test_se), .CLK(CK), .Q(n3156), .QN(n2766) );
  sdffs1 \DFF_369/Q_reg  ( .DIN(g9827), .SDIN(n3154), .SSEL(test_se), .CLK(CK), 
        .Q(n3155), .QN(n1980) );
  sdffs1 \DFF_368/Q_reg  ( .DIN(g11258), .SDIN(n3153), .SSEL(test_se), .CLK(CK), .Q(n3154), .QN(n2678) );
  sdffs1 \DFF_367/Q_reg  ( .DIN(g4189), .SDIN(n3152), .SSEL(test_se), .CLK(CK), 
        .Q(n3153), .QN(n2661) );
  sdffs1 \DFF_366/Q_reg  ( .DIN(g6308), .SDIN(n3151), .SSEL(test_se), .CLK(CK), 
        .Q(n3152), .QN(n1945) );
  sdffs1 \DFF_365/Q_reg  ( .DIN(g11400), .SDIN(n3150), .SSEL(test_se), .CLK(CK), .Q(n3151), .QN(n2788) );
  sdffs1 \DFF_364/Q_reg  ( .DIN(g7749), .SDIN(g8986), .SSEL(test_se), .CLK(CK), 
        .Q(n3150), .QN(n2817) );
  sdffs1 \DFF_363/Q_reg  ( .DIN(g7776), .SDIN(n3149), .SSEL(test_se), .CLK(CK), 
        .Q(g8986), .QN(n2022) );
  sdffs1 \DFF_362/Q_reg  ( .DIN(g9820), .SDIN(n3148), .SSEL(test_se), .CLK(CK), 
        .Q(n3149), .QN(n1978) );
  sdffs1 \DFF_361/Q_reg  ( .DIN(g8276), .SDIN(g2613), .SSEL(test_se), .CLK(CK), 
        .Q(n3148), .QN(n2602) );
  sdffs1 \DFF_360/Q_reg  ( .DIN(g8781), .SDIN(n3147), .SSEL(test_se), .CLK(CK), 
        .Q(g2613) );
  sdffs1 \DFF_359/Q_reg  ( .DIN(g9347), .SDIN(n3146), .SSEL(test_se), .CLK(CK), 
        .Q(n3147), .QN(n2009) );
  sdffs1 \DFF_358/Q_reg  ( .DIN(g9818), .SDIN(g874), .SSEL(test_se), .CLK(CK), 
        .Q(n3146), .QN(n1951) );
  sdffs1 \DFF_357/Q_reg  ( .DIN(g9821), .SDIN(g5646), .SSEL(test_se), .CLK(CK), 
        .Q(g874) );
  sdffs1 \DFF_356/Q_reg  ( .DIN(g7753), .SDIN(n3145), .SSEL(test_se), .CLK(CK), 
        .Q(g5646) );
  sdffs1 \DFF_355/Q_reg  ( .DIN(g7300), .SDIN(n3144), .SSEL(test_se), .CLK(CK), 
        .Q(n3145), .QN(n2616) );
  sdffs1 \DFF_354/Q_reg  ( .DIN(g9350), .SDIN(n3143), .SSEL(test_se), .CLK(CK), 
        .Q(n3144), .QN(n2010) );
  sdffs1 \DFF_353/Q_reg  ( .DIN(g6310), .SDIN(n2627), .SSEL(test_se), .CLK(CK), 
        .Q(n3143), .QN(n2013) );
  sdffs1 \DFF_352/Q_reg  ( .DIN(g5673), .SDIN(n3142), .SSEL(test_se), .CLK(CK), 
        .Q(n2627) );
  sdffs1 \DFF_351/Q_reg  ( .DIN(g11406), .SDIN(g37), .SSEL(test_se), .CLK(CK), 
        .Q(n3142), .QN(n2808) );
  sdffs1 \DFF_350/Q_reg  ( .DIN(n2822), .SDIN(n3141), .SSEL(test_se), .CLK(CK), 
        .Q(g37) );
  sdffs1 \DFF_349/Q_reg  ( .DIN(g8281), .SDIN(g4190), .SSEL(test_se), .CLK(CK), 
        .Q(n3141), .QN(n2509) );
  sdffs1 \DFF_347/Q_reg  ( .DIN(g8568), .SDIN(n3140), .SSEL(test_se), .CLK(CK), 
        .Q(g4190), .QN(n2492) );
  sdffs1 \DFF_346/Q_reg  ( .DIN(g8573), .SDIN(n3139), .SSEL(test_se), .CLK(CK), 
        .Q(n3140), .QN(n2628) );
  sdffs1 \DFF_345/Q_reg  ( .DIN(g7763), .SDIN(n3138), .SSEL(test_se), .CLK(CK), 
        .Q(n3139), .QN(n2753) );
  sdffs1 \DFF_344/Q_reg  ( .DIN(g11654), .SDIN(n3137), .SSEL(test_se), .CLK(CK), .Q(n3138), .QN(n2796) );
  sdffs1 \DFF_343/Q_reg  ( .DIN(g4187), .SDIN(n3136), .SSEL(test_se), .CLK(CK), 
        .Q(n3137), .QN(n2657) );
  sdffs1 \DFF_342/Q_reg  ( .DIN(g11629), .SDIN(n3135), .SSEL(test_se), .CLK(CK), .Q(n3136), .QN(n2786) );
  sdffs1 \DFF_340/Q_reg  ( .DIN(g8571), .SDIN(n3134), .SSEL(test_se), .CLK(CK), 
        .Q(n3135), .QN(n2046) );
  sdffs1 \DFF_339/Q_reg  ( .DIN(g8285), .SDIN(n3133), .SSEL(test_se), .CLK(CK), 
        .Q(n3134), .QN(n2505) );
  sdffs1 \DFF_338/Q_reg  ( .DIN(g4183), .SDIN(n3132), .SSEL(test_se), .CLK(CK), 
        .Q(n3133), .QN(n2664) );
  sdffs1 \DFF_337/Q_reg  ( .DIN(g8427), .SDIN(n3131), .SSEL(test_se), .CLK(CK), 
        .Q(n3132), .QN(n1926) );
  sdffs1 \DFF_336/Q_reg  ( .DIN(g7287), .SDIN(n3130), .SSEL(test_se), .CLK(CK), 
        .Q(n3131), .QN(\DFF_336/net623 ) );
  sdffs1 \DFF_335/Q_reg  ( .DIN(n545), .SDIN(n3129), .SSEL(test_se), .CLK(CK), 
        .Q(n3130), .QN(n2011) );
  sdffs1 \DFF_334/Q_reg  ( .DIN(g7298), .SDIN(n3128), .SSEL(test_se), .CLK(CK), 
        .Q(n3129), .QN(n2612) );
  sdffs1 \DFF_333/Q_reg  ( .DIN(g9351), .SDIN(n3127), .SSEL(test_se), .CLK(CK), 
        .Q(n3128), .QN(n1932) );
  sdffs1 \DFF_332/Q_reg  ( .DIN(g7813), .SDIN(n3126), .SSEL(test_se), .CLK(CK), 
        .Q(n3127), .QN(n1984) );
  sdffs1 \DFF_331/Q_reg  ( .DIN(g7313), .SDIN(n3125), .SSEL(test_se), .CLK(CK), 
        .Q(n3126), .QN(n1962) );
  sdffs1 \DFF_330/Q_reg  ( .DIN(g5670), .SDIN(n3124), .SSEL(test_se), .CLK(CK), 
        .Q(n3125), .QN(\DFF_330/net617 ) );
  sdffs1 \DFF_329/Q_reg  ( .DIN(g11332), .SDIN(g3069), .SSEL(test_se), .CLK(CK), .Q(n3124), .QN(n2638) );
  sdffs1 \DFF_328/Q_reg  ( .DIN(g4898), .SDIN(n2551), .SSEL(test_se), .CLK(CK), 
        .Q(g3069) );
  sdffs1 \DFF_327/Q_reg  ( .DIN(g7312), .SDIN(n3123), .SSEL(test_se), .CLK(CK), 
        .Q(n2551) );
  sdffs1 \DFF_326/Q_reg  ( .DIN(g7343), .SDIN(n3122), .SSEL(test_se), .CLK(CK), 
        .Q(n3123), .QN(n2736) );
  sdffs1 \DFF_325/Q_reg  ( .DIN(g11632), .SDIN(n3121), .SSEL(test_se), .CLK(CK), .Q(n3122), .QN(n2750) );
  sdffs1 \DFF_324/Q_reg  ( .DIN(g8280), .SDIN(n3120), .SSEL(test_se), .CLK(CK), 
        .Q(n3121), .QN(n1952) );
  sdffs1 \DFF_323/Q_reg  ( .DIN(g6845), .SDIN(n3119), .SSEL(test_se), .CLK(CK), 
        .Q(n3120), .QN(n2727) );
  sdffs1 \DFF_322/Q_reg  ( .DIN(g7303), .SDIN(n3118), .SSEL(test_se), .CLK(CK), 
        .Q(n3119), .QN(n2606) );
  sdffs1 \DFF_321/Q_reg  ( .DIN(g10882), .SDIN(g1765), .SSEL(test_se), .CLK(CK), .Q(n3118), .QN(n2746) );
  sdffs1 \DFF_320/Q_reg  ( .DIN(g3329), .SDIN(n3117), .SSEL(test_se), .CLK(CK), 
        .Q(g1765) );
  sdffs1 \DFF_319/Q_reg  ( .DIN(n2824), .SDIN(g2044), .SSEL(test_se), .CLK(CK), 
        .Q(n3117), .QN(\DFF_319/net606 ) );
  sdffs1 \DFF_318/Q_reg  ( .DIN(g6339), .SDIN(n3116), .SSEL(test_se), .CLK(CK), 
        .Q(g2044) );
  sdffs1 \DFF_317/Q_reg  ( .DIN(g11401), .SDIN(n3115), .SSEL(test_se), .CLK(CK), .Q(n3116), .QN(n2774) );
  sdffs1 \DFF_316/Q_reg  ( .DIN(g9342), .SDIN(n3114), .SSEL(test_se), .CLK(CK), 
        .Q(n3115), .QN(n1933) );
  sdffs1 \DFF_315/Q_reg  ( .DIN(g7334), .SDIN(n3113), .SSEL(test_se), .CLK(CK), 
        .Q(n3114), .QN(n2537) );
  sdffs1 \DFF_314/Q_reg  ( .DIN(g8422), .SDIN(n3112), .SSEL(test_se), .CLK(CK), 
        .Q(n3113), .QN(n2519) );
  sdffs1 \DFF_313/Q_reg  ( .DIN(g8287), .SDIN(n3111), .SSEL(test_se), .CLK(CK), 
        .Q(n3112), .QN(n2503) );
  sdffs1 \DFF_312/Q_reg  ( .DIN(g11398), .SDIN(g2731), .SSEL(test_se), .CLK(CK), .Q(n3111), .QN(n2807) );
  sdffs1 \DFF_311/Q_reg  ( .DIN(g11408), .SDIN(n3110), .SSEL(test_se), .CLK(CK), .Q(g2731) );
  sdffs1 \DFF_310/Q_reg  ( .DIN(g9819), .SDIN(n3109), .SSEL(test_se), .CLK(CK), 
        .Q(n3110), .QN(n1985) );
  sdffs1 \DFF_309/Q_reg  ( .DIN(g4184), .SDIN(n3108), .SSEL(test_se), .CLK(CK), 
        .Q(n3109), .QN(n2663) );
  sdffs1 \DFF_308/Q_reg  ( .DIN(g11512), .SDIN(n3107), .SSEL(test_se), .CLK(CK), .Q(n3108), .QN(n2591) );
  sdffs1 \DFF_307/Q_reg  ( .DIN(g7748), .SDIN(n3106), .SSEL(test_se), .CLK(CK), 
        .Q(n3107), .QN(n2521) );
  sdffs1 \DFF_306/Q_reg  ( .DIN(g8438), .SDIN(g2639), .SSEL(test_se), .CLK(CK), 
        .Q(n3106), .QN(n2528) );
  sdffs1 \DFF_304/Q_reg  ( .DIN(g2638), .SDIN(n3105), .SSEL(test_se), .CLK(CK), 
        .Q(g2639), .QN(n2577) );
  sdffs1 \DFF_303/Q_reg  ( .DIN(g7306), .SDIN(n3104), .SSEL(test_se), .CLK(CK), 
        .Q(n3105), .QN(n1939) );
  sdffs1 \DFF_302/Q_reg  ( .DIN(g9826), .SDIN(g4179), .SSEL(test_se), .CLK(CK), 
        .Q(n3104), .QN(n1953) );
  sdffs1 \DFF_301/Q_reg  ( .DIN(g8273), .SDIN(n3103), .SSEL(test_se), .CLK(CK), 
        .Q(g4179), .QN(n2056) );
  sdffs1 \DFF_300/Q_reg  ( .DIN(g9353), .SDIN(n3102), .SSEL(test_se), .CLK(CK), 
        .Q(n3103), .QN(n2028) );
  sdffs1 \DFF_299/Q_reg  ( .DIN(g1217), .SDIN(n3101), .SSEL(test_se), .CLK(CK), 
        .Q(n3102), .QN(n2578) );
  sdffs1 \DFF_297/Q_reg  ( .DIN(g9825), .SDIN(n3100), .SSEL(test_se), .CLK(CK), 
        .Q(n3101), .QN(n1986) );
  sdffs1 \DFF_296/Q_reg  ( .DIN(g7746), .SDIN(g1955), .SSEL(test_se), .CLK(CK), 
        .Q(n3100), .QN(n1925) );
  sdffs1 \DFF_295/Q_reg  ( .DIN(g6265), .SDIN(n3099), .SSEL(test_se), .CLK(CK), 
        .Q(g1955) );
  sdffs1 \DFF_294/Q_reg  ( .DIN(g11470), .SDIN(n3098), .SSEL(test_se), .CLK(CK), .Q(n3099), .QN(n2787) );
  sdffs1 \DFF_293/Q_reg  ( .DIN(g11473), .SDIN(n3097), .SSEL(test_se), .CLK(CK), .Q(n3098), .QN(n2748) );
  sdffs1 \DFF_292/Q_reg  ( .DIN(g6804), .SDIN(g2986), .SSEL(test_se), .CLK(CK), 
        .Q(n3097), .QN(n2571) );
  sdffs1 \DFF_291/Q_reg  ( .DIN(g4897), .SDIN(n3096), .SSEL(test_se), .CLK(CK), 
        .Q(g2986) );
  sdffs1 \DFF_290/Q_reg  ( .DIN(g6809), .SDIN(n2545), .SSEL(test_se), .CLK(CK), 
        .Q(n3096), .QN(n2566) );
  sdffs1 \DFF_289/Q_reg  ( .DIN(g7809), .SDIN(n3095), .SSEL(test_se), .CLK(CK), 
        .Q(n2545) );
  sdffs1 \DFF_288/Q_reg  ( .DIN(g11051), .SDIN(g8980), .SSEL(test_se), .CLK(CK), .Q(n3095), .QN(n2693) );
  sdffs1 \DFF_287/Q_reg  ( .DIN(g7780), .SDIN(n3094), .SSEL(test_se), .CLK(CK), 
        .Q(g8980), .QN(n2036) );
  sdffs1 \DFF_286/Q_reg  ( .DIN(g9346), .SDIN(n3093), .SSEL(test_se), .CLK(CK), 
        .Q(n3094), .QN(n1994) );
  sdffs1 \DFF_285/Q_reg  ( .DIN(g10875), .SDIN(n3092), .SSEL(test_se), .CLK(CK), .Q(n3093), .QN(n2720) );
  sdffs1 \DFF_284/Q_reg  ( .DIN(g6837), .SDIN(n3091), .SSEL(test_se), .CLK(CK), 
        .Q(n3092), .QN(n1946) );
  sdffs1 \DFF_283/Q_reg  ( .DIN(g11510), .SDIN(n3090), .SSEL(test_se), .CLK(CK), .Q(n3091), .QN(n2593) );
  sdffs1 \DFF_282/Q_reg  ( .DIN(g5669), .SDIN(n3089), .SSEL(test_se), .CLK(CK), 
        .Q(n3090), .QN(n2811) );
  sdffs1 \DFF_281/Q_reg  ( .DIN(g8431), .SDIN(n3088), .SSEL(test_se), .CLK(CK), 
        .Q(n3089), .QN(n2497) );
  sdffs1 \DFF_280/Q_reg  ( .DIN(g11034), .SDIN(n3087), .SSEL(test_se), .CLK(CK), .Q(n3088), .QN(n2714) );
  sdffs1 \DFF_279/Q_reg  ( .DIN(g7771), .SDIN(n3086), .SSEL(test_se), .CLK(CK), 
        .Q(n3087), .QN(n2754) );
  sdffs1 \DFF_278/Q_reg  ( .DIN(g6817), .SDIN(n3085), .SSEL(test_se), .CLK(CK), 
        .Q(n3086), .QN(n1949) );
  sdffs1 \DFF_277/Q_reg  ( .DIN(g8443), .SDIN(n3084), .SSEL(test_se), .CLK(CK), 
        .Q(n3085), .QN(n2533) );
  sdffs1 \DFF_276/Q_reg  ( .DIN(g6844), .SDIN(n3083), .SSEL(test_se), .CLK(CK), 
        .Q(n3084), .QN(n2074) );
  sdffs1 \DFF_275/Q_reg  ( .DIN(n873), .SDIN(n3082), .SSEL(test_se), .CLK(CK), 
        .Q(n3083), .QN(\DFF_275/net562 ) );
  sdffs1 \DFF_273/Q_reg  ( .DIN(g8442), .SDIN(n3081), .SSEL(test_se), .CLK(CK), 
        .Q(n3082), .QN(n2532) );
  sdffs1 \DFF_272/Q_reg  ( .DIN(g5661), .SDIN(n3080), .SSEL(test_se), .CLK(CK), 
        .Q(n3081), .QN(n2813) );
  sdffs1 \DFF_271/Q_reg  ( .DIN(g9356), .SDIN(g5644), .SSEL(test_se), .CLK(CK), 
        .Q(n3080), .QN(n2008) );
  sdffs1 \DFF_270/Q_reg  ( .DIN(g7751), .SDIN(g2648), .SSEL(test_se), .CLK(CK), 
        .Q(g5644) );
  sdffs1 \DFF_269/Q_reg  ( .DIN(n2826), .SDIN(n3079), .SSEL(test_se), .CLK(CK), 
        .Q(g2648) );
  sdffs1 \DFF_268/Q_reg  ( .DIN(g7811), .SDIN(g8), .SSEL(test_se), .CLK(CK), 
        .Q(n3079), .QN(n2620) );
  sdffs1 \DFF_267/Q_reg  ( .DIN(g2613), .SDIN(n3078), .SSEL(test_se), .CLK(CK), 
        .Q(g8) );
  sdffs1 \DFF_266/Q_reg  ( .DIN(g11642), .SDIN(n3077), .SSEL(test_se), .CLK(CK), .Q(n3078), .QN(n2580) );
  sdffs1 \DFF_265/Q_reg  ( .DIN(g5643), .SDIN(n3076), .SSEL(test_se), .CLK(CK), 
        .Q(n3077), .QN(n2669) );
  sdffs1 \DFF_264/Q_reg  ( .DIN(g11466), .SDIN(n3075), .SSEL(test_se), .CLK(CK), .Q(n3076), .QN(n2073) );
  sdffs1 \DFF_263/Q_reg  ( .DIN(g11653), .SDIN(g17), .SSEL(test_se), .CLK(CK), 
        .Q(n3075), .QN(n2579) );
  sdffs1 \DFF_262/Q_reg  ( .DIN(g4894), .SDIN(n3074), .SSEL(test_se), .CLK(CK), 
        .Q(g17) );
  sdffs1 \DFF_261/Q_reg  ( .DIN(g8780), .SDIN(n3073), .SSEL(test_se), .CLK(CK), 
        .Q(n3074), .QN(n1982) );
  sdffs1 \DFF_260/Q_reg  ( .DIN(g11049), .SDIN(n3072), .SSEL(test_se), .CLK(CK), .Q(n3073), .QN(n2695) );
  sdffs1 \DFF_259/Q_reg  ( .DIN(g7768), .SDIN(n3071), .SSEL(test_se), .CLK(CK), 
        .Q(n3072), .QN(n2794) );
  sdffs1 \DFF_258/Q_reg  ( .DIN(g7345), .SDIN(n3070), .SSEL(test_se), .CLK(CK), 
        .Q(n3071), .QN(n2805) );
  sdffs1 \DFF_256/Q_reg  ( .DIN(g7350), .SDIN(n3069), .SSEL(test_se), .CLK(CK), 
        .Q(n3070), .QN(n2741) );
  sdffs1 \DFF_255/Q_reg  ( .DIN(g11468), .SDIN(n3068), .SSEL(test_se), .CLK(CK), .Q(n3069), .QN(n1977) );
  sdffs1 \DFF_254/Q_reg  ( .DIN(g7357), .SDIN(g4176), .SSEL(test_se), .CLK(CK), 
        .Q(n3068), .QN(n2729) );
  sdffs1 \DFF_253/Q_reg  ( .DIN(g7288), .SDIN(g1850), .SSEL(test_se), .CLK(CK), 
        .Q(g4176), .QN(n2557) );
  sdffs1 \DFF_252/Q_reg  ( .DIN(g5671), .SDIN(n3067), .SSEL(test_se), .CLK(CK), 
        .Q(g1850) );
  sdffs1 \DFF_251/Q_reg  ( .DIN(g7769), .SDIN(n3066), .SSEL(test_se), .CLK(CK), 
        .Q(n3067), .QN(n2780) );
  sdffs1 \DFF_250/Q_reg  ( .DIN(g7293), .SDIN(n3065), .SSEL(test_se), .CLK(CK), 
        .Q(n3066), .QN(n2610) );
  sdffs1 \DFF_249/Q_reg  ( .DIN(g8871), .SDIN(n3064), .SSEL(test_se), .CLK(CK), 
        .Q(n3065), .QN(n2701) );
  sdffs1 \DFF_248/Q_reg  ( .DIN(g4190), .SDIN(g4178), .SSEL(test_se), .CLK(CK), 
        .Q(n3064), .QN(n2660) );
  sdffs1 \DFF_247/Q_reg  ( .DIN(g8076), .SDIN(g5652), .SSEL(test_se), .CLK(CK), 
        .Q(g4178), .QN(n2513) );
  sdffs1 \DFF_246/Q_reg  ( .DIN(g7759), .SDIN(n3063), .SSEL(test_se), .CLK(CK), 
        .Q(g5652) );
  sdffs1 \DFF_245/Q_reg  ( .DIN(g11337), .SDIN(g5650), .SSEL(test_se), .CLK(CK), .Q(n3063), .QN(n2630) );
  sdffs1 \DFF_244/Q_reg  ( .DIN(g7757), .SDIN(n3062), .SSEL(test_se), .CLK(CK), 
        .Q(g5650) );
  sdffs1 \DFF_243/Q_reg  ( .DIN(g8569), .SDIN(n3061), .SSEL(test_se), .CLK(CK), 
        .Q(n3062), .QN(n2047) );
  sdffs1 \DFF_242/Q_reg  ( .DIN(n2820), .SDIN(n3060), .SSEL(test_se), .CLK(CK), 
        .Q(n3061), .QN(\DFF_242/net529 ) );
  sdffs1 \DFF_241/Q_reg  ( .DIN(g6330), .SDIN(n2584), .SSEL(test_se), .CLK(CK), 
        .Q(n3060), .QN(n2724) );
  sdffs1 \DFF_240/Q_reg  ( .DIN(g6303), .SDIN(n3059), .SSEL(test_se), .CLK(CK), 
        .Q(n2584) );
  sdffs1 \DFF_239/Q_reg  ( .DIN(g5650), .SDIN(n3058), .SSEL(test_se), .CLK(CK), 
        .Q(n3059), .QN(n2690) );
  sdffs1 \DFF_238/Q_reg  ( .DIN(g11511), .SDIN(n3057), .SSEL(test_se), .CLK(CK), .Q(n3058), .QN(n2592) );
  sdffs1 \DFF_237/Q_reg  ( .DIN(g7326), .SDIN(n3056), .SSEL(test_se), .CLK(CK), 
        .Q(n3057), .QN(n2012) );
  sdffs1 \DFF_235/Q_reg  ( .DIN(g8990), .SDIN(n3055), .SSEL(test_se), .CLK(CK), 
        .Q(n3056), .QN(n2525) );
  sdffs1 \DFF_234/Q_reg  ( .DIN(g7800), .SDIN(n3054), .SSEL(test_se), .CLK(CK), 
        .Q(n3055), .QN(n2600) );
  sdffs1 \DFF_233/Q_reg  ( .DIN(g2044), .SDIN(n2582), .SSEL(test_se), .CLK(CK), 
        .Q(n3054), .QN(g8271) );
  sdffs1 \DFF_232/Q_reg  ( .DIN(g6301), .SDIN(n3053), .SSEL(test_se), .CLK(CK), 
        .Q(n2582) );
  sdffs1 \DFF_231/Q_reg  ( .DIN(g7299), .SDIN(n3052), .SSEL(test_se), .CLK(CK), 
        .Q(n3053), .QN(n2614) );
  sdffs1 \DFF_230/Q_reg  ( .DIN(g11513), .SDIN(n3051), .SSEL(test_se), .CLK(CK), .Q(n3052), .QN(n2590) );
  sdffs1 \DFF_229/Q_reg  ( .DIN(g7773), .SDIN(n3050), .SSEL(test_se), .CLK(CK), 
        .Q(n3051), .QN(n2733) );
  sdffs1 \DFF_228/Q_reg  ( .DIN(n2823), .SDIN(g4182), .SSEL(test_se), .CLK(CK), 
        .Q(n3050), .QN(\DFF_228/net515 ) );
  sdffs1 \DFF_227/Q_reg  ( .DIN(g6800), .SDIN(g1356), .SSEL(test_se), .CLK(CK), 
        .Q(g4182), .QN(n2573) );
  sdffs1 \DFF_226/Q_reg  ( .DIN(g6818), .SDIN(n3049), .SSEL(test_se), .CLK(CK), 
        .Q(g1356) );
  sdffs1 \DFF_225/Q_reg  ( .DIN(g5646), .SDIN(g8983), .SSEL(test_se), .CLK(CK), 
        .Q(n3049), .QN(n2665) );
  sdffs1 \DFF_224/Q_reg  ( .DIN(g7783), .SDIN(n3048), .SSEL(test_se), .CLK(CK), 
        .Q(g8983), .QN(n2018) );
  sdffs1 \DFF_223/Q_reg  ( .DIN(g8694), .SDIN(g5651), .SSEL(test_se), .CLK(CK), 
        .Q(n3048), .QN(n1983) );
  sdffs1 \DFF_222/Q_reg  ( .DIN(g7758), .SDIN(n3047), .SSEL(test_se), .CLK(CK), 
        .Q(g5651) );
  sdffs1 \DFF_221/Q_reg  ( .DIN(g11334), .SDIN(n3046), .SSEL(test_se), .CLK(CK), .Q(n3047), .QN(n2639) );
  sdffs1 \DFF_220/Q_reg  ( .DIN(g7747), .SDIN(n3045), .SSEL(test_se), .CLK(CK), 
        .Q(n3046), .QN(n2518) );
  sdffs1 \DFF_218/Q_reg  ( .DIN(g7363), .SDIN(n3044), .SSEL(test_se), .CLK(CK), 
        .Q(n3045), .QN(n2755) );
  sdffs1 \DFF_217/Q_reg  ( .DIN(g11263), .SDIN(n3043), .SSEL(test_se), .CLK(CK), .Q(n3044), .QN(n2681) );
  sdffs1 \DFF_216/Q_reg  ( .DIN(g11509), .SDIN(g1317), .SSEL(test_se), .CLK(CK), .Q(n3043), .QN(n2594) );
  sdffs1 \DFF_215/Q_reg  ( .DIN(g1356), .SDIN(n3042), .SSEL(test_se), .CLK(CK), 
        .Q(g1317) );
  sdffs1 \DFF_214/Q_reg  ( .DIN(g6299), .SDIN(g8978), .SSEL(test_se), .CLK(CK), 
        .Q(n3042), .QN(n1969) );
  sdffs1 \DFF_213/Q_reg  ( .DIN(g7778), .SDIN(n3041), .SSEL(test_se), .CLK(CK), 
        .Q(g8978), .QN(n2037) );
  sdffs1 \DFF_212/Q_reg  ( .DIN(g9355), .SDIN(n3040), .SSEL(test_se), .CLK(CK), 
        .Q(n3041), .QN(n1993) );
  sdffs1 \DFF_211/Q_reg  ( .DIN(g11052), .SDIN(n3039), .SSEL(test_se), .CLK(CK), .Q(n3040), .QN(n2692) );
  sdffs1 \DFF_210/Q_reg  ( .DIN(g11328), .SDIN(n3038), .SSEL(test_se), .CLK(CK), .Q(n3039), .QN(n2635) );
  sdffs1 \DFF_209/Q_reg  ( .DIN(g8284), .SDIN(n3037), .SSEL(test_se), .CLK(CK), 
        .Q(n3038), .QN(n2506) );
  sdffs1 \DFF_208/Q_reg  ( .DIN(g11050), .SDIN(n3036), .SSEL(test_se), .CLK(CK), .Q(n3037), .QN(n2694) );
  sdffs1 \DFF_207/Q_reg  ( .DIN(g11440), .SDIN(n3035), .SSEL(test_se), .CLK(CK), .Q(n3036), .QN(n2673) );
  sdffs1 \DFF_206/Q_reg  ( .DIN(g11040), .SDIN(n3034), .SSEL(test_se), .CLK(CK), .Q(n3035), .QN(n2704) );
  sdffs1 \DFF_205/Q_reg  ( .DIN(g11325), .SDIN(n3033), .SSEL(test_se), .CLK(CK), .Q(n3034), .QN(n2632) );
  sdffs1 \DFF_204/Q_reg  ( .DIN(g11269), .SDIN(n3032), .SSEL(test_se), .CLK(CK), .Q(n3033), .QN(n2674) );
  sdffs1 \DFF_203/Q_reg  ( .DIN(g11326), .SDIN(n3031), .SSEL(test_se), .CLK(CK), .Q(n3032), .QN(n2633) );
  sdffs1 \DFF_202/Q_reg  ( .DIN(g7297), .SDIN(n3030), .SSEL(test_se), .CLK(CK), 
        .Q(n3031), .QN(n2613) );
  sdffs1 \DFF_201/Q_reg  ( .DIN(g7329), .SDIN(n3029), .SSEL(test_se), .CLK(CK), 
        .Q(n3030), .QN(n2544) );
  sdffs1 \DFF_200/Q_reg  ( .DIN(g5666), .SDIN(n3028), .SSEL(test_se), .CLK(CK), 
        .Q(n3029), .QN(n2751) );
  sdffs1 \DFF_199/Q_reg  ( .DIN(g8873), .SDIN(n3027), .SSEL(test_se), .CLK(CK), 
        .Q(n3028), .QN(n2721) );
  sdffs1 \DFF_198/Q_reg  ( .DIN(g11656), .SDIN(n3026), .SSEL(test_se), .CLK(CK), .Q(n3027), .QN(n2000) );
  sdffs1 \DFF_197/Q_reg  ( .DIN(g7770), .SDIN(n3025), .SSEL(test_se), .CLK(CK), 
        .Q(n3026), .QN(n2768) );
  sdffs1 \DFF_196/Q_reg  ( .DIN(g8067), .SDIN(n3024), .SSEL(test_se), .CLK(CK), 
        .Q(n3025), .QN(n2514) );
  sdffs1 \DFF_195/Q_reg  ( .DIN(g11633), .SDIN(n3023), .SSEL(test_se), .CLK(CK), .Q(n3024), .QN(n2742) );
  sdffs1 \DFF_194/Q_reg  ( .DIN(g3069), .SDIN(g5648), .SSEL(test_se), .CLK(CK), 
        .Q(n3023), .QN(\DFF_194/net481 ) );
  sdffs1 \DFF_193/Q_reg  ( .DIN(g7755), .SDIN(n3022), .SSEL(test_se), .CLK(CK), 
        .Q(g5648) );
  sdffs1 \DFF_192/Q_reg  ( .DIN(g7799), .SDIN(n2558), .SSEL(test_se), .CLK(CK), 
        .Q(n3022), .QN(n2653) );
  sdffs1 \DFF_191/Q_reg  ( .DIN(g5657), .SDIN(n3021), .SSEL(test_se), .CLK(CK), 
        .Q(n2558) );
  sdffs1 \DFF_190/Q_reg  ( .DIN(g8425), .SDIN(n2552), .SSEL(test_se), .CLK(CK), 
        .Q(n3021), .QN(n1992) );
  sdffs1 \DFF_189/Q_reg  ( .DIN(g7316), .SDIN(n3020), .SSEL(test_se), .CLK(CK), 
        .Q(n2552) );
  sdffs1 \DFF_188/Q_reg  ( .DIN(g875), .SDIN(g2612), .SSEL(test_se), .CLK(CK), 
        .Q(n3020), .QN(n2618) );
  sdffs1 \DFF_187/Q_reg  ( .DIN(g6283), .SDIN(n3019), .SSEL(test_se), .CLK(CK), 
        .Q(g2612) );
  sdffs1 \DFF_186/Q_reg  ( .DIN(g11048), .SDIN(n3018), .SSEL(test_se), .CLK(CK), .Q(n3019), .QN(n2696) );
  sdffs1 \DFF_185/Q_reg  ( .DIN(g7319), .SDIN(g4187), .SSEL(test_se), .CLK(CK), 
        .Q(n3018), .QN(n1947) );
  sdffs1 \DFF_184/Q_reg  ( .DIN(g8077), .SDIN(n3017), .SSEL(test_se), .CLK(CK), 
        .Q(g4187), .QN(n2512) );
  sdffs1 \DFF_183/Q_reg  ( .DIN(g5652), .SDIN(n2546), .SSEL(test_se), .CLK(CK), 
        .Q(n3017), .QN(n2667) );
  sdffs1 \DFF_182/Q_reg  ( .DIN(g7324), .SDIN(n3016), .SSEL(test_se), .CLK(CK), 
        .Q(n2546) );
  sdffs1 \DFF_181/Q_reg  ( .DIN(g11405), .SDIN(n3015), .SSEL(test_se), .CLK(CK), .Q(n3016), .QN(n2731) );
  sdffs1 \DFF_180/Q_reg  ( .DIN(g8782), .SDIN(n3014), .SSEL(test_se), .CLK(CK), 
        .Q(n3015), .QN(n2501) );
  sdffs1 \DFF_179/Q_reg  ( .DIN(g7336), .SDIN(n3013), .SSEL(test_se), .CLK(CK), 
        .Q(n3014), .QN(n2763) );
  sdffs1 \DFF_178/Q_reg  ( .DIN(g11409), .SDIN(n3012), .SSEL(test_se), .CLK(CK), .Q(n3013), .QN(n1989) );
  sdffs1 \DFF_177/Q_reg  ( .DIN(g11266), .SDIN(n3011), .SSEL(test_se), .CLK(CK), .Q(n3012), .QN(n2685) );
  sdffs1 \DFF_176/Q_reg  ( .DIN(g7762), .SDIN(n3010), .SSEL(test_se), .CLK(CK), 
        .Q(n3011), .QN(n2767) );
  sdffs1 \DFF_175/Q_reg  ( .DIN(g5651), .SDIN(n3009), .SSEL(test_se), .CLK(CK), 
        .Q(n3010), .QN(n2688) );
  sdffs1 \DFF_174/Q_reg  ( .DIN(g6336), .SDIN(n3008), .SSEL(test_se), .CLK(CK), 
        .Q(n3009), .QN(n2061) );
  sdffs1 \DFF_173/Q_reg  ( .DIN(g6806), .SDIN(n3007), .SSEL(test_se), .CLK(CK), 
        .Q(n3008), .QN(n2569) );
  sdffs1 \DFF_172/Q_reg  ( .DIN(g8441), .SDIN(n3006), .SSEL(test_se), .CLK(CK), 
        .Q(n3007), .QN(n2531) );
  sdffs1 \DFF_171/Q_reg  ( .DIN(g11259), .SDIN(n3005), .SSEL(test_se), .CLK(CK), .Q(n3006), .QN(n2679) );
  sdffs1 \DFF_170/Q_reg  ( .DIN(g6813), .SDIN(n3004), .SSEL(test_se), .CLK(CK), 
        .Q(n3005), .QN(n2562) );
  sdffs1 \DFF_169/Q_reg  ( .DIN(g7331), .SDIN(n2790), .SSEL(test_se), .CLK(CK), 
        .Q(n3004), .QN(n2538) );
  sdffs1 \DFF_168/Q_reg  ( .DIN(n2821), .SDIN(n3003), .SSEL(test_se), .CLK(CK), 
        .Q(n2790) );
  sdffs1 \DFF_167/Q_reg  ( .DIN(g7805), .SDIN(n3002), .SSEL(test_se), .CLK(CK), 
        .Q(n3003), .QN(n2651) );
  sdffs1 \DFF_166/Q_reg  ( .DIN(g10877), .SDIN(n3001), .SSEL(test_se), .CLK(CK), .Q(n3002), .QN(n2718) );
  sdffs1 \DFF_165/Q_reg  ( .DIN(g7327), .SDIN(n3000), .SSEL(test_se), .CLK(CK), 
        .Q(n3001), .QN(n1991) );
  sdffs1 \DFF_164/Q_reg  ( .DIN(g7340), .SDIN(n2547), .SSEL(test_se), .CLK(CK), 
        .Q(n3000), .QN(n2771) );
  sdffs1 \DFF_163/Q_reg  ( .DIN(g7308), .SDIN(n2999), .SSEL(test_se), .CLK(CK), 
        .Q(n2547) );
  sdffs1 \DFF_162/Q_reg  ( .DIN(g11036), .SDIN(n2998), .SSEL(test_se), .CLK(CK), .Q(n2999), .QN(n2712) );
  sdffs1 \DFF_161/Q_reg  ( .DIN(g11180), .SDIN(n2997), .SSEL(test_se), .CLK(CK), .Q(n2998), .QN(n2726) );
  sdffs1 \DFF_159/Q_reg  ( .DIN(g11044), .SDIN(n2996), .SSEL(test_se), .CLK(CK), .Q(n2997), .QN(n2698) );
  sdffs1 \DFF_158/Q_reg  ( .DIN(g6814), .SDIN(n2995), .SSEL(test_se), .CLK(CK), 
        .Q(n2996), .QN(n1974) );
  sdffs1 \DFF_157/Q_reg  ( .DIN(g5656), .SDIN(g2638), .SSEL(test_se), .CLK(CK), 
        .Q(n2995), .QN(\DFF_157/net444 ) );
  sdffs1 \DFF_156/Q_reg  ( .DIN(g755), .SDIN(n2994), .SSEL(test_se), .CLK(CK), 
        .Q(g2638) );
  sdffs1 \DFF_155/Q_reg  ( .DIN(g8288), .SDIN(g2606), .SSEL(test_se), .CLK(CK), 
        .Q(n2994), .QN(n2502) );
  sdffs1 \DFF_154/Q_reg  ( .DIN(g6283), .SDIN(n2993), .SSEL(test_se), .CLK(CK), 
        .Q(g2606) );
  sdffs1 \DFF_153/Q_reg  ( .DIN(g7322), .SDIN(n2992), .SSEL(test_se), .CLK(CK), 
        .Q(n2993), .QN(n2555) );
  sdffs1 \DFF_152/Q_reg  ( .DIN(g11469), .SDIN(n2991), .SSEL(test_se), .CLK(CK), .Q(n2992), .QN(n1950) );
  sdffs1 \DFF_151/Q_reg  ( .DIN(g11331), .SDIN(g2603), .SSEL(test_se), .CLK(CK), .Q(n2991), .QN(n2637) );
  sdffs1 \DFF_150/Q_reg  ( .DIN(g6285), .SDIN(g4175), .SSEL(test_se), .CLK(CK), 
        .Q(g2603) );
  sdffs1 \DFF_149/Q_reg  ( .DIN(g6799), .SDIN(n2990), .SSEL(test_se), .CLK(CK), 
        .Q(g4175), .QN(n2058) );
  sdffs1 \DFF_148/Q_reg  ( .DIN(g11404), .SDIN(n2989), .SSEL(test_se), .CLK(CK), .Q(n2990), .QN(n2743) );
  sdffs1 \DFF_147/Q_reg  ( .DIN(g8426), .SDIN(n2988), .SSEL(test_se), .CLK(CK), 
        .Q(n2989), .QN(n1937) );
  sdffs1 \DFF_146/Q_reg  ( .DIN(g11635), .SDIN(n2987), .SSEL(test_se), .CLK(CK), .Q(n2988), .QN(n2809) );
  sdffs1 \DFF_145/Q_reg  ( .DIN(g6309), .SDIN(n2986), .SSEL(test_se), .CLK(CK), 
        .Q(n2987), .QN(n1971) );
  sdffs1 \DFF_143/Q_reg  ( .DIN(g11594), .SDIN(n2985), .SSEL(test_se), .CLK(CK), .Q(n2986), .QN(n2588) );
  sdffs1 \DFF_142/Q_reg  ( .DIN(g7307), .SDIN(n2984), .SSEL(test_se), .CLK(CK), 
        .Q(n2985), .QN(n2550) );
  sdffs1 \DFF_141/Q_reg  ( .DIN(g7815), .SDIN(n2983), .SSEL(test_se), .CLK(CK), 
        .Q(n2984), .QN(n2626) );
  sdffs1 \DFF_140/Q_reg  ( .DIN(g7353), .SDIN(n2982), .SSEL(test_se), .CLK(CK), 
        .Q(n2983), .QN(n2781) );
  sdffs1 \DFF_139/Q_reg  ( .DIN(g8439), .SDIN(n2981), .SSEL(test_se), .CLK(CK), 
        .Q(n2982), .QN(n2529) );
  sdffs1 \DFF_138/Q_reg  ( .DIN(g7359), .SDIN(g1217), .SSEL(test_se), .CLK(CK), 
        .Q(n2981), .QN(n2802) );
  sdffs1 \DFF_137/Q_reg  ( .DIN(g9823), .SDIN(n2980), .SSEL(test_se), .CLK(CK), 
        .Q(g1217) );
  sdffs1 \DFF_136/Q_reg  ( .DIN(g5654), .SDIN(n2979), .SSEL(test_se), .CLK(CK), 
        .Q(n2980), .QN(\DFF_136/net423 ) );
  sdffs1 \DFF_135/Q_reg  ( .DIN(g9930), .SDIN(n2978), .SSEL(test_se), .CLK(CK), 
        .Q(n2979), .QN(n1975) );
  sdffs1 \DFF_134/Q_reg  ( .DIN(g11627), .SDIN(n2977), .SSEL(test_se), .CLK(CK), .Q(n2978), .QN(n2810) );
  sdffs1 \DFF_133/Q_reg  ( .DIN(g7766), .SDIN(n2976), .SSEL(test_se), .CLK(CK), 
        .Q(n2977), .QN(n2815) );
  sdffs1 \DFF_132/Q_reg  ( .DIN(g7309), .SDIN(n2975), .SSEL(test_se), .CLK(CK), 
        .Q(n2976), .QN(n2040) );
  sdffs1 \DFF_131/Q_reg  ( .DIN(g5662), .SDIN(n2974), .SSEL(test_se), .CLK(CK), 
        .Q(n2975), .QN(n2801) );
  sdffs1 \DFF_130/Q_reg  ( .DIN(g7351), .SDIN(g2605), .SSEL(test_se), .CLK(CK), 
        .Q(n2974), .QN(n2737) );
  sdffs1 \DFF_129/Q_reg  ( .DIN(g6282), .SDIN(n2973), .SSEL(test_se), .CLK(CK), 
        .Q(g2605) );
  sdffs1 \DFF_128/Q_reg  ( .DIN(g8992), .SDIN(g4185), .SSEL(test_se), .CLK(CK), 
        .Q(n2973), .QN(n2527) );
  sdffs1 \DFF_127/Q_reg  ( .DIN(g7289), .SDIN(n2972), .SSEL(test_se), .CLK(CK), 
        .Q(g4185), .QN(n2556) );
  sdffs1 \DFF_126/Q_reg  ( .DIN(g1360), .SDIN(n2971), .SSEL(test_se), .CLK(CK), 
        .Q(n2972), .QN(\DFF_126/net413 ) );
  sdffs1 \DFF_125/Q_reg  ( .DIN(g7310), .SDIN(n2970), .SSEL(test_se), .CLK(CK), 
        .Q(n2971), .QN(n1972) );
  sdffs1 \DFF_124/Q_reg  ( .DIN(g11256), .SDIN(n2969), .SSEL(test_se), .CLK(CK), .Q(n2970), .QN(n2675) );
  sdffs1 \DFF_123/Q_reg  ( .DIN(g7767), .SDIN(g16), .SSEL(test_se), .CLK(CK), 
        .Q(n2969), .QN(n2804) );
  sdffs1 \DFF_122/Q_reg  ( .DIN(g4906), .SDIN(n2968), .SSEL(test_se), .CLK(CK), 
        .Q(g16) );
  sdffs1 \DFF_121/Q_reg  ( .DIN(g2986), .SDIN(n2967), .SSEL(test_se), .CLK(CK), 
        .Q(n2968), .QN(\DFF_121/net408 ) );
  sdffs1 \DFF_120/Q_reg  ( .DIN(g10878), .SDIN(n2966), .SSEL(test_se), .CLK(CK), .Q(n2967), .QN(n2792) );
  sdffs1 \DFF_119/Q_reg  ( .DIN(g8278), .SDIN(n2965), .SSEL(test_se), .CLK(CK), 
        .Q(n2966), .QN(n2601) );
  sdffs1 \DFF_118/Q_reg  ( .DIN(g7335), .SDIN(g632), .SSEL(test_se), .CLK(CK), 
        .Q(n2965), .QN(n2586) );
  sdffs1 \DFF_117/Q_reg  ( .DIN(g5655), .SDIN(n2964), .SSEL(test_se), .CLK(CK), 
        .Q(g632) );
  sdffs1 \DFF_116/Q_reg  ( .DIN(n2825), .SDIN(n2963), .SSEL(test_se), .CLK(CK), 
        .Q(n2964), .QN(n2732) );
  sdffs1 \DFF_115/Q_reg  ( .DIN(g7808), .SDIN(n2962), .SSEL(test_se), .CLK(CK), 
        .Q(n2963), .QN(n2652) );
  sdffs1 \DFF_114/Q_reg  ( .DIN(g11265), .SDIN(n2961), .SSEL(test_se), .CLK(CK), .Q(n2962), .QN(n2683) );
  sdffs1 \DFF_113/Q_reg  ( .DIN(g6337), .SDIN(g4173), .SSEL(test_se), .CLK(CK), 
        .Q(n2961), .QN(n1979) );
  sdffs1 \DFF_112/Q_reg  ( .DIN(g6797), .SDIN(n2960), .SSEL(test_se), .CLK(CK), 
        .Q(g4173), .QN(n2574) );
  sdffs1 \DFF_111/Q_reg  ( .DIN(g7817), .SDIN(n2959), .SSEL(test_se), .CLK(CK), 
        .Q(n2960), .QN(n2624) );
  sdffs1 \DFF_109/Q_reg  ( .DIN(g8993), .SDIN(n2958), .SSEL(test_se), .CLK(CK), 
        .Q(n2959), .QN(n2540) );
  sdffs1 \DFF_108/Q_reg  ( .DIN(g7806), .SDIN(n2957), .SSEL(test_se), .CLK(CK), 
        .Q(n2958), .QN(n2650) );
  sdffs1 \DFF_106/Q_reg  ( .DIN(g11403), .SDIN(n2956), .SSEL(test_se), .CLK(CK), .Q(n2957), .QN(n2749) );
  sdffs1 \DFF_105/Q_reg  ( .DIN(g7317), .SDIN(n2955), .SSEL(test_se), .CLK(CK), 
        .Q(n2956), .QN(n2041) );
  sdffs1 \DFF_104/Q_reg  ( .DIN(g8450), .SDIN(n2954), .SSEL(test_se), .CLK(CK), 
        .Q(n2955), .QN(n2623) );
  sdffs1 \DFF_103/Q_reg  ( .DIN(g7810), .SDIN(n2953), .SSEL(test_se), .CLK(CK), 
        .Q(n2954), .QN(n2619) );
  sdffs1 \DFF_102/Q_reg  ( .DIN(g8423), .SDIN(n2952), .SSEL(test_se), .CLK(CK), 
        .Q(n2953), .QN(n2520) );
  sdffs1 \DFF_101/Q_reg  ( .DIN(g11039), .SDIN(g2609), .SSEL(test_se), .CLK(CK), .Q(n2952), .QN(n2706) );
  sdffs1 \DFF_100/Q_reg  ( .DIN(g6253), .SDIN(g4189), .SSEL(test_se), .CLK(CK), 
        .Q(g2609) );
  sdffs1 \DFF_99/Q_reg  ( .DIN(g8437), .SDIN(n2951), .SSEL(test_se), .CLK(CK), 
        .Q(g4189), .QN(n2043) );
  sdffs1 \DFF_98/Q_reg  ( .DIN(g8440), .SDIN(n2950), .SSEL(test_se), .CLK(CK), 
        .Q(n2951), .QN(n2530) );
  sdffs1 \DFF_97/Q_reg  ( .DIN(g7328), .SDIN(n2949), .SSEL(test_se), .CLK(CK), 
        .Q(n2950), .QN(n2541) );
  sdffs1 \DFF_96/Q_reg  ( .DIN(g10881), .SDIN(n2948), .SSEL(test_se), .CLK(CK), 
        .Q(n2949), .QN(n2752) );
  sdffs1 \DFF_95/Q_reg  ( .DIN(g8444), .SDIN(n2947), .SSEL(test_se), .CLK(CK), 
        .Q(n2948), .QN(n2534) );
  sdffs1 \DFF_94/Q_reg  ( .DIN(g6808), .SDIN(n2946), .SSEL(test_se), .CLK(CK), 
        .Q(n2947), .QN(n2567) );
  sdffs1 \DFF_93/Q_reg  ( .DIN(g3007), .SDIN(n2945), .SSEL(test_se), .CLK(CK), 
        .Q(n2946), .QN(\DFF_93/net380 ) );
  sdffs1 \DFF_92/Q_reg  ( .DIN(n2819), .SDIN(g8979), .SSEL(test_se), .CLK(CK), 
        .Q(n2945), .QN(n2030) );
  sdffs1 \DFF_91/Q_reg  ( .DIN(g7779), .SDIN(n2944), .SSEL(test_se), .CLK(CK), 
        .Q(g8979), .QN(n2020) );
  sdffs1 \DFF_90/Q_reg  ( .DIN(g7332), .SDIN(g745), .SSEL(test_se), .CLK(CK), 
        .Q(n2944), .QN(n2587) );
  sdffs1 \DFF_89/Q_reg  ( .DIN(g2639), .SDIN(n2943), .SSEL(test_se), .CLK(CK), 
        .Q(g745) );
  sdffs1 \DFF_88/Q_reg  ( .DIN(g7305), .SDIN(n2942), .SSEL(test_se), .CLK(CK), 
        .Q(n2943), .QN(n2549) );
  sdffs1 \DFF_87/Q_reg  ( .DIN(g7807), .SDIN(n2941), .SSEL(test_se), .CLK(CK), 
        .Q(n2942), .QN(n2647) );
  sdffs1 \DFF_86/Q_reg  ( .DIN(g8435), .SDIN(n2940), .SSEL(test_se), .CLK(CK), 
        .Q(n2941), .QN(n2493) );
  sdffs1 \DFF_85/Q_reg  ( .DIN(g8282), .SDIN(n2939), .SSEL(test_se), .CLK(CK), 
        .Q(n2940), .QN(n2508) );
  sdffs1 \DFF_83/Q_reg  ( .DIN(g8570), .SDIN(n2938), .SSEL(test_se), .CLK(CK), 
        .Q(n2939), .QN(n2007) );
  sdffs1 \DFF_82/Q_reg  ( .DIN(g6812), .SDIN(n2937), .SSEL(test_se), .CLK(CK), 
        .Q(n2938), .QN(n2563) );
  sdffs1 \DFF_81/Q_reg  ( .DIN(g7364), .SDIN(g1957), .SSEL(test_se), .CLK(CK), 
        .Q(n2937), .QN(n2739) );
  sdffs1 \DFF_80/Q_reg  ( .DIN(g1956), .SDIN(n2936), .SSEL(test_se), .CLK(CK), 
        .Q(g1957) );
  sdffs1 \DFF_79/Q_reg  ( .DIN(g11507), .SDIN(n2935), .SSEL(test_se), .CLK(CK), 
        .Q(n2936), .QN(n2596) );
  sdffs1 \DFF_78/Q_reg  ( .DIN(g5668), .SDIN(n2934), .SSEL(test_se), .CLK(CK), 
        .Q(n2935), .QN(n2734) );
  sdffs1 \DFF_77/Q_reg  ( .DIN(g4907), .SDIN(n2933), .SSEL(test_se), .CLK(CK), 
        .Q(n2934), .QN(n2576) );
  sdffs1 \DFF_76/Q_reg  ( .DIN(g7323), .SDIN(n2932), .SSEL(test_se), .CLK(CK), 
        .Q(n2933), .QN(n1963) );
  sdffs1 \DFF_75/Q_reg  ( .DIN(g8080), .SDIN(n2931), .SSEL(test_se), .CLK(CK), 
        .Q(n2932), .QN(n2025) );
  sdffs1 \DFF_74/Q_reg  ( .DIN(g8448), .SDIN(n2930), .SSEL(test_se), .CLK(CK), 
        .Q(n2931), .QN(n2709) );
  sdffs1 \DFF_73/Q_reg  ( .DIN(g11041), .SDIN(n2929), .SSEL(test_se), .CLK(CK), 
        .Q(n2930), .QN(n2702) );
  sdffs1 \DFF_72/Q_reg  ( .DIN(g8063), .SDIN(g113), .SSEL(test_se), .CLK(CK), 
        .Q(n2929), .QN(n1981) );
  sdffs1 \DFF_71/Q_reg  ( .DIN(g7285), .SDIN(n2928), .SSEL(test_se), .CLK(CK), 
        .Q(g113) );
  sdffs1 \DFF_70/Q_reg  ( .DIN(g11508), .SDIN(n2927), .SSEL(test_se), .CLK(CK), 
        .Q(n2928), .QN(n2595) );
  sdffs1 \DFF_69/Q_reg  ( .DIN(g11038), .SDIN(g1956), .SSEL(test_se), .CLK(CK), 
        .Q(n2927), .QN(n2708) );
  sdffs1 \DFF_68/Q_reg  ( .DIN(g1955), .SDIN(n2548), .SSEL(test_se), .CLK(CK), 
        .Q(g1956) );
  sdffs1 \DFF_67/Q_reg  ( .DIN(g7311), .SDIN(n2926), .SSEL(test_se), .CLK(CK), 
        .Q(n2548) );
  sdffs1 \DFF_66/Q_reg  ( .DIN(g6836), .SDIN(n2925), .SSEL(test_se), .CLK(CK), 
        .Q(n2926), .QN(n2559) );
  sdffs1 \DFF_65/Q_reg  ( .DIN(g5649), .SDIN(n2924), .SSEL(test_se), .CLK(CK), 
        .Q(n2925), .QN(n2684) );
  sdffs1 \DFF_64/Q_reg  ( .DIN(g8065), .SDIN(g8977), .SSEL(test_se), .CLK(CK), 
        .Q(n2924), .QN(n2516) );
  sdffs1 \DFF_63/Q_reg  ( .DIN(g7777), .SDIN(g2602), .SSEL(test_se), .CLK(CK), 
        .Q(g8977), .QN(n2021) );
  sdffs1 \DFF_62/Q_reg  ( .DIN(g6284), .SDIN(n2923), .SSEL(test_se), .CLK(CK), 
        .Q(g2602) );
  sdffs1 \DFF_61/Q_reg  ( .DIN(g7292), .SDIN(n2922), .SSEL(test_se), .CLK(CK), 
        .Q(n2923), .QN(n2609) );
  sdffs1 \DFF_60/Q_reg  ( .DIN(g8429), .SDIN(n2921), .SSEL(test_se), .CLK(CK), 
        .Q(n2922), .QN(n2499) );
  sdffs1 \DFF_59/Q_reg  ( .DIN(g7814), .SDIN(n2920), .SSEL(test_se), .CLK(CK), 
        .Q(n2921), .QN(n2622) );
  sdffs1 \DFF_58/Q_reg  ( .DIN(g7302), .SDIN(n2919), .SSEL(test_se), .CLK(CK), 
        .Q(n2920), .QN(n2604) );
  sdffs1 \DFF_57/Q_reg  ( .DIN(g9344), .SDIN(n2918), .SSEL(test_se), .CLK(CK), 
        .Q(n2919), .QN(n2029) );
  sdffs1 \DFF_56/Q_reg  ( .DIN(g6811), .SDIN(n2917), .SSEL(test_se), .CLK(CK), 
        .Q(n2918), .QN(n2564) );
  sdffs1 \DFF_55/Q_reg  ( .DIN(g4182), .SDIN(n2916), .SSEL(test_se), .CLK(CK), 
        .Q(n2917), .QN(n2662) );
  sdffs1 \DFF_54/Q_reg  ( .DIN(n778), .SDIN(g3007), .SSEL(test_se), .CLK(CK), 
        .Q(n2916), .QN(n2575) );
  sdffs1 \DFF_53/Q_reg  ( .DIN(n2827), .SDIN(n2915), .SSEL(test_se), .CLK(CK), 
        .Q(g3007) );
  sdffs1 \DFF_52/Q_reg  ( .DIN(g11472), .SDIN(n2914), .SSEL(test_se), .CLK(CK), 
        .Q(n2915), .QN(n2760) );
  sdffs1 \DFF_51/Q_reg  ( .DIN(g11333), .SDIN(n2913), .SSEL(test_se), .CLK(CK), 
        .Q(n2914), .QN(n2640) );
  sdffs1 \DFF_50/Q_reg  ( .DIN(g11047), .SDIN(g8985), .SSEL(test_se), .CLK(CK), 
        .Q(n2913), .QN(n2697) );
  sdffs1 \DFF_49/Q_reg  ( .DIN(g7775), .SDIN(n2912), .SSEL(test_se), .CLK(CK), 
        .Q(g8985), .QN(n2023) );
  sdffs1 \DFF_48/Q_reg  ( .DIN(g8433), .SDIN(n2911), .SSEL(test_se), .CLK(CK), 
        .Q(n2912), .QN(n2495) );
  sdffs1 \DFF_47/Q_reg  ( .DIN(g8989), .SDIN(n2910), .SSEL(test_se), .CLK(CK), 
        .Q(n2911), .QN(n2524) );
  sdffs1 \DFF_46/Q_reg  ( .DIN(g7765), .SDIN(n2909), .SSEL(test_se), .CLK(CK), 
        .Q(n2910), .QN(n2735) );
  sdffs1 \DFF_45/Q_reg  ( .DIN(g11033), .SDIN(n2908), .SSEL(test_se), .CLK(CK), 
        .Q(n2909), .QN(n2716) );
  sdffs1 \DFF_44/Q_reg  ( .DIN(g9354), .SDIN(n2907), .SSEL(test_se), .CLK(CK), 
        .Q(n2908), .QN(n1954) );
  sdffs1 \DFF_43/Q_reg  ( .DIN(g9338), .SDIN(n2906), .SSEL(test_se), .CLK(CK), 
        .Q(n2907), .QN(n1987) );
  sdffs1 \DFF_42/Q_reg  ( .DIN(g7341), .SDIN(n2905), .SSEL(test_se), .CLK(CK), 
        .Q(n2906), .QN(n2758) );
  sdffs1 \DFF_41/Q_reg  ( .DIN(g5645), .SDIN(n2904), .SSEL(test_se), .CLK(CK), 
        .Q(n2905), .QN(n2666) );
  sdffs1 \DFF_39/Q_reg  ( .DIN(g7344), .SDIN(g4180), .SSEL(test_se), .CLK(CK), 
        .Q(n2904), .QN(n2814) );
  sdffs1 \DFF_38/Q_reg  ( .DIN(g8436), .SDIN(g757), .SSEL(test_se), .CLK(CK), 
        .Q(g4180), .QN(n2511) );
  sdffs1 \DFF_37/Q_reg  ( .DIN(n518), .SDIN(n2903), .SSEL(test_se), .CLK(CK), 
        .Q(g757) );
  sdffs1 \DFF_36/Q_reg  ( .DIN(g8987), .SDIN(n2902), .SSEL(test_se), .CLK(CK), 
        .Q(n2903), .QN(n2522) );
  sdffs1 \DFF_34/Q_reg  ( .DIN(g8447), .SDIN(n2901), .SSEL(test_se), .CLK(CK), 
        .Q(n2902), .QN(n2543) );
  sdffs1 \DFF_33/Q_reg  ( .DIN(g7325), .SDIN(n2900), .SSEL(test_se), .CLK(CK), 
        .Q(n2901), .QN(n2002) );
  sdffs1 \DFF_32/Q_reg  ( .DIN(g7290), .SDIN(n2899), .SSEL(test_se), .CLK(CK), 
        .Q(n2900), .QN(n2607) );
  sdffs1 \DFF_31/Q_reg  ( .DIN(g6815), .SDIN(g4177), .SSEL(test_se), .CLK(CK), 
        .Q(n2899), .QN(n1976) );
  sdffs1 \DFF_30/Q_reg  ( .DIN(g7785), .SDIN(n2898), .SSEL(test_se), .CLK(CK), 
        .Q(g4177), .QN(n2057) );
  sdffs1 \DFF_29/Q_reg  ( .DIN(g8079), .SDIN(n2897), .SSEL(test_se), .CLK(CK), 
        .Q(n2898), .QN(n2775) );
  sdffs1 \DFF_28/Q_reg  ( .DIN(g8279), .SDIN(n2896), .SSEL(test_se), .CLK(CK), 
        .Q(n2897), .QN(n2048) );
  sdffs1 \DFF_27/Q_reg  ( .DIN(g6805), .SDIN(n2895), .SSEL(test_se), .CLK(CK), 
        .Q(n2896), .QN(n2570) );
  sdffs1 \DFF_26/Q_reg  ( .DIN(g11037), .SDIN(g1737), .SSEL(test_se), .CLK(CK), 
        .Q(n2895), .QN(n2710) );
  sdffs1 \DFF_25/Q_reg  ( .DIN(g1736), .SDIN(n2894), .SSEL(test_se), .CLK(CK), 
        .Q(g1737) );
  sdffs1 \DFF_24/Q_reg  ( .DIN(g7330), .SDIN(n2645), .SSEL(test_se), .CLK(CK), 
        .Q(n2894), .QN(n2539) );
  sdffs1 \DFF_23/Q_reg  ( .DIN(g11182), .SDIN(n2893), .SSEL(test_se), .CLK(CK), 
        .Q(n2645) );
  sdffs1 \DFF_22/Q_reg  ( .DIN(g10774), .SDIN(g1736), .SSEL(test_se), .CLK(CK), 
        .Q(n2893), .QN(n2812) );
  sdffs1 \DFF_21/Q_reg  ( .DIN(g6846), .SDIN(n2892), .SSEL(test_se), .CLK(CK), 
        .Q(g1736) );
  sdffs1 \DFF_20/Q_reg  ( .DIN(g7356), .SDIN(n2891), .SSEL(test_se), .CLK(CK), 
        .Q(n2892), .QN(n2738) );
  sdffs1 \DFF_19/Q_reg  ( .DIN(g11439), .SDIN(n2625), .SSEL(test_se), .CLK(CK), 
        .Q(n2891), .QN(n2672) );
  sdffs1 \DFF_18/Q_reg  ( .DIN(g7816), .SDIN(n2890), .SSEL(test_se), .CLK(CK), 
        .Q(n2625) );
  sdffs1 \DFF_17/Q_reg  ( .DIN(g7354), .SDIN(n2889), .SSEL(test_se), .CLK(CK), 
        .Q(n2890), .QN(n2770) );
  sdffs1 \DFF_16/Q_reg  ( .DIN(g6810), .SDIN(n2888), .SSEL(test_se), .CLK(CK), 
        .Q(n2889), .QN(n2565) );
  sdffs1 \DFF_15/Q_reg  ( .DIN(g8432), .SDIN(n2887), .SSEL(test_se), .CLK(CK), 
        .Q(n2888), .QN(n2496) );
  sdffs1 \DFF_14/Q_reg  ( .DIN(g11471), .SDIN(n2886), .SSEL(test_se), .CLK(CK), 
        .Q(n2887), .QN(n2044) );
  sdffs1 \DFF_13/Q_reg  ( .DIN(g8572), .SDIN(n2885), .SSEL(test_se), .CLK(CK), 
        .Q(n2886), .QN(n2045) );
  sdffs1 \DFF_12/Q_reg  ( .DIN(g11467), .SDIN(n2884), .SSEL(test_se), .CLK(CK), 
        .Q(n2885), .QN(n1930) );
  sdffs1 \DFF_11/Q_reg  ( .DIN(g9343), .SDIN(n2883), .SSEL(test_se), .CLK(CK), 
        .Q(n2884), .QN(n1958) );
  sdffs1 \DFF_10/Q_reg  ( .DIN(g7349), .SDIN(n2882), .SSEL(test_se), .CLK(CK), 
        .Q(n2883), .QN(n2759) );
  sdffs1 \DFF_9/Q_reg  ( .DIN(g5663), .SDIN(n2881), .SSEL(test_se), .CLK(CK), 
        .Q(n2882), .QN(n2791) );
  sdffs1 \DFF_7/Q_reg  ( .DIN(g6304), .SDIN(n2880), .SSEL(test_se), .CLK(CK), 
        .Q(n2881), .QN(n1988) );
  sdffs1 \DFF_6/Q_reg  ( .DIN(g9345), .SDIN(n2879), .SSEL(test_se), .CLK(CK), 
        .Q(n2880), .QN(n1955) );
  sdffs1 \DFF_5/Q_reg  ( .DIN(g7315), .SDIN(n2878), .SSEL(test_se), .CLK(CK), 
        .Q(n2879), .QN(n2001) );
  sdffs1 \DFF_4/Q_reg  ( .DIN(g8272), .SDIN(n2877), .SSEL(test_se), .CLK(CK), 
        .Q(n2878), .QN(n2789) );
  sdffs1 \DFF_3/Q_reg  ( .DIN(g11257), .SDIN(n2876), .SSEL(test_se), .CLK(CK), 
        .Q(n2877), .QN(n2677) );
  sdffs1 \DFF_2/Q_reg  ( .DIN(g5644), .SDIN(n2875), .SSEL(test_se), .CLK(CK), 
        .Q(n2876), .QN(n2668) );
  sdffs1 \DFF_1/Q_reg  ( .DIN(g9349), .SDIN(n2874), .SSEL(test_se), .CLK(CK), 
        .Q(n2875), .QN(n1935) );
  sdffs1 \DFF_0/Q_reg  ( .DIN(g5660), .SDIN(test_si), .SSEL(test_se), .CLK(CK), 
        .Q(n2874), .QN(n2617) );
  i1s1 trig50_0U1 ( .DIN(trig50_0n1), .Q(Trigger_en0_0) );
  nnd2s1 trig50_0U2 ( .DIN1(trig50_0n2), .DIN2(trig50_0n3), .Q(trig50_0n1) );
  nor5s1 trig50_0U3 ( .DIN1(n592), .DIN2(trig50_0n4), .DIN3(n1466), .DIN4(n1798), .DIN5(n1698),         .Q(trig50_0n3) );
  or2s1 trig50_0U4 ( .DIN1(n762), .DIN2(n632), .Q(trig50_0n4) );
  and4s1 trig50_0U5 ( .DIN1(n920), .DIN2(n880), .DIN3(trig50_0n5), .DIN4(n1107), .Q(trig50_0n2) );
  nor2s1 trig50_0U6 ( .DIN1(n1209), .DIN2(n1045), .Q(trig50_0n5) );
  dffs2 troj12_0counter_reg_0_ ( .DIN(troj12_0n10), .CLK(CK), .Q(troj12_0counter_0_) );
  dffles2 troj12_0counter_reg_1_ ( .DIN(troj12_0N1), .EB(troj12_0n9), .CLK(CK), .QN(troj12_0n6) );
  dffles2 troj12_0counter_reg_2_ ( .DIN(troj12_0N2), .EB(troj12_0n9), .CLK(CK), .QN(troj12_0n8) );
  dffles2 troj12_0counter_reg_3_ ( .DIN(troj12_0N3), .EB(troj12_0n9), .CLK(CK), .QN(troj12_0n7) );
  dffs2 troj12_0Trojan_out0_reg ( .DIN(troj12_0N6), .CLK(CK), .Q(Trojan_out0) );
  hi1s1 troj12_0U3 ( .DIN(Trigger_en0_0), .Q(troj12_0n9) );
  xnr2s1 troj12_0U4 ( .DIN1(troj12_0n1), .DIN2(Trigger_en0_0), .Q(troj12_0n10) );
  and3s1 troj12_0U5 ( .DIN1(troj12_0n2), .DIN2(troj12_0n3), .DIN3(troj12_0n4), .Q(troj12_0N6) );
  xnr2s1 troj12_0U6 ( .DIN1(troj12_0n5), .DIN2(troj12_0n3), .Q(troj12_0N3) );
  hi1s1 troj12_0U7 ( .DIN(troj12_0n7), .Q(troj12_0n3) );
  nnd2s1 troj12_0U8 ( .DIN1(troj12_0n4), .DIN2(troj12_0n2), .Q(troj12_0n5) );
  hi1s1 troj12_0U9 ( .DIN(troj12_0n8), .Q(troj12_0n2) );
  xnr2s1 troj12_0U10 ( .DIN1(troj12_0n8), .DIN2(troj12_0n4), .Q(troj12_0N2) );
  nor2s1 troj12_0U11 ( .DIN1(troj12_0n1), .DIN2(troj12_0n6), .Q(troj12_0n4) );
  hi1s1 troj12_0U12 ( .DIN(troj12_0counter_0_), .Q(troj12_0n1) );
  xnr2s1 troj12_0U13 ( .DIN1(troj12_0counter_0_), .DIN2(troj12_0n6), .Q(troj12_0N1) );
    xor2s1 trojan12_0  (.DIN1(tempn1458), .DIN2(Trojan_out0), .Q(n1458) );

endmodule

