
module c2670 ( N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, 
    N21, N22, N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, 
    N40, N43, N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, 
    N61, N62, N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, 
    N78, N79, N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, 
    N95, N96, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, 
    N112, N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, 
    N126, N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, 
    N140, N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, 
    N253, N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, 
    N287, N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, 
    N328, N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, 
    N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, 
    N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, 
    N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, 
    N172_I, N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I, 
    N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, 
    N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, 
    N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, 
    N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, 
    N217_I, N218_I, N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, 
    N489, N490, N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, 
    N1269, N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, 
    N1969, N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, 
    N2387, N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, 
    N2971, N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, 
    N3881, N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, 
    N150_O, N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, 
    N159_O, N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, 
    N168_O, N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, 
    N177_O, N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, 
    N186_O, N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, 
    N195_O, N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, 
    N204_O, N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, 
    N213_O, N214_O, N215_O, N216_O, N217_O, N218_O );

input  N1, N2, N3, N4, N5, N6, N7, N8, N11, N14, N15, N16, N19, N20, N21, N22, 
    N23, N24, N25, N26, N27, N28, N29, N32, N33, N34, N35, N36, N37, N40, N43, 
    N44, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N60, N61, N62, 
    N63, N64, N65, N66, N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, 
    N80, N81, N82, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, 
    N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N111, N112, 
    N113, N114, N115, N116, N117, N118, N119, N120, N123, N124, N125, N126, 
    N127, N128, N129, N130, N131, N132, N135, N136, N137, N138, N139, N140, 
    N141, N142, N219, N224, N227, N230, N231, N234, N237, N241, N246, N253, 
    N256, N259, N262, N263, N266, N269, N272, N275, N278, N281, N284, N287, 
    N290, N294, N297, N301, N305, N309, N313, N316, N319, N322, N325, N328, 
    N331, N334, N337, N340, N343, N346, N349, N352, N355, N143_I, N144_I, 
    N145_I, N146_I, N147_I, N148_I, N149_I, N150_I, N151_I, N152_I, N153_I, 
    N154_I, N155_I, N156_I, N157_I, N158_I, N159_I, N160_I, N161_I, N162_I, 
    N163_I, N164_I, N165_I, N166_I, N167_I, N168_I, N169_I, N170_I, N171_I, 
    N172_I, N173_I, N174_I, N175_I, N176_I, N177_I, N178_I, N179_I, N180_I, 
    N181_I, N182_I, N183_I, N184_I, N185_I, N186_I, N187_I, N188_I, N189_I, 
    N190_I, N191_I, N192_I, N193_I, N194_I, N195_I, N196_I, N197_I, N198_I, 
    N199_I, N200_I, N201_I, N202_I, N203_I, N204_I, N205_I, N206_I, N207_I, 
    N208_I, N209_I, N210_I, N211_I, N212_I, N213_I, N214_I, N215_I, N216_I, 
    N217_I, N218_I;

output N398, N400, N401, N419, N420, N456, N457, N458, N487, N488, N489, N490, 
    N491, N492, N493, N494, N792, N799, N805, N1026, N1028, N1029, N1269, 
    N1277, N1448, N1726, N1816, N1817, N1818, N1819, N1820, N1821, N1969, 
    N1970, N1971, N2010, N2012, N2014, N2016, N2018, N2020, N2022, N2387, 
    N2388, N2389, N2390, N2496, N2643, N2644, N2891, N2925, N2970, N2971, 
    N3038, N3079, N3546, N3671, N3803, N3804, N3809, N3851, N3875, N3881, 
    N3882, N143_O, N144_O, N145_O, N146_O, N147_O, N148_O, N149_O, N150_O, 
    N151_O, N152_O, N153_O, N154_O, N155_O, N156_O, N157_O, N158_O, N159_O, 
    N160_O, N161_O, N162_O, N163_O, N164_O, N165_O, N166_O, N167_O, N168_O, 
    N169_O, N170_O, N171_O, N172_O, N173_O, N174_O, N175_O, N176_O, N177_O, 
    N178_O, N179_O, N180_O, N181_O, N182_O, N183_O, N184_O, N185_O, N186_O, 
    N187_O, N188_O, N189_O, N190_O, N191_O, N192_O, N193_O, N194_O, N195_O, 
    N196_O, N197_O, N198_O, N199_O, N200_O, N201_O, N202_O, N203_O, N204_O, 
    N205_O, N206_O, N207_O, N208_O, N209_O, N210_O, N211_O, N212_O, N213_O, 
    N214_O, N215_O, N216_O, N217_O, N218_O;

    wire n279, n280, n281, n282, n283, n284, n285, n286, n288, n289, n290, 
        n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
        n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
        n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
        n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
        n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
        n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
        n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
        n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
        n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
        n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
        n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
        n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
        n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
        n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
        n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
        n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
        n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
        n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
        n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
        n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
        n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
        n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
        n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
        n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
        n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
        n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
        n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
        n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
        n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
        n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
        n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
        n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
        n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
        n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
        n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
        n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
        n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
        n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
        n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
        n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
        n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
        n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
        n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
        n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
        n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
        n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
        n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
        n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
        n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, 
        n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, 
        n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, 
        n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
        n915;


wire Trigger_en59_0,  troj59_0n1,  troj59_0n2,  troj59_0n3,  troj59_0n4,  troj59_0n5,  troj59_0n6,  tempn391;

    assign N398 = N219;
    assign N400 = N219;
    assign N401 = N219;
    assign N419 = N253;
    assign N420 = N253;
    assign N456 = N290;
    assign N457 = N290;
    assign N458 = N290;
    assign N805 = N219;
    assign N2388 = N2387;
    assign N2390 = N2389;
    assign N2644 = N2643;
    assign N3804 = N3803;
    assign N3875 = 1'b0;
    assign N143_O = N143_I;
    assign N144_O = N144_I;
    assign N145_O = N145_I;
    assign N146_O = N146_I;
    assign N147_O = N147_I;
    assign N148_O = N148_I;
    assign N149_O = N149_I;
    assign N150_O = N150_I;
    assign N151_O = N151_I;
    assign N152_O = N152_I;
    assign N153_O = N153_I;
    assign N154_O = N154_I;
    assign N155_O = N155_I;
    assign N156_O = N156_I;
    assign N157_O = N157_I;
    assign N158_O = N158_I;
    assign N159_O = N159_I;
    assign N160_O = N160_I;
    assign N161_O = N161_I;
    assign N162_O = N162_I;
    assign N163_O = N163_I;
    assign N164_O = N164_I;
    assign N165_O = N165_I;
    assign N166_O = N166_I;
    assign N167_O = N167_I;
    assign N168_O = N168_I;
    assign N169_O = N169_I;
    assign N170_O = N170_I;
    assign N171_O = N171_I;
    assign N172_O = N172_I;
    assign N173_O = N173_I;
    assign N174_O = N174_I;
    assign N175_O = N175_I;
    assign N176_O = N176_I;
    assign N177_O = N177_I;
    assign N178_O = N178_I;
    assign N179_O = N179_I;
    assign N180_O = N180_I;
    assign N181_O = N181_I;
    assign N182_O = N182_I;
    assign N183_O = N183_I;
    assign N184_O = N184_I;
    assign N185_O = N185_I;
    assign N186_O = N186_I;
    assign N187_O = N187_I;
    assign N188_O = N188_I;
    assign N189_O = N189_I;
    assign N190_O = N190_I;
    assign N191_O = N191_I;
    assign N192_O = N192_I;
    assign N193_O = N193_I;
    assign N194_O = N194_I;
    assign N195_O = N195_I;
    assign N196_O = N196_I;
    assign N197_O = N197_I;
    assign N198_O = N198_I;
    assign N199_O = N199_I;
    assign N200_O = N200_I;
    assign N201_O = N201_I;
    assign N202_O = N202_I;
    assign N203_O = N203_I;
    assign N204_O = N204_I;
    assign N205_O = N205_I;
    assign N206_O = N206_I;
    assign N207_O = N207_I;
    assign N208_O = N208_I;
    assign N209_O = N209_I;
    assign N210_O = N210_I;
    assign N211_O = N211_I;
    assign N212_O = N212_I;
    assign N213_O = N213_I;
    assign N214_O = N214_I;
    assign N215_O = N215_I;
    assign N216_O = N216_I;
    assign N217_O = N217_I;
    assign N218_O = N218_I;
    nor2s1 U1 ( .Q(N3038), .DIN1(n279), .DIN2(n280) );
    hi1s1 U2 ( .Q(N2022), .DIN(n281) );
    hi1s1 U3 ( .Q(N2020), .DIN(n282) );
    hi1s1 U4 ( .Q(N2018), .DIN(n283) );
    hi1s1 U5 ( .Q(N2016), .DIN(N1819) );
    hi1s1 U6 ( .Q(N2014), .DIN(N1820) );
    hi1s1 U7 ( .Q(N2012), .DIN(N1821) );
    hi1s1 U8 ( .Q(N2010), .DIN(n284) );
    nor2s1 U9 ( .Q(N3881), .DIN1(n285), .DIN2(n286) );
    nnd2s1 U11 ( .Q(N3851), .DIN1(n288), .DIN2(n289) );
    hi1s1 U12 ( .Q(N3079), .DIN(N3038) );
    nnd2s1 U13 ( .Q(N2891), .DIN1(n290), .DIN2(n291) );
    nnd2s1 U14 ( .Q(N1971), .DIN1(n292), .DIN2(n293) );
    nnd2s1 U15 ( .Q(N1970), .DIN1(N36), .DIN2(n292) );
    nnd2s1 U16 ( .Q(N1969), .DIN1(N241), .DIN2(n294) );
    nor2s1 U17 ( .Q(N1277), .DIN1(n295), .DIN2(n296) );
    nnd2s1 U18 ( .Q(N1029), .DIN1(N231), .DIN2(n297) );
    nnd2s1 U19 ( .Q(N1269), .DIN1(N325), .DIN2(n297) );
    nnd2s1 U20 ( .Q(N792), .DIN1(n298), .DIN2(n299) );
    nnd2s1 U21 ( .Q(N1028), .DIN1(N7), .DIN2(N237) );
    hi1s1 U22 ( .Q(N494), .DIN(N108) );
    hi1s1 U23 ( .Q(N493), .DIN(N57) );
    hi1s1 U24 ( .Q(N492), .DIN(N120) );
    hi1s1 U25 ( .Q(N491), .DIN(N69) );
    hi1s1 U26 ( .Q(N490), .DIN(N96) );
    hi1s1 U27 ( .Q(N489), .DIN(N82) );
    hi1s1 U28 ( .Q(N488), .DIN(N132) );
    hi1s1 U29 ( .Q(N487), .DIN(N44) );
    nnd2s1 U30 ( .Q(N799), .DIN1(N237), .DIN2(n300) );
    nor2s1 U31 ( .Q(n301), .DIN1(n302), .DIN2(n303) );
    nor2s1 U32 ( .Q(N1816), .DIN1(n304), .DIN2(n305) );
    nor2s1 U33 ( .Q(N1817), .DIN1(n306), .DIN2(n307) );
    nor2s1 U34 ( .Q(n308), .DIN1(n309), .DIN2(n310) );
    nor2s1 U35 ( .Q(n311), .DIN1(n312), .DIN2(n313) );
    nor2s1 U36 ( .Q(n314), .DIN1(n315), .DIN2(n316) );
    nor2s1 U37 ( .Q(n317), .DIN1(n318), .DIN2(n319) );
    nor2s1 U38 ( .Q(n320), .DIN1(n321), .DIN2(n322) );
    nor2s1 U39 ( .Q(N1818), .DIN1(n323), .DIN2(n324) );
    nor2s1 U40 ( .Q(N1820), .DIN1(n325), .DIN2(n326) );
    nor2s1 U41 ( .Q(N1821), .DIN1(n327), .DIN2(n328) );
    nor2s1 U42 ( .Q(n329), .DIN1(n330), .DIN2(n331) );
    nor2s1 U43 ( .Q(n294), .DIN1(n332), .DIN2(n333) );
    nor2s1 U44 ( .Q(n284), .DIN1(n334), .DIN2(n335) );
    nor2s1 U45 ( .Q(n336), .DIN1(n337), .DIN2(n338) );
    nor2s1 U46 ( .Q(n281), .DIN1(n339), .DIN2(n340) );
    nor2s1 U47 ( .Q(n282), .DIN1(n341), .DIN2(n342) );
    nor2s1 U48 ( .Q(n283), .DIN1(n343), .DIN2(n344) );
    nor2s1 U49 ( .Q(N1819), .DIN1(n345), .DIN2(n346) );
    nor2s1 U50 ( .Q(n347), .DIN1(N262), .DIN2(N1818) );
    nor2s1 U51 ( .Q(n348), .DIN1(n349), .DIN2(n350) );
    nor2s1 U52 ( .Q(n351), .DIN1(n352), .DIN2(n353) );
    nor2s1 U53 ( .Q(n354), .DIN1(n352), .DIN2(n355) );
    nor2s1 U54 ( .Q(n356), .DIN1(n357), .DIN2(n358) );
    nnd2s1 U55 ( .Q(n359), .DIN1(n360), .DIN2(n361) );
    nor2s1 U56 ( .Q(n362), .DIN1(N1821), .DIN2(n363) );
    nnd2s1 U57 ( .Q(n364), .DIN1(n365), .DIN2(n366) );
    nor2s1 U58 ( .Q(n367), .DIN1(n368), .DIN2(n369) );
    nor2s1 U59 ( .Q(n370), .DIN1(n371), .DIN2(n372) );
    nor2s1 U60 ( .Q(n373), .DIN1(n367), .DIN2(n370) );
    nor2s1 U61 ( .Q(n374), .DIN1(n352), .DIN2(n375) );
    nor2s1 U62 ( .Q(n376), .DIN1(n354), .DIN2(n373) );
    nor2s1 U63 ( .Q(n377), .DIN1(n374), .DIN2(n376) );
    nor2s1 U64 ( .Q(n378), .DIN1(n352), .DIN2(n379) );
    nor2s1 U65 ( .Q(n380), .DIN1(n351), .DIN2(n377) );
    nor2s1 U66 ( .Q(n381), .DIN1(n378), .DIN2(n380) );
    nor2s1 U67 ( .Q(n382), .DIN1(n383), .DIN2(n384) );
    nor2s1 U68 ( .Q(n385), .DIN1(n386), .DIN2(n387) );
    nor2s1 U69 ( .Q(n388), .DIN1(n389), .DIN2(n390) );
    nor2s1 U70 ( .Q( tempn391 ), .DIN1(n392), .DIN2(n393) );
    nor2s1 U71 ( .Q(n394), .DIN1(n395), .DIN2(n396) );
    nnd2s1 U72 ( .Q(N2496), .DIN1(n336), .DIN2(n397) );
    nor2s1 U73 ( .Q(n398), .DIN1(n284), .DIN2(n359) );
    nor2s1 U74 ( .Q(n371), .DIN1(n356), .DIN2(n394) );
    hi1s1 U75 ( .Q(n399), .DIN(n336) );
    hi1s1 U76 ( .Q(n400), .DIN(N301) );
    hi1s1 U77 ( .Q(n401), .DIN(N297) );
    hi1s1 U78 ( .Q(n402), .DIN(N309) );
    hi1s1 U79 ( .Q(n403), .DIN(N305) );
    nor2s1 U80 ( .Q(n404), .DIN1(N319), .DIN2(N322) );
    hi1s1 U81 ( .Q(n405), .DIN(N319) );
    nor2s1 U82 ( .Q(n406), .DIN1(n405), .DIN2(N322) );
    nor2s1 U83 ( .Q(n407), .DIN1(n408), .DIN2(N319) );
    nor2s1 U84 ( .Q(n409), .DIN1(n408), .DIN2(n405) );
    hi1s1 U85 ( .Q(n410), .DIN(n314) );
    hi1s1 U86 ( .Q(n411), .DIN(n317) );
    hi1s1 U87 ( .Q(n412), .DIN(N1816) );
    hi1s1 U88 ( .Q(n413), .DIN(n308) );
    nor2s1 U89 ( .Q(n414), .DIN1(N227), .DIN2(N234) );
    hi1s1 U90 ( .Q(n415), .DIN(N227) );
    nor2s1 U91 ( .Q(n416), .DIN1(n417), .DIN2(n415) );
    nor2s1 U92 ( .Q(n418), .DIN1(n415), .DIN2(N234) );
    nor2s1 U93 ( .Q(n419), .DIN1(n417), .DIN2(N227) );
    hi1s1 U94 ( .Q(n420), .DIN(n329) );
    hi1s1 U95 ( .Q(n421), .DIN(n294) );
    hi1s1 U96 ( .Q(n422), .DIN(N294) );
    hi1s1 U97 ( .Q(n423), .DIN(N275) );
    hi1s1 U98 ( .Q(n424), .DIN(N266) );
    hi1s1 U99 ( .Q(n425), .DIN(N284) );
    hi1s1 U100 ( .Q(n426), .DIN(N287) );
    hi1s1 U101 ( .Q(n427), .DIN(N278) );
    hi1s1 U102 ( .Q(n428), .DIN(N281) );
    hi1s1 U103 ( .Q(n429), .DIN(N263) );
    nnd2s1 U104 ( .Q(n430), .DIN1(n431), .DIN2(n432) );
    nnd2s1 U105 ( .Q(n349), .DIN1(n433), .DIN2(N40) );
    hi1s1 U106 ( .Q(n357), .DIN(N8) );
    nnd2s1 U107 ( .Q(n352), .DIN1(N8), .DIN2(n434) );
    nnd2s1 U108 ( .Q(n369), .DIN1(n435), .DIN2(N8) );
    nor2s1 U109 ( .Q(n368), .DIN1(n357), .DIN2(N1819) );
    nnd2s1 U110 ( .Q(n436), .DIN1(n437), .DIN2(n294) );
    nor2s1 U111 ( .Q(n395), .DIN1(n357), .DIN2(N1820) );
    nor2s1 U112 ( .Q(n438), .DIN1(n399), .DIN2(N230) );
    nor2s1 U113 ( .Q(n292), .DIN1(n439), .DIN2(n440) );
    hi1s1 U114 ( .Q(n441), .DIN(N241) );
    nnd2s1 U115 ( .Q(n296), .DIN1(n442), .DIN2(n443) );
    nnd2s1 U116 ( .Q(n295), .DIN1(n444), .DIN2(n445) );
    nor2s1 U117 ( .Q(n446), .DIN1(n447), .DIN2(n448) );
    nor2s1 U118 ( .Q(n449), .DIN1(n450), .DIN2(n451) );
    nnd2s1 U119 ( .Q(N2971), .DIN1(n452), .DIN2(n453) );
    nnd2s1 U120 ( .Q(n454), .DIN1(n455), .DIN2(n456) );
    nnd2s1 U121 ( .Q(n457), .DIN1(n458), .DIN2(n459) );
    nnd2s1 U122 ( .Q(n460), .DIN1(n461), .DIN2(n462) );
    nnd2s1 U123 ( .Q(n463), .DIN1(n464), .DIN2(n465) );
    nnd2s1 U124 ( .Q(n466), .DIN1(n467), .DIN2(n468) );
    nnd2s1 U125 ( .Q(n469), .DIN1(n470), .DIN2(n471) );
    nnd2s1 U126 ( .Q(n472), .DIN1(n473), .DIN2(n474) );
    nnd2s1 U127 ( .Q(n475), .DIN1(n476), .DIN2(n477) );
    nnd2s1 U128 ( .Q(n478), .DIN1(n375), .DIN2(n355) );
    nnd2s1 U129 ( .Q(n479), .DIN1(n480), .DIN2(n481) );
    nnd2s1 U130 ( .Q(n482), .DIN1(n483), .DIN2(n350) );
    nnd2s1 U131 ( .Q(n484), .DIN1(n379), .DIN2(n353) );
    nnd2s1 U132 ( .Q(n363), .DIN1(n485), .DIN2(n486) );
    nnd2s1 U133 ( .Q(n358), .DIN1(n487), .DIN2(n488) );
    nnd2s1 U134 ( .Q(N3803), .DIN1(n489), .DIN2(n490) );
    nnd2s1 U135 ( .Q(n491), .DIN1(n492), .DIN2(n493) );
    nnd2s1 U136 ( .Q(N2643), .DIN1(n494), .DIN2(n495) );
    nnd2s1 U137 ( .Q(N2389), .DIN1(n496), .DIN2(n497) );
    nnd2s1 U138 ( .Q(N2387), .DIN1(n498), .DIN2(n499) );
    nnd2s1 U139 ( .Q(n500), .DIN1(N2), .DIN2(N15) );
    nor2s1 U140 ( .Q(n299), .DIN1(n400), .DIN2(n401) );
    nor2s1 U141 ( .Q(n298), .DIN1(n402), .DIN2(n403) );
    nnd2s1 U142 ( .Q(n312), .DIN1(n501), .DIN2(n502) );
    nnd2s1 U143 ( .Q(n313), .DIN1(n503), .DIN2(n504) );
    nnd2s1 U144 ( .Q(n315), .DIN1(n505), .DIN2(n506) );
    nnd2s1 U145 ( .Q(n316), .DIN1(n507), .DIN2(n508) );
    nnd2s1 U146 ( .Q(n318), .DIN1(n509), .DIN2(n510) );
    nnd2s1 U147 ( .Q(n319), .DIN1(n511), .DIN2(n512) );
    nnd2s1 U148 ( .Q(n302), .DIN1(n513), .DIN2(n514) );
    nnd2s1 U149 ( .Q(n303), .DIN1(n515), .DIN2(n516) );
    nnd2s1 U150 ( .Q(n304), .DIN1(n517), .DIN2(n518) );
    nnd2s1 U151 ( .Q(n305), .DIN1(n519), .DIN2(n520) );
    nnd2s1 U152 ( .Q(n306), .DIN1(n521), .DIN2(n522) );
    nnd2s1 U153 ( .Q(n307), .DIN1(n523), .DIN2(n524) );
    nnd2s1 U154 ( .Q(n309), .DIN1(n525), .DIN2(n526) );
    nnd2s1 U155 ( .Q(n310), .DIN1(n527), .DIN2(n528) );
    nnd2s1 U156 ( .Q(n321), .DIN1(n529), .DIN2(n530) );
    nnd2s1 U157 ( .Q(n322), .DIN1(n531), .DIN2(n532) );
    nnd2s1 U158 ( .Q(n323), .DIN1(n533), .DIN2(n534) );
    nnd2s1 U159 ( .Q(n324), .DIN1(n535), .DIN2(n536) );
    nnd2s1 U160 ( .Q(n537), .DIN1(n538), .DIN2(n539) );
    nor2s1 U161 ( .Q(n540), .DIN1(n541), .DIN2(n542) );
    nnd2s1 U162 ( .Q(n543), .DIN1(n544), .DIN2(n545) );
    nor2s1 U163 ( .Q(n546), .DIN1(n547), .DIN2(n548) );
    nor2s1 U164 ( .Q(n549), .DIN1(n550), .DIN2(n551) );
    nnd2s1 U165 ( .Q(n552), .DIN1(n553), .DIN2(n554) );
    nnd2s1 U166 ( .Q(n325), .DIN1(n555), .DIN2(n556) );
    nnd2s1 U167 ( .Q(n326), .DIN1(n557), .DIN2(n558) );
    nnd2s1 U168 ( .Q(n327), .DIN1(n559), .DIN2(n560) );
    nnd2s1 U169 ( .Q(n328), .DIN1(n561), .DIN2(n562) );
    nnd2s1 U170 ( .Q(n339), .DIN1(n563), .DIN2(n564) );
    nnd2s1 U171 ( .Q(n340), .DIN1(n565), .DIN2(n566) );
    nnd2s1 U172 ( .Q(n341), .DIN1(n567), .DIN2(n568) );
    nnd2s1 U173 ( .Q(n342), .DIN1(n569), .DIN2(n570) );
    nnd2s1 U174 ( .Q(n343), .DIN1(n571), .DIN2(n572) );
    nnd2s1 U175 ( .Q(n344), .DIN1(n573), .DIN2(n574) );
    nnd2s1 U176 ( .Q(n345), .DIN1(n575), .DIN2(n576) );
    nnd2s1 U177 ( .Q(n346), .DIN1(n577), .DIN2(n578) );
    nnd2s1 U178 ( .Q(n330), .DIN1(n579), .DIN2(n580) );
    nnd2s1 U179 ( .Q(n331), .DIN1(n581), .DIN2(n582) );
    nnd2s1 U180 ( .Q(n332), .DIN1(n583), .DIN2(n584) );
    nnd2s1 U181 ( .Q(n333), .DIN1(n585), .DIN2(n586) );
    nnd2s1 U182 ( .Q(n334), .DIN1(n587), .DIN2(n588) );
    nnd2s1 U183 ( .Q(n335), .DIN1(n589), .DIN2(n590) );
    nnd2s1 U184 ( .Q(n337), .DIN1(n591), .DIN2(n592) );
    nnd2s1 U185 ( .Q(n338), .DIN1(n593), .DIN2(n594) );
    nnd2s1 U186 ( .Q(n595), .DIN1(n596), .DIN2(n597) );
    nnd2s1 U187 ( .Q(n598), .DIN1(n599), .DIN2(n600) );
    nnd2s1 U188 ( .Q(n601), .DIN1(n602), .DIN2(n603) );
    nor2s1 U189 ( .Q(n604), .DIN1(n605), .DIN2(n606) );
    nnd2s1 U190 ( .Q(n607), .DIN1(n608), .DIN2(n609) );
    nor2s1 U191 ( .Q(n610), .DIN1(n611), .DIN2(n612) );
    nor2s1 U192 ( .Q(n613), .DIN1(n614), .DIN2(n615) );
    nnd2s1 U193 ( .Q(n616), .DIN1(n617), .DIN2(n618) );
    nnd2s1 U194 ( .Q(n619), .DIN1(n620), .DIN2(n621) );
    nnd2s1 U195 ( .Q(n622), .DIN1(n623), .DIN2(n624) );
    nnd2s1 U196 ( .Q(n625), .DIN1(n626), .DIN2(n627) );
    nor2s1 U197 ( .Q(n628), .DIN1(n629), .DIN2(n630) );
    nnd2s1 U198 ( .Q(n631), .DIN1(n632), .DIN2(n633) );
    nnd2s1 U199 ( .Q(n634), .DIN1(n635), .DIN2(n636) );
    nnd2s1 U200 ( .Q(n637), .DIN1(n638), .DIN2(n639) );
    nnd2s1 U201 ( .Q(n640), .DIN1(n641), .DIN2(n642) );
    nnd2s1 U202 ( .Q(n643), .DIN1(n644), .DIN2(n645) );
    nnd2s1 U203 ( .Q(n646), .DIN1(n647), .DIN2(n648) );
    nor2s1 U204 ( .Q(n649), .DIN1(n650), .DIN2(n651) );
    nor2s1 U205 ( .Q(n652), .DIN1(n653), .DIN2(n654) );
    nor2s1 U206 ( .Q(n443), .DIN1(N490), .DIN2(N489) );
    nor2s1 U207 ( .Q(n442), .DIN1(N488), .DIN2(N487) );
    nor2s1 U208 ( .Q(n445), .DIN1(N494), .DIN2(N493) );
    nor2s1 U209 ( .Q(n444), .DIN1(N492), .DIN2(N491) );
    nor2s1 U210 ( .Q(n655), .DIN1(N3809), .DIN2(N3671) );
    nnd2s1 U211 ( .Q(n286), .DIN1(n656), .DIN2(n655) );
    nor2s1 U212 ( .Q(n657), .DIN1(N2971), .DIN2(N2970) );
    nnd2s1 U213 ( .Q(n285), .DIN1(N1726), .DIN2(n657) );
    nor2s1 U214 ( .Q(n433), .DIN1(n347), .DIN2(n412) );
    nor2s1 U215 ( .Q(n658), .DIN1(N294), .DIN2(n411) );
    nor2s1 U216 ( .Q(n659), .DIN1(n317), .DIN2(n422) );
    nor2s1 U217 ( .Q(n660), .DIN1(n314), .DIN2(n426) );
    nor2s1 U218 ( .Q(n661), .DIN1(n308), .DIN2(n425) );
    nnd2s1 U219 ( .Q(n662), .DIN1(N1816), .DIN2(N40) );
    nor2s1 U220 ( .Q(n663), .DIN1(n362), .DIN2(n398) );
    nnd2s1 U221 ( .Q(n372), .DIN1(n664), .DIN2(n665) );
    nnd2s1 U222 ( .Q(n666), .DIN1(n667), .DIN2(n668) );
    nor2s1 U223 ( .Q(n669), .DIN1(n348), .DIN2(n381) );
    nor2s1 U224 ( .Q(n670), .DIN1(N2022), .DIN2(N281) );
    nnd2s1 U225 ( .Q(n671), .DIN1(n672), .DIN2(n673) );
    nnd2s1 U226 ( .Q(n674), .DIN1(n675), .DIN2(n676) );
    nor2s1 U227 ( .Q(n677), .DIN1(n678), .DIN2(n679) );
    nor2s1 U228 ( .Q(n680), .DIN1(n681), .DIN2(n682) );
    nnd2s1 U229 ( .Q(n386), .DIN1(n680), .DIN2(n677) );
    nor2s1 U230 ( .Q(n683), .DIN1(n684), .DIN2(n685) );
    nnd2s1 U231 ( .Q(n387), .DIN1(n683), .DIN2(N28) );
    nor2s1 U232 ( .Q(n686), .DIN1(n301), .DIN2(n454) );
    nor2s1 U233 ( .Q(n687), .DIN1(n457), .DIN2(n460) );
    nnd2s1 U234 ( .Q(n383), .DIN1(n687), .DIN2(n686) );
    nor2s1 U235 ( .Q(n688), .DIN1(n463), .DIN2(n466) );
    nnd2s1 U236 ( .Q(n384), .DIN1(n688), .DIN2(n689) );
    nnd2s1 U237 ( .Q(n690), .DIN1(n691), .DIN2(n692) );
    nor2s1 U238 ( .Q(n693), .DIN1(n694), .DIN2(n690) );
    nor2s1 U239 ( .Q(n695), .DIN1(n696), .DIN2(n697) );
    nnd2s1 U240 ( .Q(n392), .DIN1(n695), .DIN2(n693) );
    nor2s1 U241 ( .Q(n698), .DIN1(n699), .DIN2(n700) );
    nor2s1 U242 ( .Q(n701), .DIN1(n702), .DIN2(n703) );
    nnd2s1 U243 ( .Q(n393), .DIN1(n701), .DIN2(n698) );
    nnd2s1 U244 ( .Q(n704), .DIN1(n705), .DIN2(n706) );
    nor2s1 U245 ( .Q(n707), .DIN1(n469), .DIN2(n704) );
    nor2s1 U246 ( .Q(n708), .DIN1(n472), .DIN2(n475) );
    nnd2s1 U247 ( .Q(n389), .DIN1(n708), .DIN2(n707) );
    nor2s1 U248 ( .Q(n709), .DIN1(n478), .DIN2(n479) );
    nor2s1 U249 ( .Q(n710), .DIN1(n482), .DIN2(n484) );
    nnd2s1 U250 ( .Q(n390), .DIN1(n710), .DIN2(n709) );
    nnd2s1 U251 ( .Q(n279), .DIN1(n711), .DIN2(N11) );
    nnd2s1 U252 ( .Q(n280), .DIN1(n712), .DIN2(n713) );
    nnd2s1 U253 ( .Q(n439), .DIN1(N237), .DIN2(N1726) );
    hi1s1 U254 ( .Q(n714), .DIN(N256) );
    hi1s1 U255 ( .Q(n715), .DIN(N259) );
    hi1s1 U256 ( .Q(n716), .DIN(N346) );
    hi1s1 U257 ( .Q(n717), .DIN(N349) );
    nor2s1 U258 ( .Q(n718), .DIN1(N349), .DIN2(n716) );
    nor2s1 U259 ( .Q(n719), .DIN1(N346), .DIN2(n717) );
    nor2s1 U260 ( .Q(n720), .DIN1(n718), .DIN2(n719) );
    nor2s1 U261 ( .Q(n721), .DIN1(N259), .DIN2(n714) );
    nor2s1 U262 ( .Q(n722), .DIN1(N256), .DIN2(n715) );
    nor2s1 U263 ( .Q(n723), .DIN1(n721), .DIN2(n722) );
    nnd2s1 U264 ( .Q(n724), .DIN1(n725), .DIN2(n726) );
    hi1s1 U265 ( .Q(n727), .DIN(n301) );
    hi1s1 U266 ( .Q(n728), .DIN(N1817) );
    hi1s1 U267 ( .Q(n729), .DIN(n320) );
    hi1s1 U268 ( .Q(n730), .DIN(N1818) );
    nor2s1 U269 ( .Q(n731), .DIN1(n552), .DIN2(n549) );
    nnd2s1 U270 ( .Q(n732), .DIN1(n549), .DIN2(n552) );
    nnd2s1 U271 ( .Q(n733), .DIN1(n734), .DIN2(n732) );
    nor2s1 U272 ( .Q(n735), .DIN1(N2018), .DIN2(N1819) );
    nor2s1 U273 ( .Q(n736), .DIN1(N2016), .DIN2(n283) );
    nor2s1 U274 ( .Q(n737), .DIN1(n735), .DIN2(n736) );
    nor2s1 U275 ( .Q(n738), .DIN1(N2022), .DIN2(n282) );
    nor2s1 U276 ( .Q(n739), .DIN1(N2020), .DIN2(n281) );
    nor2s1 U277 ( .Q(n740), .DIN1(n738), .DIN2(n739) );
    nnd2s1 U278 ( .Q(n741), .DIN1(n742), .DIN2(n743) );
    hi1s1 U279 ( .Q(n744), .DIN(N313) );
    hi1s1 U280 ( .Q(n291), .DIN(N316) );
    hi1s1 U281 ( .Q(n745), .DIN(N272) );
    hi1s1 U282 ( .Q(n746), .DIN(N269) );
    nor2s1 U283 ( .Q(n747), .DIN1(N281), .DIN2(n427) );
    nor2s1 U284 ( .Q(n748), .DIN1(N278), .DIN2(n428) );
    nor2s1 U285 ( .Q(n749), .DIN1(n747), .DIN2(n748) );
    nor2s1 U286 ( .Q(n750), .DIN1(N287), .DIN2(n425) );
    nor2s1 U287 ( .Q(n751), .DIN1(N284), .DIN2(n426) );
    nor2s1 U288 ( .Q(n752), .DIN1(n750), .DIN2(n751) );
    nnd2s1 U289 ( .Q(n753), .DIN1(n754), .DIN2(n755) );
    nor2s1 U290 ( .Q(n756), .DIN1(n662), .DIN2(n757) );
    nor2s1 U291 ( .Q(n758), .DIN1(n756), .DIN2(n745) );
    nor2s1 U292 ( .Q(n759), .DIN1(n402), .DIN2(n434) );
    nor2s1 U293 ( .Q(n435), .DIN1(n758), .DIN2(n759) );
    nor2s1 U294 ( .Q(n760), .DIN1(n756), .DIN2(n714) );
    nor2s1 U295 ( .Q(n761), .DIN1(n426), .DIN2(n434) );
    nor2s1 U296 ( .Q(n437), .DIN1(n760), .DIN2(n761) );
    nor2s1 U297 ( .Q(n762), .DIN1(n756), .DIN2(n715) );
    nor2s1 U298 ( .Q(n763), .DIN1(n422), .DIN2(n434) );
    nor2s1 U299 ( .Q(n764), .DIN1(n762), .DIN2(n763) );
    nor2s1 U300 ( .Q(n765), .DIN1(N297), .DIN2(n434) );
    nor2s1 U301 ( .Q(n766), .DIN1(n756), .DIN2(N263) );
    nor2s1 U302 ( .Q(n767), .DIN1(n765), .DIN2(n766) );
    hi1s1 U303 ( .Q(n768), .DIN(N246) );
    nnd2s1 U304 ( .Q(n769), .DIN1(n770), .DIN2(n441) );
    nor2s1 U305 ( .Q(n771), .DIN1(n772), .DIN2(n420) );
    nor2s1 U306 ( .Q(n773), .DIN1(n329), .DIN2(n769) );
    nor2s1 U307 ( .Q(N3546), .DIN1(n771), .DIN2(n773) );
    hi1s1 U308 ( .Q(n774), .DIN(N29) );
    nor2s1 U309 ( .Q(n775), .DIN1(N32), .DIN2(n426) );
    nor2s1 U310 ( .Q(n776), .DIN1(N287), .DIN2(n777) );
    nor2s1 U311 ( .Q(n678), .DIN1(n775), .DIN2(n776) );
    nor2s1 U312 ( .Q(n778), .DIN1(N26), .DIN2(n422) );
    nor2s1 U313 ( .Q(n779), .DIN1(N294), .DIN2(n780) );
    nor2s1 U314 ( .Q(n679), .DIN1(n778), .DIN2(n779) );
    nor2s1 U315 ( .Q(n781), .DIN1(N33), .DIN2(n401) );
    nor2s1 U316 ( .Q(n782), .DIN1(N297), .DIN2(n783) );
    nor2s1 U317 ( .Q(n681), .DIN1(n781), .DIN2(n782) );
    nor2s1 U318 ( .Q(n784), .DIN1(N35), .DIN2(n402) );
    nor2s1 U319 ( .Q(n785), .DIN1(N309), .DIN2(n786) );
    nor2s1 U320 ( .Q(n682), .DIN1(n784), .DIN2(n785) );
    nor2s1 U321 ( .Q(n787), .DIN1(N27), .DIN2(n400) );
    nor2s1 U322 ( .Q(n788), .DIN1(N301), .DIN2(n789) );
    nor2s1 U323 ( .Q(n684), .DIN1(n787), .DIN2(n788) );
    nor2s1 U324 ( .Q(n790), .DIN1(N34), .DIN2(n403) );
    nor2s1 U325 ( .Q(n791), .DIN1(N305), .DIN2(n792) );
    nor2s1 U326 ( .Q(n685), .DIN1(n790), .DIN2(n791) );
    nor2s1 U327 ( .Q(n793), .DIN1(N1817), .DIN2(n402) );
    nor2s1 U328 ( .Q(n794), .DIN1(N309), .DIN2(n728) );
    nor2s1 U329 ( .Q(n689), .DIN1(n793), .DIN2(n794) );
    nor2s1 U330 ( .Q(n795), .DIN1(n382), .DIN2(n774) );
    nor2s1 U331 ( .Q(n796), .DIN1(N29), .DIN2(n385) );
    nor2s1 U332 ( .Q(n713), .DIN1(n795), .DIN2(n796) );
    nor2s1 U333 ( .Q(n797), .DIN1(N4), .DIN2(n715) );
    nor2s1 U334 ( .Q(n798), .DIN1(N259), .DIN2(n799) );
    nor2s1 U335 ( .Q(n694), .DIN1(n797), .DIN2(n798) );
    nor2s1 U336 ( .Q(n800), .DIN1(N5), .DIN2(n424) );
    nor2s1 U337 ( .Q(n801), .DIN1(N266), .DIN2(n802) );
    nor2s1 U338 ( .Q(n696), .DIN1(n800), .DIN2(n801) );
    nor2s1 U339 ( .Q(n803), .DIN1(N21), .DIN2(n746) );
    nor2s1 U340 ( .Q(n804), .DIN1(N269), .DIN2(n805) );
    nor2s1 U341 ( .Q(n697), .DIN1(n803), .DIN2(n804) );
    nor2s1 U342 ( .Q(n806), .DIN1(N22), .DIN2(n745) );
    nor2s1 U343 ( .Q(n807), .DIN1(N272), .DIN2(n808) );
    nor2s1 U344 ( .Q(n699), .DIN1(n806), .DIN2(n807) );
    nor2s1 U345 ( .Q(n809), .DIN1(N23), .DIN2(n423) );
    nor2s1 U346 ( .Q(n810), .DIN1(N275), .DIN2(n811) );
    nor2s1 U347 ( .Q(n700), .DIN1(n809), .DIN2(n810) );
    nor2s1 U348 ( .Q(n812), .DIN1(N6), .DIN2(n427) );
    nor2s1 U349 ( .Q(n813), .DIN1(N278), .DIN2(n814) );
    nor2s1 U350 ( .Q(n702), .DIN1(n812), .DIN2(n813) );
    nor2s1 U351 ( .Q(n815), .DIN1(N24), .DIN2(n428) );
    nor2s1 U352 ( .Q(n816), .DIN1(N281), .DIN2(n817) );
    nor2s1 U353 ( .Q(n703), .DIN1(n815), .DIN2(n816) );
    nor2s1 U354 ( .Q(n818), .DIN1(n284), .DIN2(n429) );
    nor2s1 U355 ( .Q(n819), .DIN1(N2010), .DIN2(N263) );
    nor2s1 U356 ( .Q(n706), .DIN1(n818), .DIN2(n819) );
    nor2s1 U357 ( .Q(n820), .DIN1(n336), .DIN2(n715) );
    nor2s1 U358 ( .Q(n821), .DIN1(N259), .DIN2(n399) );
    nor2s1 U359 ( .Q(n705), .DIN1(n820), .DIN2(n821) );
    hi1s1 U360 ( .Q(n822), .DIN(N16) );
    nor2s1 U361 ( .Q(n823), .DIN1(n388), .DIN2(n822) );
    nor2s1 U362 ( .Q(n824), .DIN1(N16), .DIN2(n391) );
    nor2s1 U363 ( .Q(n712), .DIN1(n823), .DIN2(n824) );
    nor2s1 U364 ( .Q(n825), .DIN1(n301), .DIN2(n744) );
    nor2s1 U365 ( .Q(n826), .DIN1(N313), .DIN2(n727) );
    nor2s1 U366 ( .Q(n290), .DIN1(n825), .DIN2(n826) );
    hi1s1 U367 ( .Q(N3882), .DIN(N3881) );
    hi1s1 U368 ( .Q(n434), .DIN(n756) );
    nnd2s1 U369 ( .Q(n827), .DIN1(N219), .DIN2(N94) );
    hi1s1 U370 ( .Q(N1026), .DIN(n827) );
    hi1s1 U371 ( .Q(n572), .DIN(n419) );
    nnd2s1 U372 ( .Q(n514), .DIN1(N135), .DIN2(n404) );
    nnd2s1 U373 ( .Q(n513), .DIN1(N99), .DIN2(n406) );
    nnd2s1 U374 ( .Q(n516), .DIN1(N123), .DIN2(n407) );
    nnd2s1 U375 ( .Q(n515), .DIN1(N111), .DIN2(n409) );
    nnd2s1 U376 ( .Q(n518), .DIN1(N137), .DIN2(n404) );
    nnd2s1 U377 ( .Q(n517), .DIN1(N101), .DIN2(n406) );
    nnd2s1 U378 ( .Q(n520), .DIN1(N125), .DIN2(n407) );
    nnd2s1 U379 ( .Q(n519), .DIN1(N113), .DIN2(n409) );
    nnd2s1 U380 ( .Q(n522), .DIN1(N136), .DIN2(n404) );
    nnd2s1 U381 ( .Q(n521), .DIN1(N100), .DIN2(n406) );
    nnd2s1 U382 ( .Q(n524), .DIN1(N124), .DIN2(n407) );
    nnd2s1 U383 ( .Q(n523), .DIN1(N112), .DIN2(n409) );
    nnd2s1 U384 ( .Q(n526), .DIN1(N131), .DIN2(n404) );
    nnd2s1 U385 ( .Q(n525), .DIN1(N95), .DIN2(n406) );
    nnd2s1 U386 ( .Q(n528), .DIN1(N119), .DIN2(n407) );
    nnd2s1 U387 ( .Q(n527), .DIN1(N107), .DIN2(n409) );
    nnd2s1 U388 ( .Q(n502), .DIN1(N142), .DIN2(n404) );
    nnd2s1 U389 ( .Q(n501), .DIN1(N106), .DIN2(n406) );
    nnd2s1 U390 ( .Q(n504), .DIN1(N130), .DIN2(n407) );
    nnd2s1 U391 ( .Q(n503), .DIN1(N118), .DIN2(n409) );
    nnd2s1 U392 ( .Q(n506), .DIN1(N141), .DIN2(n404) );
    nnd2s1 U393 ( .Q(n505), .DIN1(N105), .DIN2(n406) );
    nnd2s1 U394 ( .Q(n508), .DIN1(N129), .DIN2(n407) );
    nnd2s1 U395 ( .Q(n507), .DIN1(N117), .DIN2(n409) );
    nnd2s1 U396 ( .Q(n510), .DIN1(N140), .DIN2(n404) );
    nnd2s1 U397 ( .Q(n509), .DIN1(N104), .DIN2(n406) );
    nnd2s1 U398 ( .Q(n512), .DIN1(N128), .DIN2(n407) );
    nnd2s1 U399 ( .Q(n511), .DIN1(N116), .DIN2(n409) );
    nnd2s1 U400 ( .Q(n530), .DIN1(N139), .DIN2(n404) );
    nnd2s1 U401 ( .Q(n529), .DIN1(N103), .DIN2(n406) );
    nnd2s1 U402 ( .Q(n532), .DIN1(N127), .DIN2(n407) );
    nnd2s1 U403 ( .Q(n531), .DIN1(N115), .DIN2(n409) );
    nnd2s1 U404 ( .Q(n534), .DIN1(N138), .DIN2(n404) );
    nnd2s1 U405 ( .Q(n533), .DIN1(N102), .DIN2(n406) );
    nnd2s1 U406 ( .Q(n536), .DIN1(N126), .DIN2(n407) );
    nnd2s1 U407 ( .Q(n535), .DIN1(N114), .DIN2(n409) );
    nor2s1 U408 ( .Q(N3671), .DIN1(n733), .DIN2(N37) );
    nnd2s1 U409 ( .Q(n556), .DIN1(N89), .DIN2(n414) );
    nnd2s1 U410 ( .Q(n555), .DIN1(N76), .DIN2(n416) );
    nnd2s1 U411 ( .Q(n558), .DIN1(N51), .DIN2(n418) );
    nnd2s1 U412 ( .Q(n557), .DIN1(N63), .DIN2(n419) );
    nnd2s1 U413 ( .Q(n560), .DIN1(N90), .DIN2(n414) );
    nnd2s1 U414 ( .Q(n559), .DIN1(N77), .DIN2(n416) );
    nnd2s1 U415 ( .Q(n562), .DIN1(N52), .DIN2(n418) );
    nnd2s1 U416 ( .Q(n561), .DIN1(N64), .DIN2(n419) );
    nnd2s1 U417 ( .Q(n580), .DIN1(N93), .DIN2(n414) );
    nnd2s1 U418 ( .Q(n579), .DIN1(N80), .DIN2(n416) );
    nnd2s1 U419 ( .Q(n582), .DIN1(N55), .DIN2(n418) );
    nnd2s1 U420 ( .Q(n581), .DIN1(N67), .DIN2(n419) );
    nnd2s1 U421 ( .Q(n584), .DIN1(N81), .DIN2(n414) );
    nnd2s1 U422 ( .Q(n583), .DIN1(N68), .DIN2(n416) );
    nnd2s1 U423 ( .Q(n586), .DIN1(N43), .DIN2(n418) );
    nnd2s1 U424 ( .Q(n585), .DIN1(N56), .DIN2(n419) );
    nnd2s1 U425 ( .Q(n588), .DIN1(N91), .DIN2(n414) );
    nnd2s1 U426 ( .Q(n587), .DIN1(N78), .DIN2(n416) );
    nnd2s1 U427 ( .Q(n590), .DIN1(N53), .DIN2(n418) );
    nnd2s1 U428 ( .Q(n589), .DIN1(N65), .DIN2(n419) );
    nnd2s1 U429 ( .Q(n592), .DIN1(N92), .DIN2(n414) );
    nnd2s1 U430 ( .Q(n591), .DIN1(N79), .DIN2(n416) );
    nnd2s1 U431 ( .Q(n594), .DIN1(N54), .DIN2(n418) );
    nnd2s1 U432 ( .Q(n593), .DIN1(N66), .DIN2(n419) );
    nnd2s1 U433 ( .Q(n564), .DIN1(N85), .DIN2(n414) );
    nnd2s1 U434 ( .Q(n563), .DIN1(N72), .DIN2(n416) );
    nnd2s1 U435 ( .Q(n566), .DIN1(N47), .DIN2(n418) );
    nnd2s1 U436 ( .Q(n565), .DIN1(N60), .DIN2(n419) );
    nnd2s1 U437 ( .Q(n568), .DIN1(N86), .DIN2(n414) );
    nnd2s1 U438 ( .Q(n567), .DIN1(N73), .DIN2(n416) );
    nnd2s1 U439 ( .Q(n570), .DIN1(N48), .DIN2(n418) );
    nnd2s1 U440 ( .Q(n569), .DIN1(N61), .DIN2(n419) );
    nnd2s1 U441 ( .Q(n571), .DIN1(N49), .DIN2(n418) );
    nnd2s1 U442 ( .Q(n574), .DIN1(N87), .DIN2(n415) );
    nnd2s1 U443 ( .Q(n573), .DIN1(N74), .DIN2(N234) );
    nnd2s1 U444 ( .Q(n576), .DIN1(N88), .DIN2(n414) );
    nnd2s1 U445 ( .Q(n575), .DIN1(N75), .DIN2(n416) );
    nnd2s1 U446 ( .Q(n578), .DIN1(N50), .DIN2(n418) );
    nnd2s1 U447 ( .Q(n577), .DIN1(N62), .DIN2(n419) );
    nnd2s1 U448 ( .Q(n742), .DIN1(n740), .DIN2(n828) );
    nnd2s1 U449 ( .Q(n743), .DIN1(n737), .DIN2(n829) );
    hi1s1 U450 ( .Q(n830), .DIN(n741) );
    nor2s1 U451 ( .Q(N3809), .DIN1(n831), .DIN2(N37) );
    nnd2s1 U452 ( .Q(n754), .DIN1(n752), .DIN2(n832) );
    nnd2s1 U453 ( .Q(n755), .DIN1(n749), .DIN2(n833) );
    nnd2s1 U454 ( .Q(n725), .DIN1(n723), .DIN2(n834) );
    nnd2s1 U455 ( .Q(n726), .DIN1(n720), .DIN2(n835) );
    nnd2s1 U456 ( .Q(n656), .DIN1(N14), .DIN2(n836) );
    hi1s1 U457 ( .Q(N2925), .DIN(n656) );
    nnd2s1 U458 ( .Q(n432), .DIN1(N325), .DIN2(n296) );
    nnd2s1 U459 ( .Q(n431), .DIN1(N231), .DIN2(n295) );
    hi1s1 U460 ( .Q(N1726), .DIN(n430) );
    hi1s1 U461 ( .Q(n837), .DIN(n349) );
    nnd2s1 U462 ( .Q(n838), .DIN1(n659), .DIN2(n837) );
    nnd2s1 U463 ( .Q(n667), .DIN1(n660), .DIN2(n837) );
    nnd2s1 U464 ( .Q(n668), .DIN1(n661), .DIN2(n837) );
    nnd2s1 U465 ( .Q(n839), .DIN1(n399), .DIN2(n436) );
    nnd2s1 U466 ( .Q(n361), .DIN1(n764), .DIN2(n839) );
    nnd2s1 U467 ( .Q(n360), .DIN1(n840), .DIN2(n336) );
    nnd2s1 U468 ( .Q(n366), .DIN1(n663), .DIN2(n841) );
    nnd2s1 U469 ( .Q(n365), .DIN1(n363), .DIN2(N1821) );
    hi1s1 U470 ( .Q(n396), .DIN(n364) );
    nnd2s1 U471 ( .Q(n842), .DIN1(n670), .DIN2(n668) );
    nnd2s1 U472 ( .Q(n843), .DIN1(n308), .DIN2(n425) );
    nnd2s1 U473 ( .Q(n844), .DIN1(n843), .DIN2(n842) );
    nnd2s1 U474 ( .Q(n845), .DIN1(n844), .DIN2(n667) );
    nnd2s1 U475 ( .Q(n846), .DIN1(n455), .DIN2(n845) );
    nnd2s1 U476 ( .Q(n847), .DIN1(n669), .DIN2(n848) );
    nnd2s1 U477 ( .Q(n849), .DIN1(n837), .DIN2(n846) );
    nnd2s1 U478 ( .Q(n850), .DIN1(n849), .DIN2(n847) );
    nnd2s1 U479 ( .Q(n289), .DIN1(n658), .DIN2(n837) );
    nnd2s1 U480 ( .Q(n288), .DIN1(n850), .DIN2(n838) );
    hi1s1 U481 ( .Q(n851), .DIN(n438) );
    nnd2s1 U482 ( .Q(n293), .DIN1(N1), .DIN2(N3) );
    hi1s1 U483 ( .Q(N1448), .DIN(N1277) );
    hi1s1 U484 ( .Q(n297), .DIN(N1028) );
    nnd2s1 U485 ( .Q(n852), .DIN1(n359), .DIN2(n284) );
    nnd2s1 U486 ( .Q(n665), .DIN1(n368), .DIN2(n369) );
    nnd2s1 U487 ( .Q(n841), .DIN1(n767), .DIN2(n852) );
    nnd2s1 U488 ( .Q(n664), .DIN1(n395), .DIN2(n396) );
    nnd2s1 U489 ( .Q(n397), .DIN1(n851), .DIN2(n441) );
    nnd2s1 U490 ( .Q(n609), .DIN1(N340), .DIN2(n853) );
    nnd2s1 U491 ( .Q(n608), .DIN1(N343), .DIN2(n854) );
    nor2s1 U492 ( .Q(n612), .DIN1(n855), .DIN2(N337) );
    nnd2s1 U493 ( .Q(n856), .DIN1(N337), .DIN2(n855) );
    nnd2s1 U494 ( .Q(n857), .DIN1(n607), .DIN2(n610) );
    nor2s1 U495 ( .Q(n614), .DIN1(n610), .DIN2(n607) );
    nnd2s1 U496 ( .Q(n858), .DIN1(N256), .DIN2(n715) );
    nnd2s1 U497 ( .Q(n859), .DIN1(N259), .DIN2(n714) );
    nnd2s1 U498 ( .Q(n835), .DIN1(n859), .DIN2(n858) );
    nnd2s1 U499 ( .Q(n860), .DIN1(N346), .DIN2(n717) );
    nnd2s1 U500 ( .Q(n861), .DIN1(N349), .DIN2(n716) );
    nnd2s1 U501 ( .Q(n834), .DIN1(n861), .DIN2(n860) );
    nnd2s1 U502 ( .Q(n618), .DIN1(N328), .DIN2(n862) );
    nnd2s1 U503 ( .Q(n617), .DIN1(N331), .DIN2(n863) );
    nor2s1 U504 ( .Q(n864), .DIN1(n724), .DIN2(n616) );
    nnd2s1 U505 ( .Q(n620), .DIN1(n616), .DIN2(n724) );
    nor2s1 U506 ( .Q(n865), .DIN1(n613), .DIN2(n619) );
    nnd2s1 U507 ( .Q(n866), .DIN1(n619), .DIN2(n613) );
    nnd2s1 U508 ( .Q(n836), .DIN1(n866), .DIN2(n867) );
    nor2s1 U509 ( .Q(n551), .DIN1(n868), .DIN2(n314) );
    nor2s1 U510 ( .Q(n550), .DIN1(n410), .DIN2(n311) );
    nnd2s1 U511 ( .Q(n539), .DIN1(n301), .DIN2(n412) );
    nnd2s1 U512 ( .Q(n538), .DIN1(N1816), .DIN2(n727) );
    nor2s1 U513 ( .Q(n542), .DIN1(n728), .DIN2(n537) );
    nor2s1 U514 ( .Q(n541), .DIN1(n869), .DIN2(N1817) );
    hi1s1 U515 ( .Q(n870), .DIN(n540) );
    nnd2s1 U516 ( .Q(n545), .DIN1(n308), .DIN2(n729) );
    nnd2s1 U517 ( .Q(n544), .DIN1(n320), .DIN2(n413) );
    nor2s1 U518 ( .Q(n548), .DIN1(n730), .DIN2(n543) );
    nor2s1 U519 ( .Q(n547), .DIN1(n871), .DIN2(N1818) );
    nor2s1 U520 ( .Q(n448), .DIN1(n540), .DIN2(n872) );
    nor2s1 U521 ( .Q(n447), .DIN1(n546), .DIN2(n870) );
    nnd2s1 U522 ( .Q(n554), .DIN1(n446), .DIN2(n317) );
    nnd2s1 U523 ( .Q(n553), .DIN1(n873), .DIN2(n411) );
    nnd2s1 U524 ( .Q(n603), .DIN1(N2012), .DIN2(N1820) );
    nnd2s1 U525 ( .Q(n602), .DIN1(N2014), .DIN2(N1821) );
    nnd2s1 U526 ( .Q(n874), .DIN1(N2020), .DIN2(n281) );
    nnd2s1 U527 ( .Q(n875), .DIN1(N2022), .DIN2(n282) );
    nnd2s1 U528 ( .Q(n829), .DIN1(n875), .DIN2(n874) );
    nnd2s1 U529 ( .Q(n876), .DIN1(N2016), .DIN2(n283) );
    nnd2s1 U530 ( .Q(n877), .DIN1(N2018), .DIN2(N1819) );
    nnd2s1 U531 ( .Q(n828), .DIN1(n877), .DIN2(n876) );
    nnd2s1 U532 ( .Q(n597), .DIN1(n329), .DIN2(n421) );
    nnd2s1 U533 ( .Q(n596), .DIN1(n294), .DIN2(n420) );
    nnd2s1 U534 ( .Q(n600), .DIN1(n399), .DIN2(n284) );
    nnd2s1 U535 ( .Q(n599), .DIN1(n336), .DIN2(N2010) );
    nnd2s1 U536 ( .Q(n878), .DIN1(n595), .DIN2(n879) );
    nor2s1 U537 ( .Q(n450), .DIN1(n879), .DIN2(n595) );
    nnd2s1 U538 ( .Q(n880), .DIN1(n830), .DIN2(n449) );
    nor2s1 U539 ( .Q(n605), .DIN1(n449), .DIN2(n830) );
    nnd2s1 U540 ( .Q(n881), .DIN1(n601), .DIN2(n604) );
    nor2s1 U541 ( .Q(n882), .DIN1(n604), .DIN2(n601) );
    nor2s1 U542 ( .Q(n831), .DIN1(n882), .DIN2(n883) );
    nnd2s1 U543 ( .Q(n639), .DIN1(N313), .DIN2(n291) );
    nnd2s1 U544 ( .Q(n638), .DIN1(N316), .DIN2(n744) );
    nnd2s1 U545 ( .Q(n642), .DIN1(N305), .DIN2(n402) );
    nnd2s1 U546 ( .Q(n641), .DIN1(N309), .DIN2(n403) );
    nnd2s1 U547 ( .Q(n645), .DIN1(n637), .DIN2(n884) );
    nnd2s1 U548 ( .Q(n644), .DIN1(n640), .DIN2(n885) );
    nnd2s1 U549 ( .Q(n648), .DIN1(N297), .DIN2(n400) );
    nnd2s1 U550 ( .Q(n647), .DIN1(N301), .DIN2(n401) );
    nor2s1 U551 ( .Q(n651), .DIN1(n422), .DIN2(N355) );
    nor2s1 U552 ( .Q(n650), .DIN1(n886), .DIN2(N294) );
    nnd2s1 U553 ( .Q(n887), .DIN1(n646), .DIN2(n649) );
    nor2s1 U554 ( .Q(n653), .DIN1(n649), .DIN2(n646) );
    nnd2s1 U555 ( .Q(n888), .DIN1(n643), .DIN2(n652) );
    nor2s1 U556 ( .Q(n889), .DIN1(n652), .DIN2(n643) );
    nor2s1 U557 ( .Q(N2970), .DIN1(n889), .DIN2(n890) );
    nnd2s1 U558 ( .Q(n624), .DIN1(N272), .DIN2(n423) );
    nnd2s1 U559 ( .Q(n623), .DIN1(N275), .DIN2(n745) );
    nnd2s1 U560 ( .Q(n627), .DIN1(N266), .DIN2(n746) );
    nnd2s1 U561 ( .Q(n626), .DIN1(N269), .DIN2(n424) );
    nor2s1 U562 ( .Q(n630), .DIN1(n891), .DIN2(n625) );
    nnd2s1 U563 ( .Q(n892), .DIN1(n625), .DIN2(n891) );
    nnd2s1 U564 ( .Q(n893), .DIN1(N284), .DIN2(n426) );
    nnd2s1 U565 ( .Q(n894), .DIN1(N287), .DIN2(n425) );
    nnd2s1 U566 ( .Q(n833), .DIN1(n894), .DIN2(n893) );
    nnd2s1 U567 ( .Q(n895), .DIN1(N278), .DIN2(n428) );
    nnd2s1 U568 ( .Q(n896), .DIN1(N281), .DIN2(n427) );
    nnd2s1 U569 ( .Q(n832), .DIN1(n896), .DIN2(n895) );
    nnd2s1 U570 ( .Q(n633), .DIN1(N263), .DIN2(n897) );
    nnd2s1 U571 ( .Q(n632), .DIN1(N352), .DIN2(n429) );
    nor2s1 U572 ( .Q(n898), .DIN1(n753), .DIN2(n631) );
    nnd2s1 U573 ( .Q(n635), .DIN1(n631), .DIN2(n753) );
    nor2s1 U574 ( .Q(n899), .DIN1(n628), .DIN2(n634) );
    nnd2s1 U575 ( .Q(n452), .DIN1(n634), .DIN2(n628) );
    nnd2s1 U576 ( .Q(n488), .DIN1(N269), .DIN2(n434) );
    nnd2s1 U577 ( .Q(n487), .DIN1(n756), .DIN2(N305) );
    nnd2s1 U578 ( .Q(n486), .DIN1(n756), .DIN2(n400) );
    nnd2s1 U579 ( .Q(n485), .DIN1(n424), .DIN2(n434) );
    nnd2s1 U580 ( .Q(n673), .DIN1(n830), .DIN2(n851) );
    nnd2s1 U581 ( .Q(n672), .DIN1(n438), .DIN2(n741) );
    nor2s1 U582 ( .Q(n900), .DIN1(n449), .DIN2(n671) );
    nnd2s1 U583 ( .Q(n901), .DIN1(n671), .DIN2(n449) );
    nnd2s1 U584 ( .Q(n902), .DIN1(n901), .DIN2(n903) );
    nnd2s1 U585 ( .Q(n490), .DIN1(n420), .DIN2(n768) );
    nnd2s1 U586 ( .Q(n489), .DIN1(N246), .DIN2(n902) );
    nnd2s1 U587 ( .Q(n676), .DIN1(n294), .DIN2(n399) );
    nnd2s1 U588 ( .Q(n675), .DIN1(n336), .DIN2(n421) );
    nnd2s1 U589 ( .Q(n904), .DIN1(n905), .DIN2(n438) );
    nnd2s1 U590 ( .Q(n906), .DIN1(n674), .DIN2(n851) );
    nnd2s1 U591 ( .Q(n770), .DIN1(n906), .DIN2(n904) );
    nnd2s1 U592 ( .Q(n493), .DIN1(N25), .DIN2(n774) );
    nnd2s1 U593 ( .Q(n492), .DIN1(N29), .DIN2(n413) );
    nnd2s1 U594 ( .Q(n907), .DIN1(n908), .DIN2(N284) );
    nnd2s1 U595 ( .Q(n909), .DIN1(n491), .DIN2(n425) );
    nnd2s1 U596 ( .Q(n711), .DIN1(n909), .DIN2(n907) );
    nnd2s1 U597 ( .Q(n456), .DIN1(N287), .DIN2(n410) );
    nnd2s1 U598 ( .Q(n455), .DIN1(n314), .DIN2(n426) );
    nnd2s1 U599 ( .Q(n459), .DIN1(N294), .DIN2(n411) );
    nnd2s1 U600 ( .Q(n458), .DIN1(n317), .DIN2(n422) );
    nnd2s1 U601 ( .Q(n462), .DIN1(N301), .DIN2(n730) );
    nnd2s1 U602 ( .Q(n461), .DIN1(N1818), .DIN2(n400) );
    nnd2s1 U603 ( .Q(n465), .DIN1(N305), .DIN2(n412) );
    nnd2s1 U604 ( .Q(n464), .DIN1(N1816), .DIN2(n403) );
    nnd2s1 U605 ( .Q(n468), .DIN1(N297), .DIN2(n729) );
    nnd2s1 U606 ( .Q(n467), .DIN1(n320), .DIN2(n401) );
    nnd2s1 U607 ( .Q(n910), .DIN1(N263), .DIN2(n911) );
    nnd2s1 U608 ( .Q(n912), .DIN1(N20), .DIN2(n429) );
    nnd2s1 U609 ( .Q(n692), .DIN1(n912), .DIN2(n910) );
    nnd2s1 U610 ( .Q(n913), .DIN1(N256), .DIN2(n914) );
    nnd2s1 U611 ( .Q(n915), .DIN1(N19), .DIN2(n714) );
    nnd2s1 U612 ( .Q(n691), .DIN1(n915), .DIN2(n913) );
    nnd2s1 U613 ( .Q(n471), .DIN1(N256), .DIN2(n421) );
    nnd2s1 U614 ( .Q(n470), .DIN1(n294), .DIN2(n714) );
    nnd2s1 U615 ( .Q(n474), .DIN1(N269), .DIN2(N2014) );
    nnd2s1 U616 ( .Q(n473), .DIN1(n746), .DIN2(N1820) );
    nnd2s1 U617 ( .Q(n477), .DIN1(N266), .DIN2(N2012) );
    nnd2s1 U618 ( .Q(n476), .DIN1(n424), .DIN2(N1821) );
    nnd2s1 U619 ( .Q(n355), .DIN1(N275), .DIN2(N2018) );
    nnd2s1 U620 ( .Q(n375), .DIN1(n423), .DIN2(n283) );
    nnd2s1 U621 ( .Q(n481), .DIN1(N272), .DIN2(N2016) );
    nnd2s1 U622 ( .Q(n480), .DIN1(n745), .DIN2(N1819) );
    nnd2s1 U623 ( .Q(n350), .DIN1(N281), .DIN2(N2022) );
    nnd2s1 U624 ( .Q(n483), .DIN1(n428), .DIN2(n281) );
    nnd2s1 U625 ( .Q(n353), .DIN1(N278), .DIN2(N2020) );
    nnd2s1 U626 ( .Q(n379), .DIN1(n427), .DIN2(n282) );
    nnd2s1 U627 ( .Q(n495), .DIN1(n421), .DIN2(n768) );
    nnd2s1 U628 ( .Q(n494), .DIN1(N246), .DIN2(n851) );
    nnd2s1 U629 ( .Q(n497), .DIN1(N246), .DIN2(N2014) );
    nnd2s1 U630 ( .Q(n496), .DIN1(N2010), .DIN2(n768) );
    nnd2s1 U631 ( .Q(n499), .DIN1(N246), .DIN2(N2012) );
    nnd2s1 U632 ( .Q(n498), .DIN1(n399), .DIN2(n768) );
    hi1s1 U633 ( .Q(n300), .DIN(n500) );
    hi1s1 U634 ( .Q(n408), .DIN(N322) );
    hi1s1 U635 ( .Q(n848), .DIN(n666) );
    hi1s1 U636 ( .Q(n440), .DIN(N224) );
    hi1s1 U637 ( .Q(n867), .DIN(n865) );
    hi1s1 U638 ( .Q(n621), .DIN(n864) );
    hi1s1 U639 ( .Q(n890), .DIN(n888) );
    hi1s1 U640 ( .Q(n615), .DIN(n857) );
    hi1s1 U641 ( .Q(n654), .DIN(n887) );
    hi1s1 U642 ( .Q(n883), .DIN(n881) );
    hi1s1 U643 ( .Q(n734), .DIN(n731) );
    hi1s1 U644 ( .Q(n453), .DIN(n899) );
    hi1s1 U645 ( .Q(n636), .DIN(n898) );
    hi1s1 U646 ( .Q(n891), .DIN(n622) );
    hi1s1 U647 ( .Q(n885), .DIN(n637) );
    hi1s1 U648 ( .Q(n863), .DIN(N328) );
    hi1s1 U649 ( .Q(n855), .DIN(N334) );
    hi1s1 U650 ( .Q(n854), .DIN(N340) );
    hi1s1 U651 ( .Q(n879), .DIN(n598) );
    hi1s1 U652 ( .Q(n903), .DIN(n900) );
    hi1s1 U653 ( .Q(n897), .DIN(N352) );
    hi1s1 U654 ( .Q(n629), .DIN(n892) );
    hi1s1 U655 ( .Q(n886), .DIN(N355) );
    hi1s1 U656 ( .Q(n884), .DIN(n640) );
    hi1s1 U657 ( .Q(n862), .DIN(N331) );
    hi1s1 U658 ( .Q(n611), .DIN(n856) );
    hi1s1 U659 ( .Q(n853), .DIN(N343) );
    hi1s1 U660 ( .Q(n417), .DIN(N234) );
    hi1s1 U661 ( .Q(n451), .DIN(n878) );
    hi1s1 U662 ( .Q(n606), .DIN(n880) );
    hi1s1 U663 ( .Q(n871), .DIN(n543) );
    hi1s1 U664 ( .Q(n869), .DIN(n537) );
    hi1s1 U665 ( .Q(n872), .DIN(n546) );
    hi1s1 U666 ( .Q(n873), .DIN(n446) );
    hi1s1 U667 ( .Q(n868), .DIN(n311) );
    hi1s1 U668 ( .Q(n757), .DIN(n347) );
    hi1s1 U669 ( .Q(n840), .DIN(n436) );
    hi1s1 U670 ( .Q(n905), .DIN(n674) );
    hi1s1 U671 ( .Q(n772), .DIN(n769) );
    hi1s1 U672 ( .Q(n908), .DIN(n491) );
    hi1s1 U673 ( .Q(n802), .DIN(N5) );
    hi1s1 U674 ( .Q(n805), .DIN(N21) );
    hi1s1 U675 ( .Q(n799), .DIN(N4) );
    hi1s1 U676 ( .Q(n914), .DIN(N19) );
    hi1s1 U677 ( .Q(n911), .DIN(N20) );
    hi1s1 U678 ( .Q(n814), .DIN(N6) );
    hi1s1 U679 ( .Q(n817), .DIN(N24) );
    hi1s1 U680 ( .Q(n808), .DIN(N22) );
    hi1s1 U681 ( .Q(n811), .DIN(N23) );
    hi1s1 U682 ( .Q(n783), .DIN(N33) );
    hi1s1 U683 ( .Q(n786), .DIN(N35) );
    hi1s1 U684 ( .Q(n777), .DIN(N32) );
    hi1s1 U685 ( .Q(n780), .DIN(N26) );
    hi1s1 U686 ( .Q(n789), .DIN(N27) );
    hi1s1 U687 ( .Q(n792), .DIN(N34) );
  nor4s1 troj59_0U1 ( .DIN1(troj59_0n1), .DIN2(troj59_0n2), .DIN3(troj59_0n3), .DIN4(troj59_0n4), .Q(Trigger_en59_0)         );
  nnd2s1 troj59_0U2 ( .DIN1(n671), .DIN2(n665), .Q(troj59_0n4) );
  i1s1 troj59_0U3 ( .DIN(n716), .Q(troj59_0n3) );
  nnd2s1 troj59_0U4 ( .DIN1(n818), .DIN2(n784), .Q(troj59_0n2) );
  or5s1 troj59_0U5 ( .DIN1(n849), .DIN2(n847), .DIN3(n522), .DIN4(troj59_0n5), .DIN5(troj59_0n6), .Q(troj59_0n1) );
  nnd2s1 troj59_0U6 ( .DIN1(n484), .DIN2(n309), .Q(troj59_0n6) );
  i1s1 troj59_0U7 ( .DIN(n546), .Q(troj59_0n5) );
    xor2s1 trojan59_0  (.DIN1(tempn391), .DIN2(Trigger_en59_0), .Q(n391) );

endmodule

