
module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si, test_so );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so;
  wire   CRC_OUT_1_31, WX9949, WX9947, WX9945, WX9943, WX9941, WX9939, WX9937,
         WX9935, WX9933, WX9931, WX9929, WX9927, WX9925, WX9923, WX9921,
         WX9919, WX9917, WX9915, WX9913, WX9911, WX9909, WX9907, WX9905,
         WX9903, WX9901, WX9899, WX9897, WX9895, WX9893, WX9891, WX9889,
         WX9887, WX9885, WX9883, WX9881, WX9879, WX9877, WX9875, WX9873,
         WX9871, WX9869, WX9867, WX9865, WX9863, WX9861, WX9859, WX9857,
         WX9855, WX9853, WX9851, WX9849, WX9847, WX9845, WX9843, WX9841,
         WX9839, WX9837, WX9835, WX9833, WX9831, WX9829, WX9827, WX9825,
         WX9823, WX9821, WX9819, WX9817, WX9815, WX9813, WX9811, WX9809,
         WX9807, WX9805, WX9803, WX9801, WX9799, WX9797, WX9795, WX9793,
         WX9791, WX9789, WX9787, WX9785, WX9783, WX9781, WX9779, WX9777,
         WX9775, WX9773, WX9771, WX9769, WX9767, WX9765, WX9763, WX9761,
         WX9759, WX9757, WX9755, WX9753, WX9751, WX9749, WX9747, WX9745,
         WX9743, WX9741, WX9739, WX9737, WX9735, WX9733, WX9731, WX9729,
         WX9727, WX9725, WX9723, WX9721, WX9719, WX9717, WX9715, WX9713,
         WX9711, WX9709, WX9707, WX9705, WX9703, WX9701, WX9699, WX9697,
         WX9695, WX9597, WX9595, WX9593, WX9591, WX9589, WX9587, WX9585,
         WX9583, WX9581, WX9579, WX9577, WX9575, WX9573, WX9571, WX9569,
         WX9567, WX9565, WX9563, WX9561, WX9559, WX9557, WX9555, WX9553,
         WX9551, WX9549, WX9547, WX9545, WX9543, WX9541, WX9539, WX9537,
         WX9535, WX9084, WX9082, WX9080, WX9078, WX9076, WX9074, WX9072,
         WX9070, WX9068, WX9066, WX9064, WX9062, WX9060, WX9058, WX9056,
         WX9054, WX9052, WX9050, WX9048, WX9046, WX9044, WX9042, WX9040,
         WX9038, WX9036, WX9034, WX9032, WX9030, WX9028, WX9026, WX9024,
         WX9022, WX898, WX896, WX894, WX892, WX890, WX888, WX886, WX884, WX882,
         WX880, WX878, WX876, WX874, WX872, WX870, WX868, WX866, WX8656,
         WX8654, WX8652, WX8650, WX8648, WX8646, WX8644, WX8642, WX8640, WX864,
         WX8638, WX8636, WX8634, WX8632, WX8630, WX8628, WX8626, WX8624,
         WX8622, WX8620, WX862, WX8618, WX8616, WX8614, WX8612, WX8610, WX8608,
         WX8606, WX8604, WX8602, WX8600, WX860, WX8598, WX8596, WX8594, WX8592,
         WX8590, WX8588, WX8586, WX8584, WX8582, WX8580, WX858, WX8578, WX8576,
         WX8574, WX8572, WX8570, WX8568, WX8566, WX8564, WX8562, WX8560, WX856,
         WX8558, WX8556, WX8554, WX8552, WX8550, WX8548, WX8546, WX8544,
         WX8542, WX8540, WX854, WX8538, WX8536, WX8534, WX8532, WX8530, WX8528,
         WX8526, WX8524, WX8522, WX8520, WX852, WX8518, WX8516, WX8514, WX8512,
         WX8510, WX8508, WX8506, WX8504, WX8502, WX8500, WX850, WX8498, WX8496,
         WX8494, WX8492, WX8490, WX8488, WX8486, WX8484, WX8482, WX8480, WX848,
         WX8478, WX8476, WX8474, WX8472, WX8470, WX8468, WX8466, WX8464, n3205,
         WX8462, n3206, WX8460, n3207, WX846, WX8458, n3208, WX8456, n3209,
         WX8454, n3210, WX8452, n3211, WX8450, n3212, WX8448, n3213, WX8446,
         n3214, WX8444, n3215, WX8442, n3216, WX8440, n3217, WX844, WX8438,
         n3218, WX8436, n3219, WX8434, n3220, WX8432, WX8430, WX8428, WX8426,
         WX8424, WX8422, WX8420, WX842, WX8418, WX8416, WX8414, WX8412, WX8410,
         WX8408, WX8406, WX8404, WX8402, WX840, WX838, WX836, WX834, WX832,
         WX8304, WX8302, WX8300, WX830, WX8298, WX8296, WX8294, WX8292, WX8290,
         WX8288, WX8286, WX8284, WX8282, WX8280, WX828, WX8278, WX8276, WX8274,
         WX8272, WX8270, WX8268, WX8266, WX8264, WX8262, WX8260, WX826, WX8258,
         WX8256, WX8254, WX8252, WX8250, WX8248, WX8246, WX8244, WX8242, WX824,
         WX822, WX820, WX818, WX816, WX814, WX812, WX810, WX808, WX806, WX804,
         WX802, WX800, WX798, WX796, WX794, WX792, WX790, WX788, WX786, WX784,
         WX782, WX780, WX7791, WX7789, WX7787, WX7785, WX7783, WX7781, WX778,
         WX7779, WX7777, WX7775, WX7773, WX7771, WX7769, WX7767, WX7765,
         WX7763, WX7761, WX776, WX7759, WX7757, WX7755, WX7753, WX7751, WX7749,
         WX7747, WX7745, WX7743, WX7741, WX774, WX7739, WX7737, WX7735, WX7733,
         WX7731, WX7729, WX772, WX770, WX768, WX766, WX764, WX762, WX760,
         WX758, WX756, WX754, WX752, WX750, WX748, WX746, WX744, WX742, WX740,
         WX738, WX7363, WX7361, WX736, WX7359, WX7357, WX7355, WX7353, WX7351,
         WX7349, WX7347, WX7345, WX7343, WX7341, WX734, WX7339, WX7337, WX7335,
         WX7333, WX7331, WX7329, WX7327, WX7325, WX7323, WX7321, WX732, WX7319,
         WX7317, WX7315, WX7313, WX7311, WX7309, WX7307, WX7305, WX7303,
         WX7301, WX730, WX7299, WX7297, WX7295, WX7293, WX7291, WX7289, WX7287,
         WX7285, WX7283, WX7281, WX728, WX7279, WX7277, WX7275, WX7273, WX7271,
         WX7269, WX7267, WX7265, WX7263, WX7261, WX726, WX7259, WX7257, WX7255,
         WX7253, WX7251, WX7249, WX7247, WX7245, WX7243, WX7241, WX724, WX7239,
         WX7237, WX7235, WX7233, WX7231, WX7229, WX7227, WX7225, WX7223,
         WX7221, WX722, WX7219, WX7217, WX7215, WX7213, WX7211, WX7209, WX7207,
         WX7205, WX7203, WX7201, WX720, WX7199, WX7197, WX7195, WX7193, WX7191,
         WX7189, WX7187, WX7185, WX7183, WX7181, WX718, WX7179, WX7177, WX7175,
         WX7173, WX7171, n3221, WX7169, n3222, WX7167, n3223, WX7165, n3224,
         WX7163, n3225, WX7161, n3226, WX716, WX7159, n3227, WX7157, n3228,
         WX7155, n3229, WX7153, n3230, WX7151, n3231, WX7149, n3232, WX7147,
         n3233, WX7145, n3234, WX7143, n3235, WX7141, n3236, WX714, WX7139,
         WX7137, WX7135, WX7133, WX7131, WX7129, WX7127, WX7125, WX7123,
         WX7121, WX712, WX7119, WX7117, WX7115, WX7113, WX7111, WX7109, WX710,
         WX708, WX706, WX704, WX702, WX7011, WX7009, WX7007, WX7005, WX7003,
         WX7001, WX700, WX6999, WX6997, WX6995, WX6993, WX6991, WX6989, WX6987,
         WX6985, WX6983, WX6981, WX698, WX6979, WX6977, WX6975, WX6973, WX6971,
         WX6969, WX6967, WX6965, WX6963, WX6961, WX696, WX6959, WX6957, WX6955,
         WX6953, WX6951, WX6949, WX694, WX692, WX690, WX688, WX686, WX684,
         WX682, WX680, WX678, WX676, WX674, WX672, WX670, WX668, WX666, WX664,
         WX662, WX660, WX658, WX656, WX654, WX652, WX650, WX6498, WX6496,
         WX6494, WX6492, WX6490, WX6488, WX6486, WX6484, WX6482, WX6480, WX648,
         WX6478, WX6476, WX6474, WX6472, WX6470, WX6468, WX6466, WX6464,
         WX6462, WX6460, WX646, WX6458, WX6456, WX6454, WX6452, WX6450, WX6448,
         WX6446, WX6444, WX6442, WX6440, WX644, WX6438, WX6436, WX6070, WX6068,
         WX6066, WX6064, WX6062, WX6060, WX6058, WX6056, WX6054, WX6052,
         WX6050, WX6048, WX6046, WX6044, WX6042, WX6040, WX6038, WX6036,
         WX6034, WX6032, WX6030, WX6028, WX6026, WX6024, WX6022, WX6020,
         WX6018, WX6016, WX6014, WX6012, WX6010, WX6008, WX6006, WX6004,
         WX6002, WX6000, WX5998, WX5996, WX5994, WX5992, WX5990, WX5988,
         WX5986, WX5984, WX5982, WX5980, WX5978, WX5976, WX5974, WX5972,
         WX5970, WX5968, WX5966, WX5964, WX5962, WX5960, WX5958, WX5956,
         WX5954, WX5952, WX5950, WX5948, WX5946, WX5944, WX5942, WX5940,
         WX5938, WX5936, WX5934, WX5932, WX5930, WX5928, WX5926, WX5924,
         WX5922, WX5920, WX5918, WX5916, WX5914, WX5912, WX5910, WX5908,
         WX5906, WX5904, WX5902, WX5900, WX5898, WX5896, WX5894, WX5892,
         WX5890, WX5888, WX5886, WX5884, WX5882, WX5880, WX5878, n3237, WX5876,
         n3238, WX5874, n3239, WX5872, n3240, WX5870, n3241, WX5868, n3242,
         WX5866, n3243, WX5864, n3244, WX5862, n3245, WX5860, n3246, WX5858,
         n3247, WX5856, n3248, WX5854, n3249, WX5852, n3250, WX5850, n3251,
         WX5848, n3252, WX5846, WX5844, WX5842, WX5840, WX5838, WX5836, WX5834,
         WX5832, WX5830, WX5828, WX5826, WX5824, WX5822, WX5820, WX5818,
         WX5816, WX5718, WX5716, WX5714, WX5712, WX5710, WX5708, WX5706,
         WX5704, WX5702, WX5700, WX5698, WX5696, WX5694, WX5692, WX5690,
         WX5688, WX5686, WX5684, WX5682, WX5680, WX5678, WX5676, WX5674,
         WX5672, WX5670, WX5668, WX5666, WX5664, WX5662, WX5660, WX5658,
         WX5656, WX546, WX544, WX542, WX540, WX538, WX536, WX534, WX532, WX530,
         WX528, WX526, WX524, WX522, WX5205, WX5203, WX5201, WX520, WX5199,
         WX5197, WX5195, WX5193, WX5191, WX5189, WX5187, WX5185, WX5183,
         WX5181, WX518, WX5179, WX5177, WX5175, WX5173, WX5171, WX5169, WX5167,
         WX5165, WX5163, WX5161, WX516, WX5159, WX5157, WX5155, WX5153, WX5151,
         WX5149, WX5147, WX5145, WX5143, WX514, WX512, WX510, WX508, WX506,
         WX504, WX502, WX500, WX498, WX496, WX494, WX492, WX490, WX488, WX486,
         WX484, WX4777, WX4775, WX4773, WX4771, WX4769, WX4767, WX4765, WX4763,
         WX4761, WX4759, WX4757, WX4755, WX4753, WX4751, WX4749, WX4747,
         WX4745, WX4743, WX4741, WX4739, WX4737, WX4735, WX4733, WX4731,
         WX4729, WX4727, WX4725, WX4723, WX4721, WX4719, WX4717, WX4715,
         WX4713, WX4711, WX4709, WX4707, WX4705, WX4703, WX4701, WX4699,
         WX4697, WX4695, WX4693, WX4691, WX4689, WX4687, WX4685, WX4683,
         WX4681, WX4679, WX4677, WX4675, WX4673, WX4671, WX4669, WX4667,
         WX4665, WX4663, WX4661, WX4659, WX4657, WX4655, WX4653, WX4651,
         WX4649, WX4647, WX4645, WX4643, WX4641, WX4639, WX4637, WX4635,
         WX4633, WX4631, WX4629, WX4627, WX4625, WX4623, WX4621, WX4619,
         WX4617, WX4615, WX4613, WX4611, WX4609, WX4607, WX4605, WX4603,
         WX4601, WX4599, WX4597, WX4595, WX4593, WX4591, WX4589, WX4587,
         WX4585, n3253, WX4583, n3254, WX4581, n3255, WX4579, n3256, WX4577,
         n3257, WX4575, n3258, WX4573, n3259, WX4571, n3260, WX4569, n3261,
         WX4567, n3262, WX4565, n3263, WX4563, n3264, WX4561, n3265, WX4559,
         n3266, WX4557, n3267, WX4555, n3268, WX4553, WX4551, WX4549, WX4547,
         WX4545, WX4543, WX4541, WX4539, WX4537, WX4535, WX4533, WX4531,
         WX4529, WX4527, WX4525, WX4523, WX4425, WX4423, WX4421, WX4419,
         WX4417, WX4415, WX4413, WX4411, WX4409, WX4407, WX4405, WX4403,
         WX4401, WX4399, WX4397, WX4395, WX4393, WX4391, WX4389, WX4387,
         WX4385, WX4383, WX4381, WX4379, WX4377, WX4375, WX4373, WX4371,
         WX4369, WX4367, WX4365, WX4363, WX3912, WX3910, WX3908, WX3906,
         WX3904, WX3902, WX3900, WX3898, WX3896, WX3894, WX3892, WX3890,
         WX3888, WX3886, WX3884, WX3882, WX3880, WX3878, WX3876, WX3874,
         WX3872, WX3870, WX3868, WX3866, WX3864, WX3862, WX3860, WX3858,
         WX3856, WX3854, WX3852, WX3850, WX3484, WX3482, WX3480, WX3478,
         WX3476, WX3474, WX3472, WX3470, WX3468, WX3466, WX3464, WX3462,
         WX3460, WX3458, WX3456, WX3454, WX3452, WX3450, WX3448, WX3446,
         WX3444, WX3442, WX3440, WX3438, WX3436, WX3434, WX3432, WX3430,
         WX3428, WX3426, WX3424, WX3422, WX3420, WX3418, WX3416, WX3414,
         WX3412, WX3410, WX3408, WX3406, WX3404, WX3402, WX3400, WX3398,
         WX3396, WX3394, WX3392, WX3390, WX3388, WX3386, WX3384, WX3382,
         WX3380, WX3378, WX3376, WX3374, WX3372, WX3370, WX3368, WX3366,
         WX3364, WX3362, WX3360, WX3358, WX3356, WX3354, WX3352, WX3350,
         WX3348, WX3346, WX3344, WX3342, WX3340, WX3338, WX3336, WX3334,
         WX3332, WX3330, WX3328, WX3326, WX3324, WX3322, WX3320, WX3318,
         WX3316, WX3314, WX3312, WX3310, WX3308, WX3306, WX3304, WX3302,
         WX3300, WX3298, WX3296, WX3294, WX3292, n3269, WX3290, n3270, WX3288,
         n3271, WX3286, n3272, WX3284, n3273, WX3282, n3274, WX3280, n3275,
         WX3278, n3276, WX3276, n3277, WX3274, n3278, WX3272, n3279, WX3270,
         n3280, WX3268, n3281, WX3266, n3282, WX3264, n3283, WX3262, n3284,
         WX3260, WX3258, WX3256, WX3254, WX3252, WX3250, WX3248, WX3246,
         WX3244, WX3242, WX3240, WX3238, WX3236, WX3234, WX3232, WX3230,
         WX3132, WX3130, WX3128, WX3126, WX3124, WX3122, WX3120, WX3118,
         WX3116, WX3114, WX3112, WX3110, WX3108, WX3106, WX3104, WX3102,
         WX3100, WX3098, WX3096, WX3094, WX3092, WX3090, WX3088, WX3086,
         WX3084, WX3082, WX3080, WX3078, WX3076, WX3074, WX3072, WX3070,
         WX2619, WX2617, WX2615, WX2613, WX2611, WX2609, WX2607, WX2605,
         WX2603, WX2601, WX2599, WX2597, WX2595, WX2593, WX2591, WX2589,
         WX2587, WX2585, WX2583, WX2581, WX2579, WX2577, WX2575, WX2573,
         WX2571, WX2569, WX2567, WX2565, WX2563, WX2561, WX2559, WX2557,
         WX2191, WX2189, WX2187, WX2185, WX2183, WX2181, WX2179, WX2177,
         WX2175, WX2173, WX2171, WX2169, WX2167, WX2165, WX2163, WX2161,
         WX2159, WX2157, WX2155, WX2153, WX2151, WX2149, WX2147, WX2145,
         WX2143, WX2141, WX2139, WX2137, WX2135, WX2133, WX2131, WX2129,
         WX2127, WX2125, WX2123, WX2121, WX2119, WX2117, WX2115, WX2113,
         WX2111, WX2109, WX2107, WX2105, WX2103, WX2101, WX2099, WX2097,
         WX2095, WX2093, WX2091, WX2089, WX2087, WX2085, WX2083, WX2081,
         WX2079, WX2077, WX2075, WX2073, WX2071, WX2069, WX2067, WX2065,
         WX2063, WX2061, WX2059, WX2057, WX2055, WX2053, WX2051, WX2049,
         WX2047, WX2045, WX2043, WX2041, WX2039, WX2037, WX2035, WX2033,
         WX2031, WX2029, WX2027, WX2025, WX2023, WX2021, WX2019, WX2017,
         WX2015, WX2013, WX2011, WX2009, WX2007, WX2005, WX2003, WX2001,
         WX1999, n3285, n3286, WX1997, n3287, n3288, WX1995, n3289, n3290,
         WX1993, n3291, n3292, WX1991, n3293, n3294, WX1989, n3295, n3296,
         WX1987, n3297, n3298, WX1985, n3299, n3300, WX1983, n3301, n3302,
         WX1981, n3303, n3304, WX1979, n3305, n3306, WX1977, n3307, n3308,
         WX1975, n3309, n3310, WX1973, n3311, n3312, WX1971, n3313, n3314,
         WX1969, n3315, n3316, WX1967, WX1965, WX1963, WX1961, WX1959, WX1957,
         WX1955, WX1953, WX1951, WX1949, WX1947, WX1945, WX1943, WX1941,
         WX1939, WX1937, WX1839, WX1837, WX1835, WX1833, WX1831, WX1829,
         WX1827, WX1825, WX1823, WX1821, WX1819, WX1817, WX1815, WX1813,
         WX1811, WX1809, WX1807, WX1805, WX1803, WX1801, WX1799, WX1797,
         WX1795, WX1793, WX1791, WX1789, WX1787, WX1785, WX1783, WX1781,
         WX1779, WX1777, WX1326, WX1324, WX1322, WX1320, WX1318, WX1316,
         WX1314, WX1312, WX1310, WX1308, WX1306, WX1304, WX1302, WX1300,
         WX1298, WX1296, WX1294, WX1292, WX1290, WX1288, WX1286, WX1284,
         WX1282, WX1280, WX1278, WX1276, WX1274, WX1272, WX1270, WX1268,
         WX1266, WX1264, WX11670, WX11668, WX11666, WX11664, WX11662, WX11660,
         WX11658, WX11656, WX11654, WX11652, WX11650, WX11648, WX11646,
         WX11644, WX11642, WX11640, WX11638, WX11636, WX11634, WX11632,
         WX11630, WX11628, WX11626, WX11624, WX11622, WX11620, WX11618,
         WX11616, WX11614, WX11612, WX11610, WX11608, WX11242, WX11240,
         WX11238, WX11236, WX11234, WX11232, WX11230, WX11228, WX11226,
         WX11224, WX11222, WX11220, WX11218, WX11216, WX11214, WX11212,
         WX11210, WX11208, WX11206, WX11204, WX11202, WX11200, WX11198,
         WX11196, WX11194, WX11192, WX11190, WX11188, WX11186, WX11184,
         WX11182, WX11180, WX11178, WX11176, WX11174, WX11172, WX11170,
         WX11168, WX11166, WX11164, WX11162, WX11160, WX11158, WX11156,
         WX11154, WX11152, WX11150, WX11148, WX11146, WX11144, WX11142,
         WX11140, WX11138, WX11136, WX11134, WX11132, WX11130, WX11128,
         WX11126, WX11124, WX11122, WX11120, WX11118, WX11116, WX11114,
         WX11112, WX11110, WX11108, WX11106, WX11104, WX11102, WX11100,
         WX11098, WX11096, WX11094, WX11092, WX11090, WX11088, WX11086,
         WX11084, WX11082, WX11080, WX11078, WX11076, WX11074, WX11072,
         WX11070, WX11068, WX11066, WX11064, WX11062, WX11060, WX11058,
         WX11056, WX11054, WX11052, WX11050, n3317, WX11048, n3318, WX11046,
         n3319, WX11044, n3320, WX11042, n3321, WX11040, n3322, WX11038, n3323,
         WX11036, n3324, WX11034, n3325, WX11032, n3326, WX11030, n3327,
         WX11028, n3328, WX11026, n3329, WX11024, n3330, WX11022, n3331,
         WX11020, n3332, WX11018, WX11016, WX11014, WX11012, WX11010, WX11008,
         WX11006, WX11004, WX11002, WX11000, WX10998, WX10996, WX10994,
         WX10992, WX10990, WX10988, WX10890, WX10888, WX10886, WX10884,
         WX10882, WX10880, WX10878, WX10876, WX10874, WX10872, WX10870,
         WX10868, WX10866, WX10864, WX10862, WX10860, WX10858, WX10856,
         WX10854, WX10852, WX10850, WX10848, WX10846, WX10844, WX10842,
         WX10840, WX10838, WX10836, WX10834, WX10832, WX10830, WX10828,
         WX10377, WX10375, WX10373, WX10371, WX10369, WX10367, WX10365,
         WX10363, WX10361, WX10359, WX10357, WX10355, WX10353, WX10351,
         WX10349, WX10347, WX10345, WX10343, WX10341, WX10339, WX10337,
         WX10335, WX10333, WX10331, WX10329, WX10327, WX10325, WX10323,
         WX10321, WX10319, WX10317, WX10315, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994;

wire Trojan_out0,  troj11_0counter_0_,  troj11_0N1,  troj11_0N2,  troj11_0N3,  troj11_0N6,  troj11_0n1,  troj11_0n2,  troj11_0n3,  troj11_0n4,  troj11_0n5,  troj11_0n6,  troj11_0n7,  troj11_0n8,  troj11_0n9,  troj11_0n10,  Trigger_en0_0,  trig32_0n1,  trig32_0n2,  trig32_0n3,  trig32_0n4,  tempWX4567;

  assign test_so = CRC_OUT_1_31;

  nor2s3 U1 ( .DIN1(n4997), .DIN2(n6725), .Q(WX9949) );
  nor2s3 U2 ( .DIN1(n5001), .DIN2(n6712), .Q(WX9947) );
  nor2s3 U3 ( .DIN1(n5005), .DIN2(n6745), .Q(WX9945) );
  nor2s3 U4 ( .DIN1(n5009), .DIN2(n6745), .Q(WX9943) );
  nor2s3 U5 ( .DIN1(n5013), .DIN2(n6745), .Q(WX9941) );
  nor2s3 U6 ( .DIN1(n5017), .DIN2(n6744), .Q(WX9939) );
  nor2s3 U7 ( .DIN1(n5021), .DIN2(n6744), .Q(WX9937) );
  nor2s3 U8 ( .DIN1(n5025), .DIN2(n6744), .Q(WX9935) );
  nor2s3 U9 ( .DIN1(n5029), .DIN2(n6744), .Q(WX9933) );
  nor2s3 U10 ( .DIN1(n5033), .DIN2(n6744), .Q(WX9931) );
  nor2s3 U11 ( .DIN1(n5037), .DIN2(n6744), .Q(WX9929) );
  nor2s3 U12 ( .DIN1(n5041), .DIN2(n6744), .Q(WX9927) );
  nor2s3 U13 ( .DIN1(n5045), .DIN2(n6744), .Q(WX9925) );
  nor2s3 U14 ( .DIN1(n5049), .DIN2(n6744), .Q(WX9923) );
  nor2s3 U15 ( .DIN1(n5053), .DIN2(n6744), .Q(WX9921) );
  nor2s3 U16 ( .DIN1(n5057), .DIN2(n6744), .Q(WX9919) );
  nor2s3 U17 ( .DIN1(n5061), .DIN2(n6744), .Q(WX9917) );
  nor2s3 U18 ( .DIN1(n5065), .DIN2(n6743), .Q(WX9915) );
  nor2s3 U19 ( .DIN1(n5069), .DIN2(n6743), .Q(WX9913) );
  nor2s3 U20 ( .DIN1(n5073), .DIN2(n6743), .Q(WX9911) );
  nor2s3 U21 ( .DIN1(n5077), .DIN2(n6743), .Q(WX9909) );
  nor2s3 U22 ( .DIN1(n5081), .DIN2(n6743), .Q(WX9907) );
  nor2s3 U23 ( .DIN1(n5085), .DIN2(n6743), .Q(WX9905) );
  nor2s3 U24 ( .DIN1(n5089), .DIN2(n6743), .Q(WX9903) );
  nor2s3 U25 ( .DIN1(n5093), .DIN2(n6743), .Q(WX9901) );
  nor2s3 U26 ( .DIN1(n5097), .DIN2(n6743), .Q(WX9899) );
  nor2s3 U27 ( .DIN1(n5101), .DIN2(n6743), .Q(WX9897) );
  nor2s3 U28 ( .DIN1(n5105), .DIN2(n6743), .Q(WX9895) );
  nor2s3 U29 ( .DIN1(n5109), .DIN2(n6743), .Q(WX9893) );
  nor2s3 U30 ( .DIN1(n5113), .DIN2(n6742), .Q(WX9891) );
  nor2s3 U31 ( .DIN1(n5117), .DIN2(n6742), .Q(WX9889) );
  nor2s3 U32 ( .DIN1(n5121), .DIN2(n6742), .Q(WX9887) );
  nor2s3 U33 ( .DIN1(n4996), .DIN2(n6742), .Q(WX9885) );
  nor2s3 U34 ( .DIN1(n5000), .DIN2(n6742), .Q(WX9883) );
  nor2s3 U35 ( .DIN1(n5004), .DIN2(n6742), .Q(WX9881) );
  nor2s3 U36 ( .DIN1(n5008), .DIN2(n6742), .Q(WX9879) );
  nor2s3 U37 ( .DIN1(n5012), .DIN2(n6742), .Q(WX9877) );
  nor2s3 U38 ( .DIN1(n5016), .DIN2(n6742), .Q(WX9875) );
  nor2s3 U39 ( .DIN1(n5020), .DIN2(n6742), .Q(WX9873) );
  nor2s3 U40 ( .DIN1(n5024), .DIN2(n6742), .Q(WX9871) );
  nor2s3 U41 ( .DIN1(n5028), .DIN2(n6742), .Q(WX9869) );
  nor2s3 U42 ( .DIN1(n5032), .DIN2(n6741), .Q(WX9867) );
  nor2s3 U43 ( .DIN1(n5036), .DIN2(n6741), .Q(WX9865) );
  nor2s3 U44 ( .DIN1(n5040), .DIN2(n6741), .Q(WX9863) );
  nor2s3 U45 ( .DIN1(n5044), .DIN2(n6741), .Q(WX9861) );
  nor2s3 U46 ( .DIN1(n5048), .DIN2(n6741), .Q(WX9859) );
  nor2s3 U47 ( .DIN1(n5052), .DIN2(n6741), .Q(WX9857) );
  nor2s3 U48 ( .DIN1(n5056), .DIN2(n6741), .Q(WX9855) );
  and2s3 U49 ( .DIN1(RESET), .DIN2(n5060), .Q(WX9853) );
  and2s3 U50 ( .DIN1(RESET), .DIN2(n5064), .Q(WX9851) );
  and2s3 U51 ( .DIN1(RESET), .DIN2(n5068), .Q(WX9849) );
  and2s3 U52 ( .DIN1(RESET), .DIN2(n5072), .Q(WX9847) );
  and2s3 U53 ( .DIN1(RESET), .DIN2(n5076), .Q(WX9845) );
  and2s3 U54 ( .DIN1(RESET), .DIN2(n5080), .Q(WX9843) );
  and2s3 U55 ( .DIN1(RESET), .DIN2(n5084), .Q(WX9841) );
  and2s3 U56 ( .DIN1(RESET), .DIN2(n5088), .Q(WX9839) );
  and2s3 U57 ( .DIN1(RESET), .DIN2(n5092), .Q(WX9837) );
  and2s3 U58 ( .DIN1(RESET), .DIN2(n5096), .Q(WX9835) );
  and2s3 U59 ( .DIN1(RESET), .DIN2(n5100), .Q(WX9833) );
  and2s3 U60 ( .DIN1(RESET), .DIN2(n5104), .Q(WX9831) );
  and2s3 U61 ( .DIN1(RESET), .DIN2(n5108), .Q(WX9829) );
  and2s3 U62 ( .DIN1(RESET), .DIN2(n5112), .Q(WX9827) );
  and2s3 U63 ( .DIN1(RESET), .DIN2(n5116), .Q(WX9825) );
  and2s3 U64 ( .DIN1(RESET), .DIN2(n5120), .Q(WX9823) );
  and2s3 U65 ( .DIN1(RESET), .DIN2(n4995), .Q(WX9821) );
  and2s3 U66 ( .DIN1(RESET), .DIN2(n4999), .Q(WX9819) );
  and2s3 U67 ( .DIN1(RESET), .DIN2(n5003), .Q(WX9817) );
  and2s3 U68 ( .DIN1(RESET), .DIN2(n5007), .Q(WX9815) );
  and2s3 U69 ( .DIN1(RESET), .DIN2(n5011), .Q(WX9813) );
  and2s3 U70 ( .DIN1(RESET), .DIN2(n5015), .Q(WX9811) );
  and2s3 U71 ( .DIN1(RESET), .DIN2(n5019), .Q(WX9809) );
  and2s3 U72 ( .DIN1(RESET), .DIN2(n5023), .Q(WX9807) );
  and2s3 U73 ( .DIN1(RESET), .DIN2(n5027), .Q(WX9805) );
  and2s3 U74 ( .DIN1(RESET), .DIN2(n5031), .Q(WX9803) );
  and2s3 U75 ( .DIN1(RESET), .DIN2(n5035), .Q(WX9801) );
  and2s3 U76 ( .DIN1(RESET), .DIN2(n5039), .Q(WX9799) );
  and2s3 U77 ( .DIN1(RESET), .DIN2(n5043), .Q(WX9797) );
  and2s3 U78 ( .DIN1(RESET), .DIN2(n5047), .Q(WX9795) );
  and2s3 U79 ( .DIN1(RESET), .DIN2(n5051), .Q(WX9793) );
  and2s3 U80 ( .DIN1(RESET), .DIN2(n5055), .Q(WX9791) );
  nor2s3 U81 ( .DIN1(n5059), .DIN2(n6741), .Q(WX9789) );
  nor2s3 U82 ( .DIN1(n5063), .DIN2(n6741), .Q(WX9787) );
  nor2s3 U83 ( .DIN1(n5067), .DIN2(n6741), .Q(WX9785) );
  nor2s3 U84 ( .DIN1(n5071), .DIN2(n6741), .Q(WX9783) );
  nor2s3 U85 ( .DIN1(n5075), .DIN2(n6741), .Q(WX9781) );
  nor2s3 U86 ( .DIN1(n5079), .DIN2(n6740), .Q(WX9779) );
  nor2s3 U87 ( .DIN1(n5083), .DIN2(n6740), .Q(WX9777) );
  nor2s3 U88 ( .DIN1(n5087), .DIN2(n6740), .Q(WX9775) );
  nor2s3 U89 ( .DIN1(n5091), .DIN2(n6740), .Q(WX9773) );
  nor2s3 U90 ( .DIN1(n5095), .DIN2(n6740), .Q(WX9771) );
  nor2s3 U91 ( .DIN1(n5099), .DIN2(n6740), .Q(WX9769) );
  nor2s3 U92 ( .DIN1(n5103), .DIN2(n6740), .Q(WX9767) );
  nor2s3 U93 ( .DIN1(n5107), .DIN2(n6740), .Q(WX9765) );
  nor2s3 U94 ( .DIN1(n5111), .DIN2(n6740), .Q(WX9763) );
  nor2s3 U95 ( .DIN1(n5115), .DIN2(n6740), .Q(WX9761) );
  nor2s3 U96 ( .DIN1(n5119), .DIN2(n6740), .Q(WX9759) );
  nnd4s2 U97 ( .DIN1(n2308), .DIN2(n2309), .DIN3(n2310), .DIN4(n2311), .Q(
        WX9757) );
  nnd2s3 U98 ( .DIN1(n6657), .DIN2(n2313), .Q(n2311) );
  nnd2s3 U99 ( .DIN1(n6625), .DIN2(n2315), .Q(n2310) );
  nnd2s3 U100 ( .DIN1(n6616), .DIN2(n1825), .Q(n2309) );
  nnd2s3 U101 ( .DIN1(n6585), .DIN2(n1824), .Q(n2308) );
  nnd4s2 U102 ( .DIN1(n2318), .DIN2(n2319), .DIN3(n2320), .DIN4(n2321), .Q(
        WX9755) );
  nnd2s3 U103 ( .DIN1(n2322), .DIN2(n6667), .Q(n2321) );
  nnd2s3 U104 ( .DIN1(n2323), .DIN2(n6636), .Q(n2320) );
  nnd2s3 U105 ( .DIN1(n6616), .DIN2(n1826), .Q(n2319) );
  nnd2s3 U106 ( .DIN1(n6585), .DIN2(n1823), .Q(n2318) );
  nnd4s2 U107 ( .DIN1(n2324), .DIN2(n2325), .DIN3(n2326), .DIN4(n2327), .Q(
        WX9753) );
  nnd2s3 U108 ( .DIN1(n2328), .DIN2(n6666), .Q(n2327) );
  nnd2s3 U109 ( .DIN1(n2329), .DIN2(n6635), .Q(n2326) );
  nnd2s3 U110 ( .DIN1(n6615), .DIN2(n1827), .Q(n2325) );
  nnd2s3 U111 ( .DIN1(n6584), .DIN2(n1822), .Q(n2324) );
  nnd4s2 U112 ( .DIN1(n2330), .DIN2(n2331), .DIN3(n2332), .DIN4(n2333), .Q(
        WX9751) );
  nnd2s3 U113 ( .DIN1(n2334), .DIN2(n6666), .Q(n2333) );
  nnd2s3 U114 ( .DIN1(n2335), .DIN2(n6635), .Q(n2332) );
  nnd2s3 U115 ( .DIN1(n6615), .DIN2(n1828), .Q(n2331) );
  nnd2s3 U116 ( .DIN1(n6584), .DIN2(n1821), .Q(n2330) );
  nnd4s2 U117 ( .DIN1(n2336), .DIN2(n2337), .DIN3(n2338), .DIN4(n2339), .Q(
        WX9749) );
  nnd2s3 U118 ( .DIN1(n2340), .DIN2(n6666), .Q(n2339) );
  nnd2s3 U119 ( .DIN1(n2341), .DIN2(n6635), .Q(n2338) );
  nnd2s3 U120 ( .DIN1(n6615), .DIN2(n1829), .Q(n2337) );
  nnd2s3 U121 ( .DIN1(n6584), .DIN2(n1820), .Q(n2336) );
  nnd4s2 U122 ( .DIN1(n2342), .DIN2(n2343), .DIN3(n2344), .DIN4(n2345), .Q(
        WX9747) );
  nnd2s3 U123 ( .DIN1(n2346), .DIN2(n6666), .Q(n2345) );
  nnd2s3 U124 ( .DIN1(n2347), .DIN2(n6635), .Q(n2344) );
  nnd2s3 U125 ( .DIN1(n6615), .DIN2(n1830), .Q(n2343) );
  nnd2s3 U126 ( .DIN1(n6584), .DIN2(n1819), .Q(n2342) );
  nnd4s2 U127 ( .DIN1(n2348), .DIN2(n2349), .DIN3(n2350), .DIN4(n2351), .Q(
        WX9745) );
  nnd2s3 U128 ( .DIN1(n2352), .DIN2(n6666), .Q(n2351) );
  nnd2s3 U129 ( .DIN1(n2353), .DIN2(n6635), .Q(n2350) );
  nnd2s3 U130 ( .DIN1(n6615), .DIN2(n1831), .Q(n2349) );
  nnd2s3 U131 ( .DIN1(n6584), .DIN2(n1818), .Q(n2348) );
  nnd4s2 U132 ( .DIN1(n2354), .DIN2(n2355), .DIN3(n2356), .DIN4(n2357), .Q(
        WX9743) );
  nnd2s3 U133 ( .DIN1(n2358), .DIN2(n6666), .Q(n2357) );
  nnd2s3 U134 ( .DIN1(n2359), .DIN2(n6635), .Q(n2356) );
  nnd2s3 U135 ( .DIN1(n6615), .DIN2(n1832), .Q(n2355) );
  nnd2s3 U136 ( .DIN1(n6584), .DIN2(n1817), .Q(n2354) );
  nnd4s2 U137 ( .DIN1(n2360), .DIN2(n2361), .DIN3(n2362), .DIN4(n2363), .Q(
        WX9741) );
  nnd2s3 U138 ( .DIN1(n2364), .DIN2(n6666), .Q(n2363) );
  nnd2s3 U139 ( .DIN1(n2365), .DIN2(n6635), .Q(n2362) );
  nnd2s3 U140 ( .DIN1(n6615), .DIN2(n1833), .Q(n2361) );
  nnd2s3 U141 ( .DIN1(n6584), .DIN2(n1816), .Q(n2360) );
  nnd4s2 U142 ( .DIN1(n2366), .DIN2(n2367), .DIN3(n2368), .DIN4(n2369), .Q(
        WX9739) );
  nnd2s3 U143 ( .DIN1(n2370), .DIN2(n6666), .Q(n2369) );
  nnd2s3 U144 ( .DIN1(n2371), .DIN2(n6635), .Q(n2368) );
  nnd2s3 U145 ( .DIN1(n6615), .DIN2(n1834), .Q(n2367) );
  nnd2s3 U146 ( .DIN1(n6584), .DIN2(n1815), .Q(n2366) );
  nnd4s2 U147 ( .DIN1(n2372), .DIN2(n2373), .DIN3(n2374), .DIN4(n2375), .Q(
        WX9737) );
  nnd2s3 U148 ( .DIN1(n2376), .DIN2(n6666), .Q(n2375) );
  nnd2s3 U149 ( .DIN1(n2377), .DIN2(n6635), .Q(n2374) );
  nnd2s3 U150 ( .DIN1(n6615), .DIN2(n1835), .Q(n2373) );
  nnd2s3 U151 ( .DIN1(n6584), .DIN2(n1814), .Q(n2372) );
  nnd4s2 U152 ( .DIN1(n2378), .DIN2(n2379), .DIN3(n2380), .DIN4(n2381), .Q(
        WX9735) );
  nnd2s3 U153 ( .DIN1(n2382), .DIN2(n6666), .Q(n2381) );
  nnd2s3 U154 ( .DIN1(n2383), .DIN2(n6635), .Q(n2380) );
  nnd2s3 U155 ( .DIN1(n6615), .DIN2(n1836), .Q(n2379) );
  nnd2s3 U156 ( .DIN1(n6584), .DIN2(n1813), .Q(n2378) );
  nnd4s2 U157 ( .DIN1(n2384), .DIN2(n2385), .DIN3(n2386), .DIN4(n2387), .Q(
        WX9733) );
  nnd2s3 U158 ( .DIN1(n2388), .DIN2(n6666), .Q(n2387) );
  nnd2s3 U159 ( .DIN1(n2389), .DIN2(n6635), .Q(n2386) );
  nnd2s3 U160 ( .DIN1(n6615), .DIN2(n1837), .Q(n2385) );
  nnd2s3 U161 ( .DIN1(n6584), .DIN2(n1812), .Q(n2384) );
  nnd4s2 U162 ( .DIN1(n2390), .DIN2(n2391), .DIN3(n2392), .DIN4(n2393), .Q(
        WX9731) );
  nnd2s3 U163 ( .DIN1(n2394), .DIN2(n6666), .Q(n2393) );
  nnd2s3 U164 ( .DIN1(n2395), .DIN2(n6635), .Q(n2392) );
  nnd2s3 U165 ( .DIN1(n6615), .DIN2(n1838), .Q(n2391) );
  nnd2s3 U166 ( .DIN1(n6584), .DIN2(n1811), .Q(n2390) );
  nnd4s2 U167 ( .DIN1(n2396), .DIN2(n2397), .DIN3(n2398), .DIN4(n2399), .Q(
        WX9729) );
  nnd2s3 U168 ( .DIN1(n2400), .DIN2(n6666), .Q(n2399) );
  nnd2s3 U169 ( .DIN1(n2401), .DIN2(n6635), .Q(n2398) );
  nnd2s3 U170 ( .DIN1(n6615), .DIN2(n1839), .Q(n2397) );
  nnd2s3 U171 ( .DIN1(n6584), .DIN2(n1810), .Q(n2396) );
  nnd4s2 U172 ( .DIN1(n2402), .DIN2(n2403), .DIN3(n2404), .DIN4(n2405), .Q(
        WX9727) );
  nnd2s3 U173 ( .DIN1(n2406), .DIN2(n6665), .Q(n2405) );
  nnd2s3 U174 ( .DIN1(n2407), .DIN2(n6634), .Q(n2404) );
  nnd2s3 U175 ( .DIN1(n6614), .DIN2(n1840), .Q(n2403) );
  nnd2s3 U176 ( .DIN1(n6583), .DIN2(n1809), .Q(n2402) );
  nnd4s2 U177 ( .DIN1(n2408), .DIN2(n2409), .DIN3(n2410), .DIN4(n2411), .Q(
        WX9725) );
  nnd2s3 U178 ( .DIN1(n2412), .DIN2(n6665), .Q(n2411) );
  nnd2s3 U179 ( .DIN1(n2413), .DIN2(n6634), .Q(n2410) );
  nnd2s3 U180 ( .DIN1(n6614), .DIN2(n1841), .Q(n2409) );
  nnd2s3 U181 ( .DIN1(n6583), .DIN2(n1808), .Q(n2408) );
  nnd4s2 U182 ( .DIN1(n2414), .DIN2(n2415), .DIN3(n2416), .DIN4(n2417), .Q(
        WX9723) );
  nnd2s3 U183 ( .DIN1(n2418), .DIN2(n6665), .Q(n2417) );
  nnd2s3 U184 ( .DIN1(n2419), .DIN2(n6634), .Q(n2416) );
  nnd2s3 U185 ( .DIN1(n6614), .DIN2(n1842), .Q(n2415) );
  nnd2s3 U186 ( .DIN1(n6583), .DIN2(n1807), .Q(n2414) );
  nnd4s2 U187 ( .DIN1(n2420), .DIN2(n2421), .DIN3(n2422), .DIN4(n2423), .Q(
        WX9721) );
  nnd2s3 U188 ( .DIN1(n2424), .DIN2(n6665), .Q(n2423) );
  nnd2s3 U189 ( .DIN1(n2425), .DIN2(n6634), .Q(n2422) );
  nnd2s3 U190 ( .DIN1(n6614), .DIN2(n1843), .Q(n2421) );
  nnd2s3 U191 ( .DIN1(n6583), .DIN2(n1806), .Q(n2420) );
  nnd4s2 U192 ( .DIN1(n2426), .DIN2(n2427), .DIN3(n2428), .DIN4(n2429), .Q(
        WX9719) );
  nnd2s3 U193 ( .DIN1(n2430), .DIN2(n6665), .Q(n2429) );
  nnd2s3 U194 ( .DIN1(n2431), .DIN2(n6634), .Q(n2428) );
  nnd2s3 U195 ( .DIN1(n6614), .DIN2(n1844), .Q(n2427) );
  nnd2s3 U196 ( .DIN1(n6583), .DIN2(n1805), .Q(n2426) );
  nnd4s2 U197 ( .DIN1(n2432), .DIN2(n2433), .DIN3(n2434), .DIN4(n2435), .Q(
        WX9717) );
  nnd2s3 U198 ( .DIN1(n2436), .DIN2(n6665), .Q(n2435) );
  nnd2s3 U199 ( .DIN1(n2437), .DIN2(n6634), .Q(n2434) );
  nnd2s3 U200 ( .DIN1(n6614), .DIN2(n1845), .Q(n2433) );
  nnd2s3 U201 ( .DIN1(n6583), .DIN2(n1804), .Q(n2432) );
  nnd4s2 U202 ( .DIN1(n2438), .DIN2(n2439), .DIN3(n2440), .DIN4(n2441), .Q(
        WX9715) );
  nnd2s3 U203 ( .DIN1(n2442), .DIN2(n6665), .Q(n2441) );
  nnd2s3 U204 ( .DIN1(n2443), .DIN2(n6634), .Q(n2440) );
  nnd2s3 U205 ( .DIN1(n6614), .DIN2(n1846), .Q(n2439) );
  nnd2s3 U206 ( .DIN1(n6583), .DIN2(n1803), .Q(n2438) );
  nnd4s2 U207 ( .DIN1(n2444), .DIN2(n2445), .DIN3(n2446), .DIN4(n2447), .Q(
        WX9713) );
  nnd2s3 U208 ( .DIN1(n2448), .DIN2(n6665), .Q(n2447) );
  nnd2s3 U209 ( .DIN1(n2449), .DIN2(n6634), .Q(n2446) );
  nnd2s3 U210 ( .DIN1(n6614), .DIN2(n1847), .Q(n2445) );
  nnd2s3 U211 ( .DIN1(n6583), .DIN2(n1802), .Q(n2444) );
  nnd4s2 U212 ( .DIN1(n2450), .DIN2(n2451), .DIN3(n2452), .DIN4(n2453), .Q(
        WX9711) );
  nnd2s3 U213 ( .DIN1(n2454), .DIN2(n6665), .Q(n2453) );
  nnd2s3 U214 ( .DIN1(n2455), .DIN2(n6634), .Q(n2452) );
  nnd2s3 U215 ( .DIN1(n6614), .DIN2(n1848), .Q(n2451) );
  nnd2s3 U216 ( .DIN1(n6583), .DIN2(n1801), .Q(n2450) );
  nnd4s2 U217 ( .DIN1(n2456), .DIN2(n2457), .DIN3(n2458), .DIN4(n2459), .Q(
        WX9709) );
  nnd2s3 U218 ( .DIN1(n2460), .DIN2(n6665), .Q(n2459) );
  nnd2s3 U219 ( .DIN1(n2461), .DIN2(n6634), .Q(n2458) );
  nnd2s3 U220 ( .DIN1(n6614), .DIN2(n1849), .Q(n2457) );
  nnd2s3 U221 ( .DIN1(n6583), .DIN2(n1800), .Q(n2456) );
  nnd4s2 U222 ( .DIN1(n2462), .DIN2(n2463), .DIN3(n2464), .DIN4(n2465), .Q(
        WX9707) );
  nnd2s3 U223 ( .DIN1(n2466), .DIN2(n6665), .Q(n2465) );
  nnd2s3 U224 ( .DIN1(n2467), .DIN2(n6634), .Q(n2464) );
  nnd2s3 U225 ( .DIN1(n6614), .DIN2(n1850), .Q(n2463) );
  nnd2s3 U226 ( .DIN1(n6583), .DIN2(n1799), .Q(n2462) );
  nnd4s2 U227 ( .DIN1(n2468), .DIN2(n2469), .DIN3(n2470), .DIN4(n2471), .Q(
        WX9705) );
  nnd2s3 U228 ( .DIN1(n2472), .DIN2(n6665), .Q(n2471) );
  nnd2s3 U229 ( .DIN1(n2473), .DIN2(n6634), .Q(n2470) );
  nnd2s3 U230 ( .DIN1(n6614), .DIN2(n1851), .Q(n2469) );
  nnd2s3 U231 ( .DIN1(n6583), .DIN2(n1798), .Q(n2468) );
  nnd4s2 U232 ( .DIN1(n2474), .DIN2(n2475), .DIN3(n2476), .DIN4(n2477), .Q(
        WX9703) );
  nnd2s3 U233 ( .DIN1(n2478), .DIN2(n6665), .Q(n2477) );
  nnd2s3 U234 ( .DIN1(n2479), .DIN2(n6634), .Q(n2476) );
  nnd2s3 U235 ( .DIN1(n6614), .DIN2(n1852), .Q(n2475) );
  nnd2s3 U236 ( .DIN1(n6583), .DIN2(n1797), .Q(n2474) );
  nnd4s2 U237 ( .DIN1(n2480), .DIN2(n2481), .DIN3(n2482), .DIN4(n2483), .Q(
        WX9701) );
  nnd2s3 U238 ( .DIN1(n2484), .DIN2(n6664), .Q(n2483) );
  nnd2s3 U239 ( .DIN1(n2485), .DIN2(n6633), .Q(n2482) );
  nnd2s3 U240 ( .DIN1(n6613), .DIN2(n1853), .Q(n2481) );
  nnd2s3 U241 ( .DIN1(n6582), .DIN2(n1796), .Q(n2480) );
  nnd4s2 U242 ( .DIN1(n2486), .DIN2(n2487), .DIN3(n2488), .DIN4(n2489), .Q(
        WX9699) );
  nnd2s3 U243 ( .DIN1(n2490), .DIN2(n6664), .Q(n2489) );
  nnd2s3 U244 ( .DIN1(n2491), .DIN2(n6633), .Q(n2488) );
  nnd2s3 U245 ( .DIN1(n6613), .DIN2(n1854), .Q(n2487) );
  nnd2s3 U246 ( .DIN1(n6582), .DIN2(n1795), .Q(n2486) );
  nnd4s2 U247 ( .DIN1(n2492), .DIN2(n2493), .DIN3(n2494), .DIN4(n2495), .Q(
        WX9697) );
  nnd2s3 U248 ( .DIN1(n2496), .DIN2(n6664), .Q(n2495) );
  nnd2s3 U249 ( .DIN1(n2497), .DIN2(n6633), .Q(n2494) );
  nnd2s3 U250 ( .DIN1(n6613), .DIN2(n1855), .Q(n2493) );
  nnd2s3 U251 ( .DIN1(n6582), .DIN2(n1794), .Q(n2492) );
  nnd4s2 U252 ( .DIN1(n2498), .DIN2(n2499), .DIN3(n2500), .DIN4(n2501), .Q(
        WX9695) );
  nnd2s3 U253 ( .DIN1(n2502), .DIN2(n6664), .Q(n2501) );
  nnd2s3 U254 ( .DIN1(n6613), .DIN2(n1856), .Q(n2500) );
  nnd2s3 U255 ( .DIN1(n2503), .DIN2(n6633), .Q(n2499) );
  nnd2s3 U256 ( .DIN1(n6582), .DIN2(n1793), .Q(n2498) );
  nor2s3 U257 ( .DIN1(n6789), .DIN2(n1856), .Q(WX9597) );
  nor2s3 U258 ( .DIN1(n4964), .DIN2(n6740), .Q(WX9595) );
  nor2s3 U259 ( .DIN1(n4965), .DIN2(n6739), .Q(WX9593) );
  nor2s3 U260 ( .DIN1(n4966), .DIN2(n6739), .Q(WX9591) );
  nor2s3 U261 ( .DIN1(n4967), .DIN2(n6739), .Q(WX9589) );
  nor2s3 U262 ( .DIN1(n4968), .DIN2(n6739), .Q(WX9587) );
  nor2s3 U263 ( .DIN1(n4969), .DIN2(n6739), .Q(WX9585) );
  nor2s3 U264 ( .DIN1(n4970), .DIN2(n6739), .Q(WX9583) );
  nor2s3 U265 ( .DIN1(n4971), .DIN2(n6739), .Q(WX9581) );
  nor2s3 U266 ( .DIN1(n4972), .DIN2(n6739), .Q(WX9579) );
  nor2s3 U267 ( .DIN1(n4973), .DIN2(n6739), .Q(WX9577) );
  nor2s3 U268 ( .DIN1(n4974), .DIN2(n6739), .Q(WX9575) );
  nor2s3 U269 ( .DIN1(n4975), .DIN2(n6739), .Q(WX9573) );
  nor2s3 U270 ( .DIN1(n4976), .DIN2(n6738), .Q(WX9571) );
  nor2s3 U271 ( .DIN1(n4977), .DIN2(n6738), .Q(WX9569) );
  nor2s3 U272 ( .DIN1(n4978), .DIN2(n6738), .Q(WX9567) );
  nor2s3 U273 ( .DIN1(n4979), .DIN2(n6738), .Q(WX9565) );
  nor2s3 U274 ( .DIN1(n4980), .DIN2(n6738), .Q(WX9563) );
  nor2s3 U275 ( .DIN1(n4981), .DIN2(n6738), .Q(WX9561) );
  nor2s3 U276 ( .DIN1(n4982), .DIN2(n6738), .Q(WX9559) );
  nor2s3 U277 ( .DIN1(n4983), .DIN2(n6738), .Q(WX9557) );
  nor2s3 U278 ( .DIN1(n4984), .DIN2(n6738), .Q(WX9555) );
  nor2s3 U279 ( .DIN1(n4985), .DIN2(n6738), .Q(WX9553) );
  nor2s3 U280 ( .DIN1(n4986), .DIN2(n6738), .Q(WX9551) );
  nor2s3 U281 ( .DIN1(n4987), .DIN2(n6738), .Q(WX9549) );
  nor2s3 U282 ( .DIN1(n4988), .DIN2(n6737), .Q(WX9547) );
  nor2s3 U283 ( .DIN1(n4989), .DIN2(n6737), .Q(WX9545) );
  nor2s3 U284 ( .DIN1(n4990), .DIN2(n6737), .Q(WX9543) );
  nor2s3 U285 ( .DIN1(n4991), .DIN2(n6737), .Q(WX9541) );
  nor2s3 U286 ( .DIN1(n4992), .DIN2(n6737), .Q(WX9539) );
  nor2s3 U287 ( .DIN1(n4993), .DIN2(n6737), .Q(WX9537) );
  nor2s3 U288 ( .DIN1(n4994), .DIN2(n6737), .Q(WX9535) );
  nor2s3 U289 ( .DIN1(n6793), .DIN2(n2504), .Q(WX9084) );
  xor2s3 U290 ( .DIN1(n5118), .DIN2(n5297), .Q(n2504) );
  nor2s3 U291 ( .DIN1(n6793), .DIN2(n2505), .Q(WX9082) );
  xor2s3 U292 ( .DIN1(n5114), .DIN2(n5292), .Q(n2505) );
  nor2s3 U293 ( .DIN1(n6793), .DIN2(n2506), .Q(WX9080) );
  xor2s3 U294 ( .DIN1(n5110), .DIN2(n5287), .Q(n2506) );
  nor2s3 U295 ( .DIN1(n6793), .DIN2(n2507), .Q(WX9078) );
  xor2s3 U296 ( .DIN1(n5106), .DIN2(n5282), .Q(n2507) );
  nor2s3 U297 ( .DIN1(n6793), .DIN2(n2508), .Q(WX9076) );
  xor2s3 U298 ( .DIN1(n5102), .DIN2(n5277), .Q(n2508) );
  nor2s3 U299 ( .DIN1(n6793), .DIN2(n2509), .Q(WX9074) );
  xor2s3 U300 ( .DIN1(n5098), .DIN2(n5272), .Q(n2509) );
  nor2s3 U301 ( .DIN1(n6793), .DIN2(n2510), .Q(WX9072) );
  xor2s3 U302 ( .DIN1(n5094), .DIN2(n5267), .Q(n2510) );
  nor2s3 U303 ( .DIN1(n6793), .DIN2(n2511), .Q(WX9070) );
  xor2s3 U304 ( .DIN1(n5090), .DIN2(n5262), .Q(n2511) );
  nor2s3 U305 ( .DIN1(n6793), .DIN2(n2512), .Q(WX9068) );
  xor2s3 U306 ( .DIN1(n5086), .DIN2(n5257), .Q(n2512) );
  nor2s3 U307 ( .DIN1(n6792), .DIN2(n2513), .Q(WX9066) );
  xor2s3 U308 ( .DIN1(n5082), .DIN2(n5252), .Q(n2513) );
  nor2s3 U309 ( .DIN1(n6792), .DIN2(n2514), .Q(WX9064) );
  xor2s3 U310 ( .DIN1(n5078), .DIN2(n5247), .Q(n2514) );
  nor2s3 U311 ( .DIN1(n6792), .DIN2(n2515), .Q(WX9062) );
  xor2s3 U312 ( .DIN1(n5074), .DIN2(n5242), .Q(n2515) );
  nor2s3 U313 ( .DIN1(n6792), .DIN2(n2516), .Q(WX9060) );
  xor2s3 U314 ( .DIN1(n5070), .DIN2(n5237), .Q(n2516) );
  nor2s3 U315 ( .DIN1(n6792), .DIN2(n2517), .Q(WX9058) );
  xor2s3 U316 ( .DIN1(n5066), .DIN2(n5232), .Q(n2517) );
  nor2s3 U317 ( .DIN1(n6792), .DIN2(n2518), .Q(WX9056) );
  xor2s3 U318 ( .DIN1(n5062), .DIN2(n5227), .Q(n2518) );
  nor2s3 U319 ( .DIN1(n2519), .DIN2(n6737), .Q(WX9054) );
  xnr2s3 U320 ( .DIN1(n5222), .DIN2(n2520), .Q(n2519) );
  xor2s3 U321 ( .DIN1(n5058), .DIN2(n5122), .Q(n2520) );
  nor2s3 U322 ( .DIN1(n6792), .DIN2(n2521), .Q(WX9052) );
  xor2s3 U323 ( .DIN1(n5054), .DIN2(n3236), .Q(n2521) );
  nor2s3 U324 ( .DIN1(n6792), .DIN2(n2522), .Q(WX9050) );
  xor2s3 U325 ( .DIN1(n5050), .DIN2(n3235), .Q(n2522) );
  nor2s3 U326 ( .DIN1(n6792), .DIN2(n2523), .Q(WX9048) );
  xor2s3 U327 ( .DIN1(n5046), .DIN2(n3234), .Q(n2523) );
  nor2s3 U328 ( .DIN1(n6792), .DIN2(n2524), .Q(WX9046) );
  xor2s3 U329 ( .DIN1(n5042), .DIN2(n3233), .Q(n2524) );
  nor2s3 U330 ( .DIN1(n2525), .DIN2(n6737), .Q(WX9044) );
  xnr2s3 U331 ( .DIN1(n3232), .DIN2(n2526), .Q(n2525) );
  xor2s3 U332 ( .DIN1(n5038), .DIN2(n5122), .Q(n2526) );
  nor2s3 U333 ( .DIN1(n6792), .DIN2(n2527), .Q(WX9042) );
  xor2s3 U334 ( .DIN1(n5034), .DIN2(n3231), .Q(n2527) );
  nor2s3 U335 ( .DIN1(n6791), .DIN2(n2528), .Q(WX9040) );
  xor2s3 U336 ( .DIN1(n5030), .DIN2(n3230), .Q(n2528) );
  nor2s3 U337 ( .DIN1(n6791), .DIN2(n2529), .Q(WX9038) );
  xor2s3 U338 ( .DIN1(n5026), .DIN2(n3229), .Q(n2529) );
  nor2s3 U339 ( .DIN1(n6791), .DIN2(n2530), .Q(WX9036) );
  xor2s3 U340 ( .DIN1(n5022), .DIN2(n3228), .Q(n2530) );
  nor2s3 U341 ( .DIN1(n6790), .DIN2(n2531), .Q(WX9034) );
  xor2s3 U342 ( .DIN1(n5018), .DIN2(n3227), .Q(n2531) );
  nor2s3 U343 ( .DIN1(n6790), .DIN2(n2532), .Q(WX9032) );
  xor2s3 U344 ( .DIN1(n5014), .DIN2(n3226), .Q(n2532) );
  nor2s3 U345 ( .DIN1(n2533), .DIN2(n6737), .Q(WX9030) );
  xnr2s3 U346 ( .DIN1(n3225), .DIN2(n2534), .Q(n2533) );
  xor2s3 U347 ( .DIN1(n5010), .DIN2(n5122), .Q(n2534) );
  nor2s3 U348 ( .DIN1(n6790), .DIN2(n2535), .Q(WX9028) );
  xor2s3 U349 ( .DIN1(n5006), .DIN2(n3224), .Q(n2535) );
  nor2s3 U350 ( .DIN1(n6790), .DIN2(n2536), .Q(WX9026) );
  xor2s3 U351 ( .DIN1(n5002), .DIN2(n3223), .Q(n2536) );
  nor2s3 U352 ( .DIN1(n6790), .DIN2(n2537), .Q(WX9024) );
  xor2s3 U353 ( .DIN1(n4998), .DIN2(n3222), .Q(n2537) );
  nor2s3 U354 ( .DIN1(n6790), .DIN2(n2538), .Q(WX9022) );
  xor2s3 U355 ( .DIN1(n5122), .DIN2(n3221), .Q(n2538) );
  nor2s3 U356 ( .DIN1(n6463), .DIN2(n6737), .Q(WX898) );
  nor2s3 U357 ( .DIN1(n6527), .DIN2(n6737), .Q(WX896) );
  nor2s3 U358 ( .DIN1(n6436), .DIN2(n6736), .Q(WX894) );
  nor2s3 U359 ( .DIN1(n6469), .DIN2(n6736), .Q(WX892) );
  nor2s3 U360 ( .DIN1(n6472), .DIN2(n6736), .Q(WX890) );
  nor2s3 U361 ( .DIN1(n6460), .DIN2(n6736), .Q(WX888) );
  nor2s3 U362 ( .DIN1(n6442), .DIN2(n6736), .Q(WX886) );
  nor2s3 U363 ( .DIN1(n6466), .DIN2(n6736), .Q(WX884) );
  nor2s3 U364 ( .DIN1(n6454), .DIN2(n6736), .Q(WX882) );
  nor2s3 U365 ( .DIN1(n6504), .DIN2(n6736), .Q(WX880) );
  nor2s3 U366 ( .DIN1(n6451), .DIN2(n6736), .Q(WX878) );
  nor2s3 U367 ( .DIN1(n6445), .DIN2(n6736), .Q(WX876) );
  nor2s3 U368 ( .DIN1(n6457), .DIN2(n6736), .Q(WX874) );
  nor2s3 U369 ( .DIN1(n6448), .DIN2(n6736), .Q(WX872) );
  nor2s3 U370 ( .DIN1(n6523), .DIN2(n6735), .Q(WX870) );
  nor2s3 U371 ( .DIN1(n6439), .DIN2(n6735), .Q(WX868) );
  nor2s3 U372 ( .DIN1(n6539), .DIN2(n6735), .Q(WX866) );
  nor2s3 U373 ( .DIN1(n5157), .DIN2(n6735), .Q(WX8656) );
  nor2s3 U374 ( .DIN1(n5161), .DIN2(n6735), .Q(WX8654) );
  nor2s3 U375 ( .DIN1(n5165), .DIN2(n6735), .Q(WX8652) );
  nor2s3 U376 ( .DIN1(n5169), .DIN2(n6735), .Q(WX8650) );
  nor2s3 U377 ( .DIN1(n5173), .DIN2(n6735), .Q(WX8648) );
  nor2s3 U378 ( .DIN1(n5177), .DIN2(n6735), .Q(WX8646) );
  nor2s3 U379 ( .DIN1(n5181), .DIN2(n6735), .Q(WX8644) );
  nor2s3 U380 ( .DIN1(n5185), .DIN2(n6735), .Q(WX8642) );
  nor2s3 U381 ( .DIN1(n5189), .DIN2(n6735), .Q(WX8640) );
  nor2s3 U382 ( .DIN1(n6496), .DIN2(n6734), .Q(WX864) );
  nor2s3 U383 ( .DIN1(n5193), .DIN2(n6734), .Q(WX8638) );
  nor2s3 U384 ( .DIN1(n5197), .DIN2(n6734), .Q(WX8636) );
  nor2s3 U385 ( .DIN1(n5201), .DIN2(n6734), .Q(WX8634) );
  nor2s3 U386 ( .DIN1(n5205), .DIN2(n6734), .Q(WX8632) );
  nor2s3 U387 ( .DIN1(n5209), .DIN2(n6734), .Q(WX8630) );
  nor2s3 U388 ( .DIN1(n5213), .DIN2(n6734), .Q(WX8628) );
  nor2s3 U389 ( .DIN1(n5217), .DIN2(n6734), .Q(WX8626) );
  nor2s3 U390 ( .DIN1(n5221), .DIN2(n6734), .Q(WX8624) );
  nor2s3 U391 ( .DIN1(n5226), .DIN2(n6734), .Q(WX8622) );
  nor2s3 U392 ( .DIN1(n5231), .DIN2(n6739), .Q(WX8620) );
  nor2s3 U393 ( .DIN1(n6544), .DIN2(n6756), .Q(WX862) );
  nor2s3 U394 ( .DIN1(n5236), .DIN2(n6756), .Q(WX8618) );
  nor2s3 U395 ( .DIN1(n5241), .DIN2(n6756), .Q(WX8616) );
  nor2s3 U396 ( .DIN1(n5246), .DIN2(n6755), .Q(WX8614) );
  nor2s3 U397 ( .DIN1(n5251), .DIN2(n6755), .Q(WX8612) );
  nor2s3 U398 ( .DIN1(n5256), .DIN2(n6755), .Q(WX8610) );
  nor2s3 U399 ( .DIN1(n5261), .DIN2(n6755), .Q(WX8608) );
  nor2s3 U400 ( .DIN1(n5266), .DIN2(n6755), .Q(WX8606) );
  nor2s3 U401 ( .DIN1(n5271), .DIN2(n6755), .Q(WX8604) );
  nor2s3 U402 ( .DIN1(n5276), .DIN2(n6755), .Q(WX8602) );
  nor2s3 U403 ( .DIN1(n5281), .DIN2(n6755), .Q(WX8600) );
  nor2s3 U404 ( .DIN1(n6478), .DIN2(n6755), .Q(WX860) );
  nor2s3 U405 ( .DIN1(n5286), .DIN2(n6755), .Q(WX8598) );
  nor2s3 U406 ( .DIN1(n5291), .DIN2(n6755), .Q(WX8596) );
  nor2s3 U407 ( .DIN1(n5296), .DIN2(n6755), .Q(WX8594) );
  nor2s3 U408 ( .DIN1(n5156), .DIN2(n6754), .Q(WX8592) );
  nor2s3 U409 ( .DIN1(n5160), .DIN2(n6754), .Q(WX8590) );
  nor2s3 U410 ( .DIN1(n5164), .DIN2(n6754), .Q(WX8588) );
  nor2s3 U411 ( .DIN1(n5168), .DIN2(n6754), .Q(WX8586) );
  nor2s3 U412 ( .DIN1(n5172), .DIN2(n6754), .Q(WX8584) );
  nor2s3 U413 ( .DIN1(n5176), .DIN2(n6754), .Q(WX8582) );
  nor2s3 U414 ( .DIN1(n5180), .DIN2(n6754), .Q(WX8580) );
  nor2s3 U415 ( .DIN1(n6535), .DIN2(n6754), .Q(WX858) );
  nor2s3 U416 ( .DIN1(n5184), .DIN2(n6754), .Q(WX8578) );
  nor2s3 U417 ( .DIN1(n5188), .DIN2(n6754), .Q(WX8576) );
  nor2s3 U418 ( .DIN1(n5192), .DIN2(n6754), .Q(WX8574) );
  nor2s3 U419 ( .DIN1(n5196), .DIN2(n6754), .Q(WX8572) );
  nor2s3 U420 ( .DIN1(n5200), .DIN2(n6753), .Q(WX8570) );
  nor2s3 U421 ( .DIN1(n5204), .DIN2(n6753), .Q(WX8568) );
  nor2s3 U422 ( .DIN1(n5208), .DIN2(n6753), .Q(WX8566) );
  nor2s3 U423 ( .DIN1(n5212), .DIN2(n6753), .Q(WX8564) );
  nor2s3 U424 ( .DIN1(n5216), .DIN2(n6753), .Q(WX8562) );
  and2s3 U425 ( .DIN1(RESET), .DIN2(n5220), .Q(WX8560) );
  nor2s3 U426 ( .DIN1(n6518), .DIN2(n6753), .Q(WX856) );
  and2s3 U427 ( .DIN1(RESET), .DIN2(n5225), .Q(WX8558) );
  and2s3 U428 ( .DIN1(RESET), .DIN2(n5230), .Q(WX8556) );
  and2s3 U429 ( .DIN1(RESET), .DIN2(n5235), .Q(WX8554) );
  and2s3 U430 ( .DIN1(RESET), .DIN2(n5240), .Q(WX8552) );
  and2s3 U431 ( .DIN1(RESET), .DIN2(n5245), .Q(WX8550) );
  and2s3 U432 ( .DIN1(RESET), .DIN2(n5250), .Q(WX8548) );
  and2s3 U433 ( .DIN1(RESET), .DIN2(n5255), .Q(WX8546) );
  and2s3 U434 ( .DIN1(RESET), .DIN2(n5260), .Q(WX8544) );
  and2s3 U435 ( .DIN1(RESET), .DIN2(n5265), .Q(WX8542) );
  and2s3 U436 ( .DIN1(RESET), .DIN2(n5270), .Q(WX8540) );
  nor2s3 U437 ( .DIN1(n6537), .DIN2(n6753), .Q(WX854) );
  and2s3 U438 ( .DIN1(RESET), .DIN2(n5275), .Q(WX8538) );
  and2s3 U439 ( .DIN1(RESET), .DIN2(n5280), .Q(WX8536) );
  and2s3 U440 ( .DIN1(RESET), .DIN2(n5285), .Q(WX8534) );
  and2s3 U441 ( .DIN1(RESET), .DIN2(n5290), .Q(WX8532) );
  and2s3 U442 ( .DIN1(RESET), .DIN2(n5295), .Q(WX8530) );
  and2s3 U443 ( .DIN1(RESET), .DIN2(n5155), .Q(WX8528) );
  and2s3 U444 ( .DIN1(RESET), .DIN2(n5159), .Q(WX8526) );
  and2s3 U445 ( .DIN1(RESET), .DIN2(n5163), .Q(WX8524) );
  and2s3 U446 ( .DIN1(RESET), .DIN2(n5167), .Q(WX8522) );
  and2s3 U447 ( .DIN1(RESET), .DIN2(n5171), .Q(WX8520) );
  nor2s3 U448 ( .DIN1(n6512), .DIN2(n6753), .Q(WX852) );
  and2s3 U449 ( .DIN1(RESET), .DIN2(n5175), .Q(WX8518) );
  and2s3 U450 ( .DIN1(RESET), .DIN2(n5179), .Q(WX8516) );
  and2s3 U451 ( .DIN1(RESET), .DIN2(n5183), .Q(WX8514) );
  and2s3 U452 ( .DIN1(RESET), .DIN2(n5187), .Q(WX8512) );
  and2s3 U453 ( .DIN1(RESET), .DIN2(n5191), .Q(WX8510) );
  and2s3 U454 ( .DIN1(RESET), .DIN2(n5195), .Q(WX8508) );
  and2s3 U455 ( .DIN1(RESET), .DIN2(n5199), .Q(WX8506) );
  and2s3 U456 ( .DIN1(RESET), .DIN2(n5203), .Q(WX8504) );
  and2s3 U457 ( .DIN1(RESET), .DIN2(n5207), .Q(WX8502) );
  and2s3 U458 ( .DIN1(RESET), .DIN2(n5211), .Q(WX8500) );
  nor2s3 U459 ( .DIN1(n6502), .DIN2(n6753), .Q(WX850) );
  and2s3 U460 ( .DIN1(RESET), .DIN2(n5215), .Q(WX8498) );
  nor2s3 U461 ( .DIN1(n5219), .DIN2(n6753), .Q(WX8496) );
  nor2s3 U462 ( .DIN1(n5224), .DIN2(n6753), .Q(WX8494) );
  nor2s3 U463 ( .DIN1(n5229), .DIN2(n6753), .Q(WX8492) );
  nor2s3 U464 ( .DIN1(n5234), .DIN2(n6752), .Q(WX8490) );
  nor2s3 U465 ( .DIN1(n5239), .DIN2(n6752), .Q(WX8488) );
  nor2s3 U466 ( .DIN1(n5244), .DIN2(n6752), .Q(WX8486) );
  nor2s3 U467 ( .DIN1(n5249), .DIN2(n6752), .Q(WX8484) );
  nor2s3 U468 ( .DIN1(n5254), .DIN2(n6752), .Q(WX8482) );
  nor2s3 U469 ( .DIN1(n5259), .DIN2(n6752), .Q(WX8480) );
  nor2s3 U470 ( .DIN1(n6541), .DIN2(n6752), .Q(WX848) );
  nor2s3 U471 ( .DIN1(n5264), .DIN2(n6752), .Q(WX8478) );
  nor2s3 U472 ( .DIN1(n5269), .DIN2(n6752), .Q(WX8476) );
  nor2s3 U473 ( .DIN1(n5274), .DIN2(n6752), .Q(WX8474) );
  nor2s3 U474 ( .DIN1(n5279), .DIN2(n6752), .Q(WX8472) );
  nor2s3 U475 ( .DIN1(n5284), .DIN2(n6752), .Q(WX8470) );
  nor2s3 U476 ( .DIN1(n5289), .DIN2(n6751), .Q(WX8468) );
  nor2s3 U477 ( .DIN1(n5294), .DIN2(n6751), .Q(WX8466) );
  nnd4s2 U478 ( .DIN1(n2539), .DIN2(n2540), .DIN3(n2541), .DIN4(n2542), .Q(
        WX8464) );
  nnd2s3 U479 ( .DIN1(n6625), .DIN2(n2313), .Q(n2542) );
  xor2s3 U480 ( .DIN1(n2543), .DIN2(n2544), .Q(n2313) );
  xor2s3 U481 ( .DIN1(n4995), .DIN2(n4996), .Q(n2544) );
  xnr2s3 U482 ( .DIN1(n3205), .DIN2(n4997), .Q(n2543) );
  nnd2s3 U483 ( .DIN1(n2545), .DIN2(n6664), .Q(n2541) );
  nnd2s3 U484 ( .DIN1(n6613), .DIN2(n1889), .Q(n2540) );
  nnd2s3 U485 ( .DIN1(n6582), .DIN2(n1888), .Q(n2539) );
  nnd4s2 U486 ( .DIN1(n2546), .DIN2(n2547), .DIN3(n2548), .DIN4(n2549), .Q(
        WX8462) );
  nnd2s3 U487 ( .DIN1(n2322), .DIN2(n6633), .Q(n2549) );
  xor2s3 U488 ( .DIN1(n2550), .DIN2(n2551), .Q(n2322) );
  xor2s3 U489 ( .DIN1(n4999), .DIN2(n5000), .Q(n2551) );
  xnr2s3 U490 ( .DIN1(n3206), .DIN2(n5001), .Q(n2550) );
  nnd2s3 U491 ( .DIN1(n2552), .DIN2(n6664), .Q(n2548) );
  nnd2s3 U492 ( .DIN1(n6613), .DIN2(n1890), .Q(n2547) );
  nnd2s3 U493 ( .DIN1(n6582), .DIN2(n1887), .Q(n2546) );
  nnd4s2 U494 ( .DIN1(n2553), .DIN2(n2554), .DIN3(n2555), .DIN4(n2556), .Q(
        WX8460) );
  nnd2s3 U495 ( .DIN1(n2328), .DIN2(n6633), .Q(n2556) );
  xor2s3 U496 ( .DIN1(n2557), .DIN2(n2558), .Q(n2328) );
  xor2s3 U497 ( .DIN1(n5003), .DIN2(n5004), .Q(n2558) );
  xnr2s3 U498 ( .DIN1(n3207), .DIN2(n5005), .Q(n2557) );
  nnd2s3 U499 ( .DIN1(n2559), .DIN2(n6664), .Q(n2555) );
  nnd2s3 U500 ( .DIN1(n6613), .DIN2(n1891), .Q(n2554) );
  nnd2s3 U501 ( .DIN1(n6582), .DIN2(n1886), .Q(n2553) );
  nor2s3 U502 ( .DIN1(n6493), .DIN2(n6751), .Q(WX846) );
  nnd4s2 U503 ( .DIN1(n2560), .DIN2(n2561), .DIN3(n2562), .DIN4(n2563), .Q(
        WX8458) );
  nnd2s3 U504 ( .DIN1(n2334), .DIN2(n6633), .Q(n2563) );
  xor2s3 U505 ( .DIN1(n2564), .DIN2(n2565), .Q(n2334) );
  xor2s3 U506 ( .DIN1(n5007), .DIN2(n5008), .Q(n2565) );
  xnr2s3 U507 ( .DIN1(n3208), .DIN2(n5009), .Q(n2564) );
  nnd2s3 U508 ( .DIN1(n2566), .DIN2(n6664), .Q(n2562) );
  nnd2s3 U509 ( .DIN1(n6613), .DIN2(n1892), .Q(n2561) );
  nnd2s3 U510 ( .DIN1(n6582), .DIN2(n1885), .Q(n2560) );
  nnd4s2 U511 ( .DIN1(n2567), .DIN2(n2568), .DIN3(n2569), .DIN4(n2570), .Q(
        WX8456) );
  nnd2s3 U512 ( .DIN1(n2340), .DIN2(n6633), .Q(n2570) );
  xor2s3 U513 ( .DIN1(n2571), .DIN2(n2572), .Q(n2340) );
  xor2s3 U514 ( .DIN1(n5011), .DIN2(n5012), .Q(n2572) );
  xnr2s3 U515 ( .DIN1(n3209), .DIN2(n5013), .Q(n2571) );
  nnd2s3 U516 ( .DIN1(n2573), .DIN2(n6664), .Q(n2569) );
  nnd2s3 U517 ( .DIN1(n6613), .DIN2(n1893), .Q(n2568) );
  nnd2s3 U518 ( .DIN1(n6582), .DIN2(n1884), .Q(n2567) );
  nnd4s2 U519 ( .DIN1(n2574), .DIN2(n2575), .DIN3(n2576), .DIN4(n2577), .Q(
        WX8454) );
  nnd2s3 U520 ( .DIN1(n2346), .DIN2(n6633), .Q(n2577) );
  xor2s3 U521 ( .DIN1(n2578), .DIN2(n2579), .Q(n2346) );
  xor2s3 U522 ( .DIN1(n5015), .DIN2(n5016), .Q(n2579) );
  xnr2s3 U523 ( .DIN1(n3210), .DIN2(n5017), .Q(n2578) );
  nnd2s3 U524 ( .DIN1(n2580), .DIN2(n6664), .Q(n2576) );
  nnd2s3 U525 ( .DIN1(n6613), .DIN2(n1894), .Q(n2575) );
  nnd2s3 U526 ( .DIN1(n6582), .DIN2(n1883), .Q(n2574) );
  nnd4s2 U527 ( .DIN1(n2581), .DIN2(n2582), .DIN3(n2583), .DIN4(n2584), .Q(
        WX8452) );
  nnd2s3 U528 ( .DIN1(n2352), .DIN2(n6633), .Q(n2584) );
  xor2s3 U529 ( .DIN1(n2585), .DIN2(n2586), .Q(n2352) );
  xor2s3 U530 ( .DIN1(n5019), .DIN2(n5020), .Q(n2586) );
  xnr2s3 U531 ( .DIN1(n3211), .DIN2(n5021), .Q(n2585) );
  nnd2s3 U532 ( .DIN1(n2587), .DIN2(n6664), .Q(n2583) );
  nnd2s3 U533 ( .DIN1(n6613), .DIN2(n1895), .Q(n2582) );
  nnd2s3 U534 ( .DIN1(n6582), .DIN2(n1882), .Q(n2581) );
  nnd4s2 U535 ( .DIN1(n2588), .DIN2(n2589), .DIN3(n2590), .DIN4(n2591), .Q(
        WX8450) );
  nnd2s3 U536 ( .DIN1(n2358), .DIN2(n6633), .Q(n2591) );
  xor2s3 U537 ( .DIN1(n2592), .DIN2(n2593), .Q(n2358) );
  xor2s3 U538 ( .DIN1(n5023), .DIN2(n5024), .Q(n2593) );
  xnr2s3 U539 ( .DIN1(n3212), .DIN2(n5025), .Q(n2592) );
  nnd2s3 U540 ( .DIN1(n2594), .DIN2(n6664), .Q(n2590) );
  nnd2s3 U541 ( .DIN1(n6613), .DIN2(n1896), .Q(n2589) );
  nnd2s3 U542 ( .DIN1(n6582), .DIN2(n1881), .Q(n2588) );
  nnd4s2 U543 ( .DIN1(n2595), .DIN2(n2596), .DIN3(n2597), .DIN4(n2598), .Q(
        WX8448) );
  nnd2s3 U544 ( .DIN1(n2364), .DIN2(n6633), .Q(n2598) );
  xor2s3 U545 ( .DIN1(n2599), .DIN2(n2600), .Q(n2364) );
  xor2s3 U546 ( .DIN1(n5027), .DIN2(n5028), .Q(n2600) );
  xnr2s3 U547 ( .DIN1(n3213), .DIN2(n5029), .Q(n2599) );
  nnd2s3 U548 ( .DIN1(n2601), .DIN2(n6664), .Q(n2597) );
  nnd2s3 U549 ( .DIN1(n6613), .DIN2(n1897), .Q(n2596) );
  nnd2s3 U550 ( .DIN1(n6582), .DIN2(n1880), .Q(n2595) );
  nnd4s2 U551 ( .DIN1(n2602), .DIN2(n2603), .DIN3(n2604), .DIN4(n2605), .Q(
        WX8446) );
  nnd2s3 U552 ( .DIN1(n2370), .DIN2(n6633), .Q(n2605) );
  xor2s3 U553 ( .DIN1(n2606), .DIN2(n2607), .Q(n2370) );
  xor2s3 U554 ( .DIN1(n5031), .DIN2(n5032), .Q(n2607) );
  xnr2s3 U555 ( .DIN1(n3214), .DIN2(n5033), .Q(n2606) );
  nnd2s3 U556 ( .DIN1(n2608), .DIN2(n6663), .Q(n2604) );
  nnd2s3 U557 ( .DIN1(n6612), .DIN2(n1898), .Q(n2603) );
  nnd2s3 U558 ( .DIN1(n6581), .DIN2(n1879), .Q(n2602) );
  nnd4s2 U559 ( .DIN1(n2609), .DIN2(n2610), .DIN3(n2611), .DIN4(n2612), .Q(
        WX8444) );
  nnd2s3 U560 ( .DIN1(n2376), .DIN2(n6632), .Q(n2612) );
  xor2s3 U561 ( .DIN1(n2613), .DIN2(n2614), .Q(n2376) );
  xor2s3 U562 ( .DIN1(n5035), .DIN2(n5036), .Q(n2614) );
  xnr2s3 U563 ( .DIN1(n3215), .DIN2(n5037), .Q(n2613) );
  nnd2s3 U564 ( .DIN1(n2615), .DIN2(n6663), .Q(n2611) );
  nnd2s3 U565 ( .DIN1(n6612), .DIN2(n1899), .Q(n2610) );
  nnd2s3 U566 ( .DIN1(n6581), .DIN2(n1878), .Q(n2609) );
  nnd4s2 U567 ( .DIN1(n2616), .DIN2(n2617), .DIN3(n2618), .DIN4(n2619), .Q(
        WX8442) );
  nnd2s3 U568 ( .DIN1(n2382), .DIN2(n6632), .Q(n2619) );
  xor2s3 U569 ( .DIN1(n2620), .DIN2(n2621), .Q(n2382) );
  xor2s3 U570 ( .DIN1(n5039), .DIN2(n5040), .Q(n2621) );
  xnr2s3 U571 ( .DIN1(n3216), .DIN2(n5041), .Q(n2620) );
  nnd2s3 U572 ( .DIN1(n2622), .DIN2(n6663), .Q(n2618) );
  nnd2s3 U573 ( .DIN1(n6612), .DIN2(n1900), .Q(n2617) );
  nnd2s3 U574 ( .DIN1(n6581), .DIN2(n1877), .Q(n2616) );
  nnd4s2 U575 ( .DIN1(n2623), .DIN2(n2624), .DIN3(n2625), .DIN4(n2626), .Q(
        WX8440) );
  nnd2s3 U576 ( .DIN1(n2388), .DIN2(n6632), .Q(n2626) );
  xor2s3 U577 ( .DIN1(n2627), .DIN2(n2628), .Q(n2388) );
  xor2s3 U578 ( .DIN1(n5043), .DIN2(n5044), .Q(n2628) );
  xnr2s3 U579 ( .DIN1(n3217), .DIN2(n5045), .Q(n2627) );
  nnd2s3 U580 ( .DIN1(n2629), .DIN2(n6663), .Q(n2625) );
  nnd2s3 U581 ( .DIN1(n6612), .DIN2(n1901), .Q(n2624) );
  nnd2s3 U582 ( .DIN1(n6581), .DIN2(n1876), .Q(n2623) );
  nor2s3 U583 ( .DIN1(n6487), .DIN2(n6751), .Q(WX844) );
  nnd4s2 U584 ( .DIN1(n2630), .DIN2(n2631), .DIN3(n2632), .DIN4(n2633), .Q(
        WX8438) );
  nnd2s3 U585 ( .DIN1(n2394), .DIN2(n6632), .Q(n2633) );
  xor2s3 U586 ( .DIN1(n2634), .DIN2(n2635), .Q(n2394) );
  xor2s3 U587 ( .DIN1(n5047), .DIN2(n5048), .Q(n2635) );
  xnr2s3 U588 ( .DIN1(n3218), .DIN2(n5049), .Q(n2634) );
  nnd2s3 U589 ( .DIN1(n2636), .DIN2(n6663), .Q(n2632) );
  nnd2s3 U590 ( .DIN1(n6612), .DIN2(n1902), .Q(n2631) );
  nnd2s3 U591 ( .DIN1(n6581), .DIN2(n1875), .Q(n2630) );
  nnd4s2 U592 ( .DIN1(n2637), .DIN2(n2638), .DIN3(n2639), .DIN4(n2640), .Q(
        WX8436) );
  nnd2s3 U593 ( .DIN1(n2400), .DIN2(n6632), .Q(n2640) );
  xor2s3 U594 ( .DIN1(n2641), .DIN2(n2642), .Q(n2400) );
  xor2s3 U595 ( .DIN1(n5051), .DIN2(n5052), .Q(n2642) );
  xnr2s3 U596 ( .DIN1(n3219), .DIN2(n5053), .Q(n2641) );
  nnd2s3 U597 ( .DIN1(n2643), .DIN2(n6663), .Q(n2639) );
  nnd2s3 U598 ( .DIN1(n6612), .DIN2(n1903), .Q(n2638) );
  nnd2s3 U599 ( .DIN1(n6581), .DIN2(n1874), .Q(n2637) );
  nnd4s2 U600 ( .DIN1(n2644), .DIN2(n2645), .DIN3(n2646), .DIN4(n2647), .Q(
        WX8434) );
  nnd2s3 U601 ( .DIN1(n2406), .DIN2(n6632), .Q(n2647) );
  xor2s3 U602 ( .DIN1(n2648), .DIN2(n2649), .Q(n2406) );
  xor2s3 U603 ( .DIN1(n5055), .DIN2(n5056), .Q(n2649) );
  xnr2s3 U604 ( .DIN1(n3220), .DIN2(n5057), .Q(n2648) );
  nnd2s3 U605 ( .DIN1(n2650), .DIN2(n6663), .Q(n2646) );
  nnd2s3 U606 ( .DIN1(n6612), .DIN2(n1904), .Q(n2645) );
  nnd2s3 U607 ( .DIN1(n6581), .DIN2(n1873), .Q(n2644) );
  nnd4s2 U608 ( .DIN1(n2651), .DIN2(n2652), .DIN3(n2653), .DIN4(n2654), .Q(
        WX8432) );
  nnd2s3 U609 ( .DIN1(n2412), .DIN2(n6632), .Q(n2654) );
  xor2s3 U610 ( .DIN1(n2655), .DIN2(n2656), .Q(n2412) );
  xor2s3 U611 ( .DIN1(n5061), .DIN2(n2657), .Q(n2656) );
  xor2s3 U612 ( .DIN1(n5059), .DIN2(n5060), .Q(n2657) );
  xor2s3 U613 ( .DIN1(n6414), .DIN2(n6692), .Q(n2655) );
  nnd2s3 U614 ( .DIN1(n2658), .DIN2(n6663), .Q(n2653) );
  nnd2s3 U615 ( .DIN1(n6612), .DIN2(n1905), .Q(n2652) );
  nnd2s3 U616 ( .DIN1(n6581), .DIN2(n1872), .Q(n2651) );
  nnd4s2 U617 ( .DIN1(n2659), .DIN2(n2660), .DIN3(n2661), .DIN4(n2662), .Q(
        WX8430) );
  nnd2s3 U618 ( .DIN1(n2418), .DIN2(n6632), .Q(n2662) );
  xor2s3 U619 ( .DIN1(n2663), .DIN2(n2664), .Q(n2418) );
  xor2s3 U620 ( .DIN1(n5065), .DIN2(n2665), .Q(n2664) );
  xor2s3 U621 ( .DIN1(n5063), .DIN2(n5064), .Q(n2665) );
  xor2s3 U622 ( .DIN1(n6412), .DIN2(n6687), .Q(n2663) );
  nnd2s3 U623 ( .DIN1(n2666), .DIN2(n6663), .Q(n2661) );
  nnd2s3 U624 ( .DIN1(n6612), .DIN2(n1906), .Q(n2660) );
  nnd2s3 U625 ( .DIN1(n6581), .DIN2(n1871), .Q(n2659) );
  nnd4s2 U626 ( .DIN1(n2667), .DIN2(n2668), .DIN3(n2669), .DIN4(n2670), .Q(
        WX8428) );
  nnd2s3 U627 ( .DIN1(n2424), .DIN2(n6632), .Q(n2670) );
  xor2s3 U628 ( .DIN1(n2671), .DIN2(n2672), .Q(n2424) );
  xor2s3 U629 ( .DIN1(n5069), .DIN2(n2673), .Q(n2672) );
  xor2s3 U630 ( .DIN1(n5067), .DIN2(n5068), .Q(n2673) );
  xor2s3 U631 ( .DIN1(n6410), .DIN2(n6687), .Q(n2671) );
  nnd2s3 U632 ( .DIN1(n2674), .DIN2(n6663), .Q(n2669) );
  nnd2s3 U633 ( .DIN1(n6612), .DIN2(n1907), .Q(n2668) );
  nnd2s3 U634 ( .DIN1(n6581), .DIN2(n1870), .Q(n2667) );
  nnd4s2 U635 ( .DIN1(n2675), .DIN2(n2676), .DIN3(n2677), .DIN4(n2678), .Q(
        WX8426) );
  nnd2s3 U636 ( .DIN1(n2430), .DIN2(n6632), .Q(n2678) );
  xor2s3 U637 ( .DIN1(n2679), .DIN2(n2680), .Q(n2430) );
  xor2s3 U638 ( .DIN1(n5073), .DIN2(n2681), .Q(n2680) );
  xor2s3 U639 ( .DIN1(n5071), .DIN2(n5072), .Q(n2681) );
  xor2s3 U640 ( .DIN1(n6408), .DIN2(n6687), .Q(n2679) );
  nnd2s3 U641 ( .DIN1(n2682), .DIN2(n6663), .Q(n2677) );
  nnd2s3 U642 ( .DIN1(n6612), .DIN2(n1908), .Q(n2676) );
  nnd2s3 U643 ( .DIN1(n6581), .DIN2(n1869), .Q(n2675) );
  nnd4s2 U644 ( .DIN1(n2683), .DIN2(n2684), .DIN3(n2685), .DIN4(n2686), .Q(
        WX8424) );
  nnd2s3 U645 ( .DIN1(n2436), .DIN2(n6632), .Q(n2686) );
  xor2s3 U646 ( .DIN1(n2687), .DIN2(n2688), .Q(n2436) );
  xor2s3 U647 ( .DIN1(n5077), .DIN2(n2689), .Q(n2688) );
  xor2s3 U648 ( .DIN1(n5075), .DIN2(n5076), .Q(n2689) );
  xor2s3 U649 ( .DIN1(n6406), .DIN2(n6687), .Q(n2687) );
  nnd2s3 U650 ( .DIN1(n2690), .DIN2(n6663), .Q(n2685) );
  nnd2s3 U651 ( .DIN1(n6612), .DIN2(n1909), .Q(n2684) );
  nnd2s3 U652 ( .DIN1(n6581), .DIN2(n1868), .Q(n2683) );
  nnd4s2 U653 ( .DIN1(n2691), .DIN2(n2692), .DIN3(n2693), .DIN4(n2694), .Q(
        WX8422) );
  nnd2s3 U654 ( .DIN1(n2442), .DIN2(n6632), .Q(n2694) );
  xor2s3 U655 ( .DIN1(n2695), .DIN2(n2696), .Q(n2442) );
  xor2s3 U656 ( .DIN1(n5081), .DIN2(n2697), .Q(n2696) );
  xor2s3 U657 ( .DIN1(n5079), .DIN2(n5080), .Q(n2697) );
  xor2s3 U658 ( .DIN1(n6404), .DIN2(n6687), .Q(n2695) );
  nnd2s3 U659 ( .DIN1(n2698), .DIN2(n6663), .Q(n2693) );
  nnd2s3 U660 ( .DIN1(n6612), .DIN2(n1910), .Q(n2692) );
  nnd2s3 U661 ( .DIN1(n6581), .DIN2(n1867), .Q(n2691) );
  nnd4s2 U662 ( .DIN1(n2699), .DIN2(n2700), .DIN3(n2701), .DIN4(n2702), .Q(
        WX8420) );
  nnd2s3 U663 ( .DIN1(n2448), .DIN2(n6632), .Q(n2702) );
  xor2s3 U664 ( .DIN1(n2703), .DIN2(n2704), .Q(n2448) );
  xor2s3 U665 ( .DIN1(n5085), .DIN2(n2705), .Q(n2704) );
  xor2s3 U666 ( .DIN1(n5083), .DIN2(n5084), .Q(n2705) );
  xor2s3 U667 ( .DIN1(n6402), .DIN2(n6687), .Q(n2703) );
  nnd2s3 U668 ( .DIN1(n2706), .DIN2(n6662), .Q(n2701) );
  nnd2s3 U669 ( .DIN1(n6611), .DIN2(n1911), .Q(n2700) );
  nnd2s3 U670 ( .DIN1(n6580), .DIN2(n1866), .Q(n2699) );
  nor2s3 U671 ( .DIN1(n6484), .DIN2(n6751), .Q(WX842) );
  nnd4s2 U672 ( .DIN1(n2707), .DIN2(n2708), .DIN3(n2709), .DIN4(n2710), .Q(
        WX8418) );
  nnd2s3 U673 ( .DIN1(n2454), .DIN2(n6631), .Q(n2710) );
  xor2s3 U674 ( .DIN1(n2711), .DIN2(n2712), .Q(n2454) );
  xor2s3 U675 ( .DIN1(n5089), .DIN2(n2713), .Q(n2712) );
  xor2s3 U676 ( .DIN1(n5087), .DIN2(n5088), .Q(n2713) );
  xor2s3 U677 ( .DIN1(n6400), .DIN2(n6687), .Q(n2711) );
  nnd2s3 U678 ( .DIN1(n2714), .DIN2(n6662), .Q(n2709) );
  nnd2s3 U679 ( .DIN1(n6611), .DIN2(n1912), .Q(n2708) );
  nnd2s3 U680 ( .DIN1(n6580), .DIN2(n1865), .Q(n2707) );
  nnd4s2 U681 ( .DIN1(n2715), .DIN2(n2716), .DIN3(n2717), .DIN4(n2718), .Q(
        WX8416) );
  nnd2s3 U682 ( .DIN1(n2460), .DIN2(n6631), .Q(n2718) );
  xor2s3 U683 ( .DIN1(n2719), .DIN2(n2720), .Q(n2460) );
  xor2s3 U684 ( .DIN1(n5093), .DIN2(n2721), .Q(n2720) );
  xor2s3 U685 ( .DIN1(n5091), .DIN2(n5092), .Q(n2721) );
  xor2s3 U686 ( .DIN1(n6398), .DIN2(n6687), .Q(n2719) );
  nnd2s3 U687 ( .DIN1(n2722), .DIN2(n6662), .Q(n2717) );
  nnd2s3 U688 ( .DIN1(n6611), .DIN2(n1913), .Q(n2716) );
  nnd2s3 U689 ( .DIN1(n6580), .DIN2(n1864), .Q(n2715) );
  nnd4s2 U690 ( .DIN1(n2723), .DIN2(n2724), .DIN3(n2725), .DIN4(n2726), .Q(
        WX8414) );
  nnd2s3 U691 ( .DIN1(n2466), .DIN2(n6631), .Q(n2726) );
  xor2s3 U692 ( .DIN1(n2727), .DIN2(n2728), .Q(n2466) );
  xor2s3 U693 ( .DIN1(n5097), .DIN2(n2729), .Q(n2728) );
  xor2s3 U694 ( .DIN1(n5095), .DIN2(n5096), .Q(n2729) );
  xor2s3 U695 ( .DIN1(n6396), .DIN2(n6687), .Q(n2727) );
  nnd2s3 U696 ( .DIN1(n2730), .DIN2(n6662), .Q(n2725) );
  nnd2s3 U697 ( .DIN1(n6611), .DIN2(n1914), .Q(n2724) );
  nnd2s3 U698 ( .DIN1(n6580), .DIN2(n1863), .Q(n2723) );
  nnd4s2 U699 ( .DIN1(n2731), .DIN2(n2732), .DIN3(n2733), .DIN4(n2734), .Q(
        WX8412) );
  nnd2s3 U700 ( .DIN1(n2472), .DIN2(n6631), .Q(n2734) );
  xor2s3 U701 ( .DIN1(n2735), .DIN2(n2736), .Q(n2472) );
  xor2s3 U702 ( .DIN1(n5101), .DIN2(n2737), .Q(n2736) );
  xor2s3 U703 ( .DIN1(n5099), .DIN2(n5100), .Q(n2737) );
  xor2s3 U704 ( .DIN1(n6394), .DIN2(n6687), .Q(n2735) );
  nnd2s3 U705 ( .DIN1(n2738), .DIN2(n6662), .Q(n2733) );
  nnd2s3 U706 ( .DIN1(n6611), .DIN2(n1915), .Q(n2732) );
  nnd2s3 U707 ( .DIN1(n6580), .DIN2(n1862), .Q(n2731) );
  nnd4s2 U708 ( .DIN1(n2739), .DIN2(n2740), .DIN3(n2741), .DIN4(n2742), .Q(
        WX8410) );
  nnd2s3 U709 ( .DIN1(n2478), .DIN2(n6631), .Q(n2742) );
  xor2s3 U710 ( .DIN1(n2743), .DIN2(n2744), .Q(n2478) );
  xor2s3 U711 ( .DIN1(n5105), .DIN2(n2745), .Q(n2744) );
  xor2s3 U712 ( .DIN1(n5103), .DIN2(n5104), .Q(n2745) );
  xor2s3 U713 ( .DIN1(n6392), .DIN2(n6687), .Q(n2743) );
  nnd2s3 U714 ( .DIN1(n2746), .DIN2(n6662), .Q(n2741) );
  nnd2s3 U715 ( .DIN1(n6611), .DIN2(n1916), .Q(n2740) );
  nnd2s3 U716 ( .DIN1(n6580), .DIN2(n1861), .Q(n2739) );
  nnd4s2 U717 ( .DIN1(n2747), .DIN2(n2748), .DIN3(n2749), .DIN4(n2750), .Q(
        WX8408) );
  nnd2s3 U718 ( .DIN1(n2484), .DIN2(n6631), .Q(n2750) );
  xor2s3 U719 ( .DIN1(n2751), .DIN2(n2752), .Q(n2484) );
  xor2s3 U720 ( .DIN1(n5109), .DIN2(n2753), .Q(n2752) );
  xor2s3 U721 ( .DIN1(n5107), .DIN2(n5108), .Q(n2753) );
  xor2s3 U722 ( .DIN1(n6390), .DIN2(n6687), .Q(n2751) );
  nnd2s3 U723 ( .DIN1(n2754), .DIN2(n6662), .Q(n2749) );
  nnd2s3 U724 ( .DIN1(n6611), .DIN2(n1917), .Q(n2748) );
  nnd2s3 U725 ( .DIN1(n6580), .DIN2(n1860), .Q(n2747) );
  nnd4s2 U726 ( .DIN1(n2755), .DIN2(n2756), .DIN3(n2757), .DIN4(n2758), .Q(
        WX8406) );
  nnd2s3 U727 ( .DIN1(n2490), .DIN2(n6631), .Q(n2758) );
  xor2s3 U728 ( .DIN1(n2759), .DIN2(n2760), .Q(n2490) );
  xor2s3 U729 ( .DIN1(n5113), .DIN2(n2761), .Q(n2760) );
  xor2s3 U730 ( .DIN1(n5111), .DIN2(n5112), .Q(n2761) );
  xor2s3 U731 ( .DIN1(n6388), .DIN2(n6688), .Q(n2759) );
  nnd2s3 U732 ( .DIN1(n2762), .DIN2(n6662), .Q(n2757) );
  nnd2s3 U733 ( .DIN1(n6611), .DIN2(n1918), .Q(n2756) );
  nnd2s3 U734 ( .DIN1(n6580), .DIN2(n1859), .Q(n2755) );
  nnd4s2 U735 ( .DIN1(n2763), .DIN2(n2764), .DIN3(n2765), .DIN4(n2766), .Q(
        WX8404) );
  nnd2s3 U736 ( .DIN1(n2496), .DIN2(n6631), .Q(n2766) );
  xor2s3 U737 ( .DIN1(n2767), .DIN2(n2768), .Q(n2496) );
  xor2s3 U738 ( .DIN1(n5117), .DIN2(n2769), .Q(n2768) );
  xor2s3 U739 ( .DIN1(n5115), .DIN2(n5116), .Q(n2769) );
  xor2s3 U740 ( .DIN1(n6386), .DIN2(n6688), .Q(n2767) );
  nnd2s3 U741 ( .DIN1(n2770), .DIN2(n6662), .Q(n2765) );
  nnd2s3 U742 ( .DIN1(n6611), .DIN2(n1919), .Q(n2764) );
  nnd2s3 U743 ( .DIN1(n6580), .DIN2(n1858), .Q(n2763) );
  nnd4s2 U744 ( .DIN1(n2771), .DIN2(n2772), .DIN3(n2773), .DIN4(n2774), .Q(
        WX8402) );
  nnd2s3 U745 ( .DIN1(n2502), .DIN2(n6631), .Q(n2774) );
  xor2s3 U746 ( .DIN1(n2775), .DIN2(n2776), .Q(n2502) );
  xor2s3 U747 ( .DIN1(n5121), .DIN2(n2777), .Q(n2776) );
  xor2s3 U748 ( .DIN1(n5119), .DIN2(n5120), .Q(n2777) );
  xor2s3 U749 ( .DIN1(n6384), .DIN2(n6688), .Q(n2775) );
  nnd2s3 U750 ( .DIN1(n2778), .DIN2(n6662), .Q(n2773) );
  nnd2s3 U751 ( .DIN1(n6611), .DIN2(n1920), .Q(n2772) );
  nnd2s3 U752 ( .DIN1(n6580), .DIN2(n1857), .Q(n2771) );
  nor2s3 U753 ( .DIN1(n6547), .DIN2(n6751), .Q(WX840) );
  nor2s3 U754 ( .DIN1(n6475), .DIN2(n6751), .Q(WX838) );
  nor2s3 U755 ( .DIN1(n6531), .DIN2(n6751), .Q(WX836) );
  nor2s3 U756 ( .DIN1(n6464), .DIN2(n6751), .Q(WX834) );
  nor2s3 U757 ( .DIN1(n6528), .DIN2(n6751), .Q(WX832) );
  nor2s3 U758 ( .DIN1(n6805), .DIN2(n1920), .Q(WX8304) );
  nor2s3 U759 ( .DIN1(n5124), .DIN2(n6751), .Q(WX8302) );
  nor2s3 U760 ( .DIN1(n5125), .DIN2(n6751), .Q(WX8300) );
  nor2s3 U761 ( .DIN1(n6562), .DIN2(n6750), .Q(WX830) );
  nor2s3 U762 ( .DIN1(n5126), .DIN2(n6750), .Q(WX8298) );
  nor2s3 U763 ( .DIN1(n5127), .DIN2(n6750), .Q(WX8296) );
  nor2s3 U764 ( .DIN1(n5128), .DIN2(n6750), .Q(WX8294) );
  nor2s3 U765 ( .DIN1(n5129), .DIN2(n6750), .Q(WX8292) );
  nor2s3 U766 ( .DIN1(n5130), .DIN2(n6750), .Q(WX8290) );
  nor2s3 U767 ( .DIN1(n5131), .DIN2(n6750), .Q(WX8288) );
  nor2s3 U768 ( .DIN1(n5132), .DIN2(n6750), .Q(WX8286) );
  nor2s3 U769 ( .DIN1(n5133), .DIN2(n6750), .Q(WX8284) );
  nor2s3 U770 ( .DIN1(n5134), .DIN2(n6750), .Q(WX8282) );
  nor2s3 U771 ( .DIN1(n5135), .DIN2(n6750), .Q(WX8280) );
  nor2s3 U772 ( .DIN1(n6470), .DIN2(n6749), .Q(WX828) );
  nor2s3 U773 ( .DIN1(n5136), .DIN2(n6749), .Q(WX8278) );
  nor2s3 U774 ( .DIN1(n5137), .DIN2(n6749), .Q(WX8276) );
  nor2s3 U775 ( .DIN1(n5138), .DIN2(n6749), .Q(WX8274) );
  nor2s3 U776 ( .DIN1(n5139), .DIN2(n6749), .Q(WX8272) );
  nor2s3 U777 ( .DIN1(n5140), .DIN2(n6749), .Q(WX8270) );
  nor2s3 U778 ( .DIN1(n5141), .DIN2(n6749), .Q(WX8268) );
  nor2s3 U779 ( .DIN1(n5142), .DIN2(n6749), .Q(WX8266) );
  nor2s3 U780 ( .DIN1(n5143), .DIN2(n6749), .Q(WX8264) );
  nor2s3 U781 ( .DIN1(n5144), .DIN2(n6749), .Q(WX8262) );
  nor2s3 U782 ( .DIN1(n5145), .DIN2(n6749), .Q(WX8260) );
  nor2s3 U783 ( .DIN1(n6473), .DIN2(n6749), .Q(WX826) );
  nor2s3 U784 ( .DIN1(n5146), .DIN2(n6748), .Q(WX8258) );
  nor2s3 U785 ( .DIN1(n5147), .DIN2(n6748), .Q(WX8256) );
  nor2s3 U786 ( .DIN1(n5148), .DIN2(n6748), .Q(WX8254) );
  nor2s3 U787 ( .DIN1(n5149), .DIN2(n6748), .Q(WX8252) );
  nor2s3 U788 ( .DIN1(n5150), .DIN2(n6748), .Q(WX8250) );
  nor2s3 U789 ( .DIN1(n5151), .DIN2(n6748), .Q(WX8248) );
  nor2s3 U790 ( .DIN1(n5152), .DIN2(n6748), .Q(WX8246) );
  nor2s3 U791 ( .DIN1(n5153), .DIN2(n6748), .Q(WX8244) );
  nor2s3 U792 ( .DIN1(n5154), .DIN2(n6748), .Q(WX8242) );
  nor2s3 U793 ( .DIN1(n6461), .DIN2(n6748), .Q(WX824) );
  nor2s3 U794 ( .DIN1(n6443), .DIN2(n6748), .Q(WX822) );
  nor2s3 U795 ( .DIN1(n6467), .DIN2(n6748), .Q(WX820) );
  nor2s3 U796 ( .DIN1(n6455), .DIN2(n6747), .Q(WX818) );
  nor2s3 U797 ( .DIN1(n6505), .DIN2(n6747), .Q(WX816) );
  nor2s3 U798 ( .DIN1(n6452), .DIN2(n6747), .Q(WX814) );
  nor2s3 U799 ( .DIN1(n6446), .DIN2(n6747), .Q(WX812) );
  nor2s3 U800 ( .DIN1(n6458), .DIN2(n6747), .Q(WX810) );
  nor2s3 U801 ( .DIN1(n6449), .DIN2(n6747), .Q(WX808) );
  nor2s3 U802 ( .DIN1(n6524), .DIN2(n6747), .Q(WX806) );
  nor2s3 U803 ( .DIN1(n6440), .DIN2(n6747), .Q(WX804) );
  nor2s3 U804 ( .DIN1(n6508), .DIN2(n6747), .Q(WX802) );
  nor2s3 U805 ( .DIN1(n6497), .DIN2(n6747), .Q(WX800) );
  nor2s3 U806 ( .DIN1(n6489), .DIN2(n6747), .Q(WX798) );
  nor2s3 U807 ( .DIN1(n6479), .DIN2(n6747), .Q(WX796) );
  nor2s3 U808 ( .DIN1(n6520), .DIN2(n6746), .Q(WX794) );
  nor2s3 U809 ( .DIN1(n6519), .DIN2(n6746), .Q(WX792) );
  nor2s3 U810 ( .DIN1(n6514), .DIN2(n6746), .Q(WX790) );
  nor2s3 U811 ( .DIN1(n6513), .DIN2(n6746), .Q(WX788) );
  nor2s3 U812 ( .DIN1(n6503), .DIN2(n6746), .Q(WX786) );
  nor2s3 U813 ( .DIN1(n6498), .DIN2(n6746), .Q(WX784) );
  nor2s3 U814 ( .DIN1(n6494), .DIN2(n6746), .Q(WX782) );
  nor2s3 U815 ( .DIN1(n6488), .DIN2(n6746), .Q(WX780) );
  nor2s3 U816 ( .DIN1(n6802), .DIN2(n2779), .Q(WX7791) );
  xor2s3 U817 ( .DIN1(n5293), .DIN2(n5473), .Q(n2779) );
  nor2s3 U818 ( .DIN1(n6802), .DIN2(n2780), .Q(WX7789) );
  xor2s3 U819 ( .DIN1(n5288), .DIN2(n5468), .Q(n2780) );
  nor2s3 U820 ( .DIN1(n6802), .DIN2(n2781), .Q(WX7787) );
  xor2s3 U821 ( .DIN1(n5283), .DIN2(n5463), .Q(n2781) );
  nor2s3 U822 ( .DIN1(n6802), .DIN2(n2782), .Q(WX7785) );
  xor2s3 U823 ( .DIN1(n5278), .DIN2(n5458), .Q(n2782) );
  nor2s3 U824 ( .DIN1(n6802), .DIN2(n2783), .Q(WX7783) );
  xor2s3 U825 ( .DIN1(n5273), .DIN2(n5453), .Q(n2783) );
  nor2s3 U826 ( .DIN1(n6802), .DIN2(n2784), .Q(WX7781) );
  xor2s3 U827 ( .DIN1(n5268), .DIN2(n5448), .Q(n2784) );
  nor2s3 U828 ( .DIN1(n6485), .DIN2(n6746), .Q(WX778) );
  nor2s3 U829 ( .DIN1(n6802), .DIN2(n2785), .Q(WX7779) );
  xor2s3 U830 ( .DIN1(n5263), .DIN2(n5443), .Q(n2785) );
  nor2s3 U831 ( .DIN1(n6802), .DIN2(n2786), .Q(WX7777) );
  xor2s3 U832 ( .DIN1(n5258), .DIN2(n5438), .Q(n2786) );
  nor2s3 U833 ( .DIN1(n6801), .DIN2(n2787), .Q(WX7775) );
  xor2s3 U834 ( .DIN1(n5253), .DIN2(n5433), .Q(n2787) );
  nor2s3 U835 ( .DIN1(n6801), .DIN2(n2788), .Q(WX7773) );
  xor2s3 U836 ( .DIN1(n5248), .DIN2(n5428), .Q(n2788) );
  nor2s3 U837 ( .DIN1(n6801), .DIN2(n2789), .Q(WX7771) );
  xor2s3 U838 ( .DIN1(n5243), .DIN2(n5423), .Q(n2789) );
  nor2s3 U839 ( .DIN1(n6801), .DIN2(n2790), .Q(WX7769) );
  xor2s3 U840 ( .DIN1(n5238), .DIN2(n5418), .Q(n2790) );
  nor2s3 U841 ( .DIN1(n6801), .DIN2(n2791), .Q(WX7767) );
  xor2s3 U842 ( .DIN1(n5233), .DIN2(n5413), .Q(n2791) );
  nor2s3 U843 ( .DIN1(n6801), .DIN2(n2792), .Q(WX7765) );
  xor2s3 U844 ( .DIN1(n5228), .DIN2(n5408), .Q(n2792) );
  nor2s3 U845 ( .DIN1(n6801), .DIN2(n2793), .Q(WX7763) );
  xor2s3 U846 ( .DIN1(n5223), .DIN2(n5403), .Q(n2793) );
  nor2s3 U847 ( .DIN1(n2794), .DIN2(n6746), .Q(WX7761) );
  xnr2s3 U848 ( .DIN1(n5398), .DIN2(n2795), .Q(n2794) );
  xor2s3 U849 ( .DIN1(n5218), .DIN2(n5298), .Q(n2795) );
  nor2s3 U850 ( .DIN1(n6480), .DIN2(n6746), .Q(WX776) );
  nor2s3 U851 ( .DIN1(n6801), .DIN2(n2796), .Q(WX7759) );
  xor2s3 U852 ( .DIN1(n5214), .DIN2(n3252), .Q(n2796) );
  nor2s3 U853 ( .DIN1(n6801), .DIN2(n2797), .Q(WX7757) );
  xor2s3 U854 ( .DIN1(n5210), .DIN2(n3251), .Q(n2797) );
  nor2s3 U855 ( .DIN1(n6801), .DIN2(n2798), .Q(WX7755) );
  xor2s3 U856 ( .DIN1(n5206), .DIN2(n3250), .Q(n2798) );
  nor2s3 U857 ( .DIN1(n6801), .DIN2(n2799), .Q(WX7753) );
  xor2s3 U858 ( .DIN1(n5202), .DIN2(n3249), .Q(n2799) );
  nor2s3 U859 ( .DIN1(n2800), .DIN2(n6746), .Q(WX7751) );
  xnr2s3 U860 ( .DIN1(n3248), .DIN2(n2801), .Q(n2800) );
  xor2s3 U861 ( .DIN1(n5198), .DIN2(n5298), .Q(n2801) );
  nor2s3 U862 ( .DIN1(n6801), .DIN2(n2802), .Q(WX7749) );
  xor2s3 U863 ( .DIN1(n5194), .DIN2(n3247), .Q(n2802) );
  nor2s3 U864 ( .DIN1(n6801), .DIN2(n2803), .Q(WX7747) );
  xor2s3 U865 ( .DIN1(n5190), .DIN2(n3246), .Q(n2803) );
  nor2s3 U866 ( .DIN1(n6800), .DIN2(n2804), .Q(WX7745) );
  xor2s3 U867 ( .DIN1(n5186), .DIN2(n3245), .Q(n2804) );
  nor2s3 U868 ( .DIN1(n6800), .DIN2(n2805), .Q(WX7743) );
  xor2s3 U869 ( .DIN1(n5182), .DIN2(n3244), .Q(n2805) );
  nor2s3 U870 ( .DIN1(n6795), .DIN2(n2806), .Q(WX7741) );
  xor2s3 U871 ( .DIN1(n5178), .DIN2(n3243), .Q(n2806) );
  nor2s3 U872 ( .DIN1(n6476), .DIN2(n6745), .Q(WX774) );
  nor2s3 U873 ( .DIN1(n6800), .DIN2(n2807), .Q(WX7739) );
  xor2s3 U874 ( .DIN1(n5174), .DIN2(n3242), .Q(n2807) );
  nor2s3 U875 ( .DIN1(n2808), .DIN2(n6745), .Q(WX7737) );
  xnr2s3 U876 ( .DIN1(n3241), .DIN2(n2809), .Q(n2808) );
  xor2s3 U877 ( .DIN1(n5170), .DIN2(n5298), .Q(n2809) );
  nor2s3 U878 ( .DIN1(n6800), .DIN2(n2810), .Q(WX7735) );
  xor2s3 U879 ( .DIN1(n5166), .DIN2(n3240), .Q(n2810) );
  nor2s3 U880 ( .DIN1(n6800), .DIN2(n2811), .Q(WX7733) );
  xor2s3 U881 ( .DIN1(n5162), .DIN2(n3239), .Q(n2811) );
  nor2s3 U882 ( .DIN1(n6800), .DIN2(n2812), .Q(WX7731) );
  xor2s3 U883 ( .DIN1(n5158), .DIN2(n3238), .Q(n2812) );
  nor2s3 U884 ( .DIN1(n6800), .DIN2(n2813), .Q(WX7729) );
  xor2s3 U885 ( .DIN1(n5298), .DIN2(n3237), .Q(n2813) );
  nor2s3 U886 ( .DIN1(n6532), .DIN2(n6745), .Q(WX772) );
  nor2s3 U887 ( .DIN1(n6553), .DIN2(n6745), .Q(WX770) );
  nor2s3 U888 ( .DIN1(n6529), .DIN2(n6745), .Q(WX768) );
  nor2s3 U889 ( .DIN1(n6435), .DIN2(n6745), .Q(WX766) );
  nor2s3 U890 ( .DIN1(n6551), .DIN2(n6745), .Q(WX764) );
  nor2s3 U891 ( .DIN1(n6550), .DIN2(n6745), .Q(WX762) );
  nor2s3 U892 ( .DIN1(n6554), .DIN2(n6745), .Q(WX760) );
  nor2s3 U893 ( .DIN1(n6560), .DIN2(n6750), .Q(WX758) );
  nor2s3 U894 ( .DIN1(n6552), .DIN2(n6723), .Q(WX756) );
  nor2s3 U895 ( .DIN1(n6556), .DIN2(n6722), .Q(WX754) );
  nor2s3 U896 ( .DIN1(n6507), .DIN2(n6722), .Q(WX752) );
  nor2s3 U897 ( .DIN1(n6557), .DIN2(n6722), .Q(WX750) );
  nor2s3 U898 ( .DIN1(n6559), .DIN2(n6722), .Q(WX748) );
  nor2s3 U899 ( .DIN1(n6555), .DIN2(n6722), .Q(WX746) );
  nor2s3 U900 ( .DIN1(n6558), .DIN2(n6722), .Q(WX744) );
  nor2s3 U901 ( .DIN1(n6526), .DIN2(n6722), .Q(WX742) );
  nor2s3 U902 ( .DIN1(n6561), .DIN2(n6722), .Q(WX740) );
  nor2s3 U903 ( .DIN1(n6509), .DIN2(n6722), .Q(WX738) );
  nor2s3 U904 ( .DIN1(n5333), .DIN2(n6722), .Q(WX7363) );
  nor2s3 U905 ( .DIN1(n5337), .DIN2(n6722), .Q(WX7361) );
  nor2s3 U906 ( .DIN1(n6542), .DIN2(n6722), .Q(WX736) );
  nor2s3 U907 ( .DIN1(n5341), .DIN2(n6721), .Q(WX7359) );
  nor2s3 U908 ( .DIN1(n5345), .DIN2(n6721), .Q(WX7357) );
  nor2s3 U909 ( .DIN1(n5349), .DIN2(n6721), .Q(WX7355) );
  nor2s3 U910 ( .DIN1(n5353), .DIN2(n6721), .Q(WX7353) );
  nor2s3 U911 ( .DIN1(n5357), .DIN2(n6721), .Q(WX7351) );
  nor2s3 U912 ( .DIN1(n5361), .DIN2(n6721), .Q(WX7349) );
  nor2s3 U913 ( .DIN1(n5365), .DIN2(n6721), .Q(WX7347) );
  nor2s3 U914 ( .DIN1(n5369), .DIN2(n6721), .Q(WX7345) );
  nor2s3 U915 ( .DIN1(n5373), .DIN2(n6721), .Q(WX7343) );
  nor2s3 U916 ( .DIN1(n5377), .DIN2(n6721), .Q(WX7341) );
  nor2s3 U917 ( .DIN1(n6490), .DIN2(n6721), .Q(WX734) );
  nor2s3 U918 ( .DIN1(n5381), .DIN2(n6721), .Q(WX7339) );
  nor2s3 U919 ( .DIN1(n5385), .DIN2(n6720), .Q(WX7337) );
  nor2s3 U920 ( .DIN1(n5389), .DIN2(n6720), .Q(WX7335) );
  nor2s3 U921 ( .DIN1(n5393), .DIN2(n6720), .Q(WX7333) );
  nor2s3 U922 ( .DIN1(n5397), .DIN2(n6720), .Q(WX7331) );
  nor2s3 U923 ( .DIN1(n5402), .DIN2(n6720), .Q(WX7329) );
  nor2s3 U924 ( .DIN1(n5407), .DIN2(n6720), .Q(WX7327) );
  nor2s3 U925 ( .DIN1(n5412), .DIN2(n6720), .Q(WX7325) );
  nor2s3 U926 ( .DIN1(n5417), .DIN2(n6720), .Q(WX7323) );
  nor2s3 U927 ( .DIN1(n5422), .DIN2(n6720), .Q(WX7321) );
  nor2s3 U928 ( .DIN1(n6548), .DIN2(n6720), .Q(WX732) );
  nor2s3 U929 ( .DIN1(n5427), .DIN2(n6720), .Q(WX7319) );
  nor2s3 U930 ( .DIN1(n5432), .DIN2(n6720), .Q(WX7317) );
  nor2s3 U931 ( .DIN1(n5437), .DIN2(n6719), .Q(WX7315) );
  nor2s3 U932 ( .DIN1(n5442), .DIN2(n6719), .Q(WX7313) );
  nor2s3 U933 ( .DIN1(n5447), .DIN2(n6719), .Q(WX7311) );
  nor2s3 U934 ( .DIN1(n5452), .DIN2(n6719), .Q(WX7309) );
  nor2s3 U935 ( .DIN1(n5457), .DIN2(n6719), .Q(WX7307) );
  nor2s3 U936 ( .DIN1(n5462), .DIN2(n6719), .Q(WX7305) );
  nor2s3 U937 ( .DIN1(n5467), .DIN2(n6719), .Q(WX7303) );
  nor2s3 U938 ( .DIN1(n5472), .DIN2(n6719), .Q(WX7301) );
  nor2s3 U939 ( .DIN1(n6521), .DIN2(n6719), .Q(WX730) );
  nor2s3 U940 ( .DIN1(n5332), .DIN2(n6719), .Q(WX7299) );
  nor2s3 U941 ( .DIN1(n5336), .DIN2(n6719), .Q(WX7297) );
  nor2s3 U942 ( .DIN1(n5340), .DIN2(n6719), .Q(WX7295) );
  nor2s3 U943 ( .DIN1(n5344), .DIN2(n6718), .Q(WX7293) );
  nor2s3 U944 ( .DIN1(n5348), .DIN2(n6718), .Q(WX7291) );
  nor2s3 U945 ( .DIN1(n5352), .DIN2(n6718), .Q(WX7289) );
  nor2s3 U946 ( .DIN1(n5356), .DIN2(n6718), .Q(WX7287) );
  nor2s3 U947 ( .DIN1(n5360), .DIN2(n6718), .Q(WX7285) );
  nor2s3 U948 ( .DIN1(n5364), .DIN2(n6718), .Q(WX7283) );
  nor2s3 U949 ( .DIN1(n5368), .DIN2(n6718), .Q(WX7281) );
  nor2s3 U950 ( .DIN1(n6536), .DIN2(n6718), .Q(WX728) );
  nor2s3 U951 ( .DIN1(n5372), .DIN2(n6718), .Q(WX7279) );
  nor2s3 U952 ( .DIN1(n5376), .DIN2(n6718), .Q(WX7277) );
  nor2s3 U953 ( .DIN1(n5380), .DIN2(n6718), .Q(WX7275) );
  nor2s3 U954 ( .DIN1(n5384), .DIN2(n6718), .Q(WX7273) );
  nor2s3 U955 ( .DIN1(n5388), .DIN2(n6717), .Q(WX7271) );
  nor2s3 U956 ( .DIN1(n5392), .DIN2(n6717), .Q(WX7269) );
  and2s3 U957 ( .DIN1(RESET), .DIN2(n5396), .Q(WX7267) );
  and2s3 U958 ( .DIN1(RESET), .DIN2(n5401), .Q(WX7265) );
  and2s3 U959 ( .DIN1(RESET), .DIN2(n5406), .Q(WX7263) );
  and2s3 U960 ( .DIN1(RESET), .DIN2(n5411), .Q(WX7261) );
  nor2s3 U961 ( .DIN1(n6515), .DIN2(n6717), .Q(WX726) );
  and2s3 U962 ( .DIN1(RESET), .DIN2(n5416), .Q(WX7259) );
  and2s3 U963 ( .DIN1(RESET), .DIN2(n5421), .Q(WX7257) );
  and2s3 U964 ( .DIN1(RESET), .DIN2(n5426), .Q(WX7255) );
  and2s3 U965 ( .DIN1(RESET), .DIN2(n5431), .Q(WX7253) );
  and2s3 U966 ( .DIN1(RESET), .DIN2(n5436), .Q(WX7251) );
  and2s3 U967 ( .DIN1(RESET), .DIN2(n5441), .Q(WX7249) );
  and2s3 U968 ( .DIN1(RESET), .DIN2(n5446), .Q(WX7247) );
  and2s3 U969 ( .DIN1(RESET), .DIN2(n5451), .Q(WX7245) );
  and2s3 U970 ( .DIN1(RESET), .DIN2(n5456), .Q(WX7243) );
  and2s3 U971 ( .DIN1(RESET), .DIN2(n5461), .Q(WX7241) );
  nor2s3 U972 ( .DIN1(n6538), .DIN2(n6717), .Q(WX724) );
  and2s3 U973 ( .DIN1(RESET), .DIN2(n5466), .Q(WX7239) );
  and2s3 U974 ( .DIN1(RESET), .DIN2(n5471), .Q(WX7237) );
  and2s3 U975 ( .DIN1(RESET), .DIN2(n5331), .Q(WX7235) );
  and2s3 U976 ( .DIN1(RESET), .DIN2(n5335), .Q(WX7233) );
  and2s3 U977 ( .DIN1(RESET), .DIN2(n5339), .Q(WX7231) );
  and2s3 U978 ( .DIN1(RESET), .DIN2(n5343), .Q(WX7229) );
  and2s3 U979 ( .DIN1(RESET), .DIN2(n5347), .Q(WX7227) );
  and2s3 U980 ( .DIN1(RESET), .DIN2(n5351), .Q(WX7225) );
  and2s3 U981 ( .DIN1(RESET), .DIN2(n5355), .Q(WX7223) );
  and2s3 U982 ( .DIN1(RESET), .DIN2(n5359), .Q(WX7221) );
  nor2s3 U983 ( .DIN1(n6540), .DIN2(n6717), .Q(WX722) );
  and2s3 U984 ( .DIN1(RESET), .DIN2(n5363), .Q(WX7219) );
  and2s3 U985 ( .DIN1(RESET), .DIN2(n5367), .Q(WX7217) );
  and2s3 U986 ( .DIN1(RESET), .DIN2(n5371), .Q(WX7215) );
  and2s3 U987 ( .DIN1(RESET), .DIN2(n5375), .Q(WX7213) );
  and2s3 U988 ( .DIN1(RESET), .DIN2(n5379), .Q(WX7211) );
  and2s3 U989 ( .DIN1(RESET), .DIN2(n5383), .Q(WX7209) );
  and2s3 U990 ( .DIN1(RESET), .DIN2(n5387), .Q(WX7207) );
  and2s3 U991 ( .DIN1(RESET), .DIN2(n5391), .Q(WX7205) );
  nor2s3 U992 ( .DIN1(n5395), .DIN2(n6717), .Q(WX7203) );
  nor2s3 U993 ( .DIN1(n5400), .DIN2(n6717), .Q(WX7201) );
  nor2s3 U994 ( .DIN1(n6499), .DIN2(n6717), .Q(WX720) );
  nor2s3 U995 ( .DIN1(n5405), .DIN2(n6717), .Q(WX7199) );
  nor2s3 U996 ( .DIN1(n5410), .DIN2(n6717), .Q(WX7197) );
  nor2s3 U997 ( .DIN1(n5415), .DIN2(n6717), .Q(WX7195) );
  nor2s3 U998 ( .DIN1(n5420), .DIN2(n6716), .Q(WX7193) );
  nor2s3 U999 ( .DIN1(n5425), .DIN2(n6716), .Q(WX7191) );
  nor2s3 U1000 ( .DIN1(n5430), .DIN2(n6716), .Q(WX7189) );
  nor2s3 U1001 ( .DIN1(n5435), .DIN2(n6716), .Q(WX7187) );
  nor2s3 U1002 ( .DIN1(n5440), .DIN2(n6716), .Q(WX7185) );
  nor2s3 U1003 ( .DIN1(n5445), .DIN2(n6716), .Q(WX7183) );
  nor2s3 U1004 ( .DIN1(n5450), .DIN2(n6716), .Q(WX7181) );
  nor2s3 U1005 ( .DIN1(n6543), .DIN2(n6716), .Q(WX718) );
  nor2s3 U1006 ( .DIN1(n5455), .DIN2(n6716), .Q(WX7179) );
  nor2s3 U1007 ( .DIN1(n5460), .DIN2(n6716), .Q(WX7177) );
  nor2s3 U1008 ( .DIN1(n5465), .DIN2(n6716), .Q(WX7175) );
  nor2s3 U1009 ( .DIN1(n5470), .DIN2(n6716), .Q(WX7173) );
  nnd4s2 U1010 ( .DIN1(n2814), .DIN2(n2815), .DIN3(n2816), .DIN4(n2817), .Q(
        WX7171) );
  nnd2s3 U1011 ( .DIN1(n2545), .DIN2(n6631), .Q(n2817) );
  xor2s3 U1012 ( .DIN1(n2818), .DIN2(n2819), .Q(n2545) );
  xor2s3 U1013 ( .DIN1(n5155), .DIN2(n5156), .Q(n2819) );
  xnr2s3 U1014 ( .DIN1(n3221), .DIN2(n5157), .Q(n2818) );
  nnd2s3 U1015 ( .DIN1(n2820), .DIN2(n6662), .Q(n2816) );
  nnd2s3 U1016 ( .DIN1(n6611), .DIN2(n1953), .Q(n2815) );
  nnd2s3 U1017 ( .DIN1(n6580), .DIN2(n1952), .Q(n2814) );
  nnd4s2 U1018 ( .DIN1(n2821), .DIN2(n2822), .DIN3(n2823), .DIN4(n2824), .Q(
        WX7169) );
  nnd2s3 U1019 ( .DIN1(n2552), .DIN2(n6631), .Q(n2824) );
  xor2s3 U1020 ( .DIN1(n2825), .DIN2(n2826), .Q(n2552) );
  xor2s3 U1021 ( .DIN1(n5159), .DIN2(n5160), .Q(n2826) );
  xnr2s3 U1022 ( .DIN1(n3222), .DIN2(n5161), .Q(n2825) );
  nnd2s3 U1023 ( .DIN1(n2827), .DIN2(n6662), .Q(n2823) );
  nnd2s3 U1024 ( .DIN1(n6611), .DIN2(n1954), .Q(n2822) );
  nnd2s3 U1025 ( .DIN1(n6580), .DIN2(n1951), .Q(n2821) );
  nnd4s2 U1026 ( .DIN1(n2828), .DIN2(n2829), .DIN3(n2830), .DIN4(n2831), .Q(
        WX7167) );
  nnd2s3 U1027 ( .DIN1(n2559), .DIN2(n6631), .Q(n2831) );
  xor2s3 U1028 ( .DIN1(n2832), .DIN2(n2833), .Q(n2559) );
  xor2s3 U1029 ( .DIN1(n5163), .DIN2(n5164), .Q(n2833) );
  xnr2s3 U1030 ( .DIN1(n3223), .DIN2(n5165), .Q(n2832) );
  nnd2s3 U1031 ( .DIN1(n2834), .DIN2(n6662), .Q(n2830) );
  nnd2s3 U1032 ( .DIN1(n6611), .DIN2(n1955), .Q(n2829) );
  nnd2s3 U1033 ( .DIN1(n6580), .DIN2(n1950), .Q(n2828) );
  nnd4s2 U1034 ( .DIN1(n2835), .DIN2(n2836), .DIN3(n2837), .DIN4(n2838), .Q(
        WX7165) );
  nnd2s3 U1035 ( .DIN1(n2566), .DIN2(n6631), .Q(n2838) );
  xor2s3 U1036 ( .DIN1(n2839), .DIN2(n2840), .Q(n2566) );
  xor2s3 U1037 ( .DIN1(n5167), .DIN2(n5168), .Q(n2840) );
  xnr2s3 U1038 ( .DIN1(n3224), .DIN2(n5169), .Q(n2839) );
  nnd2s3 U1039 ( .DIN1(n2841), .DIN2(n6661), .Q(n2837) );
  nnd2s3 U1040 ( .DIN1(n6610), .DIN2(n1956), .Q(n2836) );
  nnd2s3 U1041 ( .DIN1(n6579), .DIN2(n1949), .Q(n2835) );
  nnd4s2 U1042 ( .DIN1(n2842), .DIN2(n2843), .DIN3(n2844), .DIN4(n2845), .Q(
        WX7163) );
  nnd2s3 U1043 ( .DIN1(n2573), .DIN2(n6630), .Q(n2845) );
  xor2s3 U1044 ( .DIN1(n2846), .DIN2(n2847), .Q(n2573) );
  xor2s3 U1045 ( .DIN1(n5171), .DIN2(n5172), .Q(n2847) );
  xnr2s3 U1046 ( .DIN1(n3225), .DIN2(n5173), .Q(n2846) );
  nnd2s3 U1047 ( .DIN1(n2848), .DIN2(n6661), .Q(n2844) );
  nnd2s3 U1048 ( .DIN1(n6610), .DIN2(n1957), .Q(n2843) );
  nnd2s3 U1049 ( .DIN1(n6579), .DIN2(n1948), .Q(n2842) );
  nnd4s2 U1050 ( .DIN1(n2849), .DIN2(n2850), .DIN3(n2851), .DIN4(n2852), .Q(
        WX7161) );
  nnd2s3 U1051 ( .DIN1(n2580), .DIN2(n6630), .Q(n2852) );
  xor2s3 U1052 ( .DIN1(n2853), .DIN2(n2854), .Q(n2580) );
  xor2s3 U1053 ( .DIN1(n5175), .DIN2(n5176), .Q(n2854) );
  xnr2s3 U1054 ( .DIN1(n3226), .DIN2(n5177), .Q(n2853) );
  nnd2s3 U1055 ( .DIN1(n2855), .DIN2(n6661), .Q(n2851) );
  nnd2s3 U1056 ( .DIN1(n6610), .DIN2(n1958), .Q(n2850) );
  nnd2s3 U1057 ( .DIN1(n6579), .DIN2(n1947), .Q(n2849) );
  nor2s3 U1058 ( .DIN1(n6545), .DIN2(n6715), .Q(WX716) );
  nnd4s2 U1059 ( .DIN1(n2856), .DIN2(n2857), .DIN3(n2858), .DIN4(n2859), .Q(
        WX7159) );
  nnd2s3 U1060 ( .DIN1(n2587), .DIN2(n6630), .Q(n2859) );
  xor2s3 U1061 ( .DIN1(n2860), .DIN2(n2861), .Q(n2587) );
  xor2s3 U1062 ( .DIN1(n5179), .DIN2(n5180), .Q(n2861) );
  xnr2s3 U1063 ( .DIN1(n3227), .DIN2(n5181), .Q(n2860) );
  nnd2s3 U1064 ( .DIN1(n2862), .DIN2(n6661), .Q(n2858) );
  nnd2s3 U1065 ( .DIN1(n6610), .DIN2(n1959), .Q(n2857) );
  nnd2s3 U1066 ( .DIN1(n6579), .DIN2(n1946), .Q(n2856) );
  nnd4s2 U1067 ( .DIN1(n2863), .DIN2(n2864), .DIN3(n2865), .DIN4(n2866), .Q(
        WX7157) );
  nnd2s3 U1068 ( .DIN1(n2594), .DIN2(n6630), .Q(n2866) );
  xor2s3 U1069 ( .DIN1(n2867), .DIN2(n2868), .Q(n2594) );
  xor2s3 U1070 ( .DIN1(n5183), .DIN2(n5184), .Q(n2868) );
  xnr2s3 U1071 ( .DIN1(n3228), .DIN2(n5185), .Q(n2867) );
  nnd2s3 U1072 ( .DIN1(n2869), .DIN2(n6661), .Q(n2865) );
  nnd2s3 U1073 ( .DIN1(n6610), .DIN2(n1960), .Q(n2864) );
  nnd2s3 U1074 ( .DIN1(n6579), .DIN2(n1945), .Q(n2863) );
  nnd4s2 U1075 ( .DIN1(n2870), .DIN2(n2871), .DIN3(n2872), .DIN4(n2873), .Q(
        WX7155) );
  nnd2s3 U1076 ( .DIN1(n2601), .DIN2(n6636), .Q(n2873) );
  xor2s3 U1077 ( .DIN1(n2874), .DIN2(n2875), .Q(n2601) );
  xor2s3 U1078 ( .DIN1(n5187), .DIN2(n5188), .Q(n2875) );
  xnr2s3 U1079 ( .DIN1(n3229), .DIN2(n5189), .Q(n2874) );
  nnd2s3 U1080 ( .DIN1(n2876), .DIN2(n6667), .Q(n2872) );
  nnd2s3 U1081 ( .DIN1(n6610), .DIN2(n1961), .Q(n2871) );
  nnd2s3 U1082 ( .DIN1(n6579), .DIN2(n1944), .Q(n2870) );
  nnd4s2 U1083 ( .DIN1(n2877), .DIN2(n2878), .DIN3(n2879), .DIN4(n2880), .Q(
        WX7153) );
  nnd2s3 U1084 ( .DIN1(n2608), .DIN2(n6630), .Q(n2880) );
  xor2s3 U1085 ( .DIN1(n2881), .DIN2(n2882), .Q(n2608) );
  xor2s3 U1086 ( .DIN1(n5191), .DIN2(n5192), .Q(n2882) );
  xnr2s3 U1087 ( .DIN1(n3230), .DIN2(n5193), .Q(n2881) );
  nnd2s3 U1088 ( .DIN1(n2883), .DIN2(n6661), .Q(n2879) );
  nnd2s3 U1089 ( .DIN1(n6610), .DIN2(n1962), .Q(n2878) );
  nnd2s3 U1090 ( .DIN1(n6579), .DIN2(n1943), .Q(n2877) );
  nnd4s2 U1091 ( .DIN1(n2884), .DIN2(n2885), .DIN3(n2886), .DIN4(n2887), .Q(
        WX7151) );
  nnd2s3 U1092 ( .DIN1(n2615), .DIN2(n6630), .Q(n2887) );
  xor2s3 U1093 ( .DIN1(n2888), .DIN2(n2889), .Q(n2615) );
  xor2s3 U1094 ( .DIN1(n5195), .DIN2(n5196), .Q(n2889) );
  xnr2s3 U1095 ( .DIN1(n3231), .DIN2(n5197), .Q(n2888) );
  nnd2s3 U1096 ( .DIN1(n2890), .DIN2(n6661), .Q(n2886) );
  nnd2s3 U1097 ( .DIN1(n6610), .DIN2(n1963), .Q(n2885) );
  nnd2s3 U1098 ( .DIN1(n6579), .DIN2(n1942), .Q(n2884) );
  nnd4s2 U1099 ( .DIN1(n2891), .DIN2(n2892), .DIN3(n2893), .DIN4(n2894), .Q(
        WX7149) );
  nnd2s3 U1100 ( .DIN1(n2622), .DIN2(n6630), .Q(n2894) );
  xor2s3 U1101 ( .DIN1(n2895), .DIN2(n2896), .Q(n2622) );
  xor2s3 U1102 ( .DIN1(n5199), .DIN2(n5200), .Q(n2896) );
  xnr2s3 U1103 ( .DIN1(n3232), .DIN2(n5201), .Q(n2895) );
  nnd2s3 U1104 ( .DIN1(n2897), .DIN2(n6661), .Q(n2893) );
  nnd2s3 U1105 ( .DIN1(n6610), .DIN2(n1964), .Q(n2892) );
  nnd2s3 U1106 ( .DIN1(n6579), .DIN2(n1941), .Q(n2891) );
  nnd4s2 U1107 ( .DIN1(n2898), .DIN2(n2899), .DIN3(n2900), .DIN4(n2901), .Q(
        WX7147) );
  nnd2s3 U1108 ( .DIN1(n2629), .DIN2(n6630), .Q(n2901) );
  xor2s3 U1109 ( .DIN1(n2902), .DIN2(n2903), .Q(n2629) );
  xor2s3 U1110 ( .DIN1(n5203), .DIN2(n5204), .Q(n2903) );
  xnr2s3 U1111 ( .DIN1(n3233), .DIN2(n5205), .Q(n2902) );
  nnd2s3 U1112 ( .DIN1(n2904), .DIN2(n6661), .Q(n2900) );
  nnd2s3 U1113 ( .DIN1(n6610), .DIN2(n1965), .Q(n2899) );
  nnd2s3 U1114 ( .DIN1(n6579), .DIN2(n1940), .Q(n2898) );
  nnd4s2 U1115 ( .DIN1(n2905), .DIN2(n2906), .DIN3(n2907), .DIN4(n2908), .Q(
        WX7145) );
  nnd2s3 U1116 ( .DIN1(n2636), .DIN2(n6630), .Q(n2908) );
  xor2s3 U1117 ( .DIN1(n2909), .DIN2(n2910), .Q(n2636) );
  xor2s3 U1118 ( .DIN1(n5207), .DIN2(n5208), .Q(n2910) );
  xnr2s3 U1119 ( .DIN1(n3234), .DIN2(n5209), .Q(n2909) );
  nnd2s3 U1120 ( .DIN1(n2911), .DIN2(n6661), .Q(n2907) );
  nnd2s3 U1121 ( .DIN1(n6610), .DIN2(n1966), .Q(n2906) );
  nnd2s3 U1122 ( .DIN1(n6579), .DIN2(n1939), .Q(n2905) );
  nnd4s2 U1123 ( .DIN1(n2912), .DIN2(n2913), .DIN3(n2914), .DIN4(n2915), .Q(
        WX7143) );
  nnd2s3 U1124 ( .DIN1(n2643), .DIN2(n6630), .Q(n2915) );
  xor2s3 U1125 ( .DIN1(n2916), .DIN2(n2917), .Q(n2643) );
  xor2s3 U1126 ( .DIN1(n5211), .DIN2(n5212), .Q(n2917) );
  xnr2s3 U1127 ( .DIN1(n3235), .DIN2(n5213), .Q(n2916) );
  nnd2s3 U1128 ( .DIN1(n2918), .DIN2(n6661), .Q(n2914) );
  nnd2s3 U1129 ( .DIN1(n6610), .DIN2(n1967), .Q(n2913) );
  nnd2s3 U1130 ( .DIN1(n6579), .DIN2(n1938), .Q(n2912) );
  nnd4s2 U1131 ( .DIN1(n2919), .DIN2(n2920), .DIN3(n2921), .DIN4(n2922), .Q(
        WX7141) );
  nnd2s3 U1132 ( .DIN1(n2650), .DIN2(n6630), .Q(n2922) );
  xor2s3 U1133 ( .DIN1(n2923), .DIN2(n2924), .Q(n2650) );
  xor2s3 U1134 ( .DIN1(n5215), .DIN2(n5216), .Q(n2924) );
  xnr2s3 U1135 ( .DIN1(n3236), .DIN2(n5217), .Q(n2923) );
  nnd2s3 U1136 ( .DIN1(n2925), .DIN2(n6660), .Q(n2921) );
  nnd2s3 U1137 ( .DIN1(n6610), .DIN2(n1968), .Q(n2920) );
  nnd2s3 U1138 ( .DIN1(n6579), .DIN2(n1937), .Q(n2919) );
  nor2s3 U1139 ( .DIN1(n6546), .DIN2(n6715), .Q(WX714) );
  nnd4s2 U1140 ( .DIN1(n2926), .DIN2(n2927), .DIN3(n2928), .DIN4(n2929), .Q(
        WX7139) );
  nnd2s3 U1141 ( .DIN1(n2658), .DIN2(n6629), .Q(n2929) );
  xor2s3 U1142 ( .DIN1(n2930), .DIN2(n2931), .Q(n2658) );
  xor2s3 U1143 ( .DIN1(n5221), .DIN2(n2932), .Q(n2931) );
  xor2s3 U1144 ( .DIN1(n5219), .DIN2(n5220), .Q(n2932) );
  xor2s3 U1145 ( .DIN1(n5222), .DIN2(n6688), .Q(n2930) );
  nnd2s3 U1146 ( .DIN1(n2933), .DIN2(n6660), .Q(n2928) );
  nnd2s3 U1147 ( .DIN1(n6609), .DIN2(n1969), .Q(n2927) );
  nnd2s3 U1148 ( .DIN1(n6578), .DIN2(n1936), .Q(n2926) );
  nnd4s2 U1149 ( .DIN1(n2934), .DIN2(n2935), .DIN3(n2936), .DIN4(n2937), .Q(
        WX7137) );
  nnd2s3 U1150 ( .DIN1(n2666), .DIN2(n6629), .Q(n2937) );
  xor2s3 U1151 ( .DIN1(n2938), .DIN2(n2939), .Q(n2666) );
  xor2s3 U1152 ( .DIN1(n5226), .DIN2(n2940), .Q(n2939) );
  xor2s3 U1153 ( .DIN1(n5224), .DIN2(n5225), .Q(n2940) );
  xor2s3 U1154 ( .DIN1(n5227), .DIN2(n6688), .Q(n2938) );
  nnd2s3 U1155 ( .DIN1(n2941), .DIN2(n6660), .Q(n2936) );
  nnd2s3 U1156 ( .DIN1(n6609), .DIN2(n1970), .Q(n2935) );
  nnd2s3 U1157 ( .DIN1(n6578), .DIN2(n1935), .Q(n2934) );
  nnd4s2 U1158 ( .DIN1(n2942), .DIN2(n2943), .DIN3(n2944), .DIN4(n2945), .Q(
        WX7135) );
  nnd2s3 U1159 ( .DIN1(n2674), .DIN2(n6629), .Q(n2945) );
  xor2s3 U1160 ( .DIN1(n2946), .DIN2(n2947), .Q(n2674) );
  xor2s3 U1161 ( .DIN1(n5231), .DIN2(n2948), .Q(n2947) );
  xor2s3 U1162 ( .DIN1(n5229), .DIN2(n5230), .Q(n2948) );
  xor2s3 U1163 ( .DIN1(n5232), .DIN2(n6688), .Q(n2946) );
  nnd2s3 U1164 ( .DIN1(n2949), .DIN2(n6660), .Q(n2944) );
  nnd2s3 U1165 ( .DIN1(n6609), .DIN2(n1971), .Q(n2943) );
  nnd2s3 U1166 ( .DIN1(n6578), .DIN2(n1934), .Q(n2942) );
  nnd4s2 U1167 ( .DIN1(n2950), .DIN2(n2951), .DIN3(n2952), .DIN4(n2953), .Q(
        WX7133) );
  nnd2s3 U1168 ( .DIN1(n2682), .DIN2(n6629), .Q(n2953) );
  xor2s3 U1169 ( .DIN1(n2954), .DIN2(n2955), .Q(n2682) );
  xor2s3 U1170 ( .DIN1(n5236), .DIN2(n2956), .Q(n2955) );
  xor2s3 U1171 ( .DIN1(n5234), .DIN2(n5235), .Q(n2956) );
  xor2s3 U1172 ( .DIN1(n5237), .DIN2(n6688), .Q(n2954) );
  nnd2s3 U1173 ( .DIN1(n2957), .DIN2(n6660), .Q(n2952) );
  nnd2s3 U1174 ( .DIN1(n6609), .DIN2(n1972), .Q(n2951) );
  nnd2s3 U1175 ( .DIN1(n6578), .DIN2(n1933), .Q(n2950) );
  nnd4s2 U1176 ( .DIN1(n2958), .DIN2(n2959), .DIN3(n2960), .DIN4(n2961), .Q(
        WX7131) );
  nnd2s3 U1177 ( .DIN1(n2690), .DIN2(n6629), .Q(n2961) );
  xor2s3 U1178 ( .DIN1(n2962), .DIN2(n2963), .Q(n2690) );
  xor2s3 U1179 ( .DIN1(n5241), .DIN2(n2964), .Q(n2963) );
  xor2s3 U1180 ( .DIN1(n5239), .DIN2(n5240), .Q(n2964) );
  xor2s3 U1181 ( .DIN1(n5242), .DIN2(n6688), .Q(n2962) );
  nnd2s3 U1182 ( .DIN1(n2965), .DIN2(n6660), .Q(n2960) );
  nnd2s3 U1183 ( .DIN1(n6609), .DIN2(n1973), .Q(n2959) );
  nnd2s3 U1184 ( .DIN1(n6578), .DIN2(n1932), .Q(n2958) );
  nnd4s2 U1185 ( .DIN1(n2966), .DIN2(n2967), .DIN3(n2968), .DIN4(n2969), .Q(
        WX7129) );
  nnd2s3 U1186 ( .DIN1(n2698), .DIN2(n6629), .Q(n2969) );
  xor2s3 U1187 ( .DIN1(n2970), .DIN2(n2971), .Q(n2698) );
  xor2s3 U1188 ( .DIN1(n5246), .DIN2(n2972), .Q(n2971) );
  xor2s3 U1189 ( .DIN1(n5244), .DIN2(n5245), .Q(n2972) );
  xor2s3 U1190 ( .DIN1(n5247), .DIN2(n6688), .Q(n2970) );
  nnd2s3 U1191 ( .DIN1(n2973), .DIN2(n6660), .Q(n2968) );
  nnd2s3 U1192 ( .DIN1(n6609), .DIN2(n1974), .Q(n2967) );
  nnd2s3 U1193 ( .DIN1(n6578), .DIN2(n1931), .Q(n2966) );
  nnd4s2 U1194 ( .DIN1(n2974), .DIN2(n2975), .DIN3(n2976), .DIN4(n2977), .Q(
        WX7127) );
  nnd2s3 U1195 ( .DIN1(n2706), .DIN2(n6629), .Q(n2977) );
  xor2s3 U1196 ( .DIN1(n2978), .DIN2(n2979), .Q(n2706) );
  xor2s3 U1197 ( .DIN1(n5251), .DIN2(n2980), .Q(n2979) );
  xor2s3 U1198 ( .DIN1(n5249), .DIN2(n5250), .Q(n2980) );
  xor2s3 U1199 ( .DIN1(n5252), .DIN2(n6688), .Q(n2978) );
  nnd2s3 U1200 ( .DIN1(n2981), .DIN2(n6660), .Q(n2976) );
  nnd2s3 U1201 ( .DIN1(n6609), .DIN2(n1975), .Q(n2975) );
  nnd2s3 U1202 ( .DIN1(n6578), .DIN2(n1930), .Q(n2974) );
  nnd4s2 U1203 ( .DIN1(n2982), .DIN2(n2983), .DIN3(n2984), .DIN4(n2985), .Q(
        WX7125) );
  nnd2s3 U1204 ( .DIN1(n2714), .DIN2(n6629), .Q(n2985) );
  xor2s3 U1205 ( .DIN1(n2986), .DIN2(n2987), .Q(n2714) );
  xor2s3 U1206 ( .DIN1(n5256), .DIN2(n2988), .Q(n2987) );
  xor2s3 U1207 ( .DIN1(n5254), .DIN2(n5255), .Q(n2988) );
  xor2s3 U1208 ( .DIN1(n5257), .DIN2(n6688), .Q(n2986) );
  nnd2s3 U1209 ( .DIN1(n2989), .DIN2(n6660), .Q(n2984) );
  nnd2s3 U1210 ( .DIN1(n6609), .DIN2(n1976), .Q(n2983) );
  nnd2s3 U1211 ( .DIN1(n6578), .DIN2(n1929), .Q(n2982) );
  nnd4s2 U1212 ( .DIN1(n2990), .DIN2(n2991), .DIN3(n2992), .DIN4(n2993), .Q(
        WX7123) );
  nnd2s3 U1213 ( .DIN1(n2722), .DIN2(n6629), .Q(n2993) );
  xor2s3 U1214 ( .DIN1(n2994), .DIN2(n2995), .Q(n2722) );
  xor2s3 U1215 ( .DIN1(n5261), .DIN2(n2996), .Q(n2995) );
  xor2s3 U1216 ( .DIN1(n5259), .DIN2(n5260), .Q(n2996) );
  xor2s3 U1217 ( .DIN1(n5262), .DIN2(n6688), .Q(n2994) );
  nnd2s3 U1218 ( .DIN1(n2997), .DIN2(n6660), .Q(n2992) );
  nnd2s3 U1219 ( .DIN1(n6609), .DIN2(n1977), .Q(n2991) );
  nnd2s3 U1220 ( .DIN1(n6578), .DIN2(n1928), .Q(n2990) );
  nnd4s2 U1221 ( .DIN1(n2998), .DIN2(n2999), .DIN3(n3000), .DIN4(n3001), .Q(
        WX7121) );
  nnd2s3 U1222 ( .DIN1(n2730), .DIN2(n6629), .Q(n3001) );
  xor2s3 U1223 ( .DIN1(n3002), .DIN2(n3003), .Q(n2730) );
  xor2s3 U1224 ( .DIN1(n5266), .DIN2(n3004), .Q(n3003) );
  xor2s3 U1225 ( .DIN1(n5264), .DIN2(n5265), .Q(n3004) );
  xor2s3 U1226 ( .DIN1(n5267), .DIN2(n6688), .Q(n3002) );
  nnd2s3 U1227 ( .DIN1(n3005), .DIN2(n6660), .Q(n3000) );
  nnd2s3 U1228 ( .DIN1(n6609), .DIN2(n1978), .Q(n2999) );
  nnd2s3 U1229 ( .DIN1(n6578), .DIN2(n1927), .Q(n2998) );
  nor2s3 U1230 ( .DIN1(n6481), .DIN2(n6715), .Q(WX712) );
  nnd4s2 U1231 ( .DIN1(n3006), .DIN2(n3007), .DIN3(n3008), .DIN4(n3009), .Q(
        WX7119) );
  nnd2s3 U1232 ( .DIN1(n2738), .DIN2(n6629), .Q(n3009) );
  xor2s3 U1233 ( .DIN1(n3010), .DIN2(n3011), .Q(n2738) );
  xor2s3 U1234 ( .DIN1(n5271), .DIN2(n3012), .Q(n3011) );
  xor2s3 U1235 ( .DIN1(n5269), .DIN2(n5270), .Q(n3012) );
  xor2s3 U1236 ( .DIN1(n5272), .DIN2(n6689), .Q(n3010) );
  nnd2s3 U1237 ( .DIN1(n3013), .DIN2(n6660), .Q(n3008) );
  nnd2s3 U1238 ( .DIN1(n6609), .DIN2(n1979), .Q(n3007) );
  nnd2s3 U1239 ( .DIN1(n6578), .DIN2(n1926), .Q(n3006) );
  nnd4s2 U1240 ( .DIN1(n3014), .DIN2(n3015), .DIN3(n3016), .DIN4(n3017), .Q(
        WX7117) );
  nnd2s3 U1241 ( .DIN1(n2746), .DIN2(n6629), .Q(n3017) );
  xor2s3 U1242 ( .DIN1(n3018), .DIN2(n3019), .Q(n2746) );
  xor2s3 U1243 ( .DIN1(n5276), .DIN2(n3020), .Q(n3019) );
  xor2s3 U1244 ( .DIN1(n5274), .DIN2(n5275), .Q(n3020) );
  xor2s3 U1245 ( .DIN1(n5277), .DIN2(n6689), .Q(n3018) );
  nnd2s3 U1246 ( .DIN1(n3021), .DIN2(n6660), .Q(n3016) );
  nnd2s3 U1247 ( .DIN1(n6609), .DIN2(n1980), .Q(n3015) );
  nnd2s3 U1248 ( .DIN1(n6578), .DIN2(n1925), .Q(n3014) );
  nnd4s2 U1249 ( .DIN1(n3022), .DIN2(n3023), .DIN3(n3024), .DIN4(n3025), .Q(
        WX7115) );
  nnd2s3 U1250 ( .DIN1(n2754), .DIN2(n6629), .Q(n3025) );
  xor2s3 U1251 ( .DIN1(n3026), .DIN2(n3027), .Q(n2754) );
  xor2s3 U1252 ( .DIN1(n5281), .DIN2(n3028), .Q(n3027) );
  xor2s3 U1253 ( .DIN1(n5279), .DIN2(n5280), .Q(n3028) );
  xor2s3 U1254 ( .DIN1(n5282), .DIN2(n6689), .Q(n3026) );
  nnd2s3 U1255 ( .DIN1(n3029), .DIN2(n6659), .Q(n3024) );
  nnd2s3 U1256 ( .DIN1(n6609), .DIN2(n1981), .Q(n3023) );
  nnd2s3 U1257 ( .DIN1(n6578), .DIN2(n1924), .Q(n3022) );
  nnd4s2 U1258 ( .DIN1(n3030), .DIN2(n3031), .DIN3(n3032), .DIN4(n3033), .Q(
        WX7113) );
  nnd2s3 U1259 ( .DIN1(n2762), .DIN2(n6628), .Q(n3033) );
  xor2s3 U1260 ( .DIN1(n3034), .DIN2(n3035), .Q(n2762) );
  xor2s3 U1261 ( .DIN1(n5286), .DIN2(n3036), .Q(n3035) );
  xor2s3 U1262 ( .DIN1(n5284), .DIN2(n5285), .Q(n3036) );
  xor2s3 U1263 ( .DIN1(n5287), .DIN2(n6689), .Q(n3034) );
  nnd2s3 U1264 ( .DIN1(n3037), .DIN2(n6659), .Q(n3032) );
  nnd2s3 U1265 ( .DIN1(n6608), .DIN2(n1982), .Q(n3031) );
  nnd2s3 U1266 ( .DIN1(n6577), .DIN2(n1923), .Q(n3030) );
  nnd4s2 U1267 ( .DIN1(n3038), .DIN2(n3039), .DIN3(n3040), .DIN4(n3041), .Q(
        WX7111) );
  nnd2s3 U1268 ( .DIN1(n2770), .DIN2(n6628), .Q(n3041) );
  xor2s3 U1269 ( .DIN1(n3042), .DIN2(n3043), .Q(n2770) );
  xor2s3 U1270 ( .DIN1(n5291), .DIN2(n3044), .Q(n3043) );
  xor2s3 U1271 ( .DIN1(n5289), .DIN2(n5290), .Q(n3044) );
  xor2s3 U1272 ( .DIN1(n5292), .DIN2(n6689), .Q(n3042) );
  nnd2s3 U1273 ( .DIN1(n3045), .DIN2(n6659), .Q(n3040) );
  nnd2s3 U1274 ( .DIN1(n6608), .DIN2(n1983), .Q(n3039) );
  nnd2s3 U1275 ( .DIN1(n6577), .DIN2(n1922), .Q(n3038) );
  nnd4s2 U1276 ( .DIN1(n3046), .DIN2(n3047), .DIN3(n3048), .DIN4(n3049), .Q(
        WX7109) );
  nnd2s3 U1277 ( .DIN1(n2778), .DIN2(n6628), .Q(n3049) );
  xor2s3 U1278 ( .DIN1(n3050), .DIN2(n3051), .Q(n2778) );
  xor2s3 U1279 ( .DIN1(n5296), .DIN2(n3052), .Q(n3051) );
  xor2s3 U1280 ( .DIN1(n5294), .DIN2(n5295), .Q(n3052) );
  xor2s3 U1281 ( .DIN1(n5297), .DIN2(n6689), .Q(n3050) );
  nnd2s3 U1282 ( .DIN1(n3053), .DIN2(n6659), .Q(n3048) );
  nnd2s3 U1283 ( .DIN1(n6608), .DIN2(n1984), .Q(n3047) );
  nnd2s3 U1284 ( .DIN1(n6577), .DIN2(n1921), .Q(n3046) );
  nor2s3 U1285 ( .DIN1(n6549), .DIN2(n6715), .Q(WX710) );
  nor2s3 U1286 ( .DIN1(n6533), .DIN2(n6715), .Q(WX708) );
  nnd4s2 U1287 ( .DIN1(n3054), .DIN2(n3055), .DIN3(n3056), .DIN4(n3057), .Q(
        WX706) );
  nnd2s3 U1288 ( .DIN1(n3058), .DIN2(n6628), .Q(n3057) );
  nnd2s3 U1289 ( .DIN1(n6608), .DIN2(n2273), .Q(n3056) );
  nnd2s3 U1290 ( .DIN1(n6577), .DIN2(n2272), .Q(n3055) );
  nnd2s3 U1291 ( .DIN1(n6657), .DIN2(n3059), .Q(n3054) );
  nnd4s2 U1292 ( .DIN1(n3060), .DIN2(n3061), .DIN3(n3062), .DIN4(n3063), .Q(
        WX704) );
  nnd2s3 U1293 ( .DIN1(n3064), .DIN2(n6628), .Q(n3063) );
  nnd2s3 U1294 ( .DIN1(n6608), .DIN2(n2274), .Q(n3062) );
  nnd2s3 U1295 ( .DIN1(n6577), .DIN2(n2271), .Q(n3061) );
  nnd2s3 U1296 ( .DIN1(n6658), .DIN2(n3065), .Q(n3060) );
  nnd4s2 U1297 ( .DIN1(n3066), .DIN2(n3067), .DIN3(n3068), .DIN4(n3069), .Q(
        WX702) );
  nnd2s3 U1298 ( .DIN1(n3070), .DIN2(n6628), .Q(n3069) );
  nnd2s3 U1299 ( .DIN1(n6608), .DIN2(n2275), .Q(n3068) );
  nnd2s3 U1300 ( .DIN1(n6577), .DIN2(n2270), .Q(n3067) );
  nnd2s3 U1301 ( .DIN1(n6657), .DIN2(n3071), .Q(n3066) );
  nor2s3 U1302 ( .DIN1(n6790), .DIN2(n1984), .Q(WX7011) );
  nor2s3 U1303 ( .DIN1(n5300), .DIN2(n6715), .Q(WX7009) );
  nor2s3 U1304 ( .DIN1(n5301), .DIN2(n6715), .Q(WX7007) );
  nor2s3 U1305 ( .DIN1(n5302), .DIN2(n6715), .Q(WX7005) );
  nor2s3 U1306 ( .DIN1(n5303), .DIN2(n6715), .Q(WX7003) );
  nor2s3 U1307 ( .DIN1(n5304), .DIN2(n6715), .Q(WX7001) );
  nnd4s2 U1308 ( .DIN1(n3072), .DIN2(n3073), .DIN3(n3074), .DIN4(n3075), .Q(
        WX700) );
  nnd2s3 U1309 ( .DIN1(n3076), .DIN2(n6628), .Q(n3075) );
  nnd2s3 U1310 ( .DIN1(n6608), .DIN2(n2276), .Q(n3074) );
  nnd2s3 U1311 ( .DIN1(n6577), .DIN2(n2269), .Q(n3073) );
  nnd2s3 U1312 ( .DIN1(n6658), .DIN2(n3077), .Q(n3072) );
  nor2s3 U1313 ( .DIN1(n5305), .DIN2(n6715), .Q(WX6999) );
  nor2s3 U1314 ( .DIN1(n5306), .DIN2(n6715), .Q(WX6997) );
  nor2s3 U1315 ( .DIN1(n5307), .DIN2(n6714), .Q(WX6995) );
  nor2s3 U1316 ( .DIN1(n5308), .DIN2(n6714), .Q(WX6993) );
  nor2s3 U1317 ( .DIN1(n5309), .DIN2(n6714), .Q(WX6991) );
  nor2s3 U1318 ( .DIN1(n5310), .DIN2(n6714), .Q(WX6989) );
  nor2s3 U1319 ( .DIN1(n5311), .DIN2(n6714), .Q(WX6987) );
  nor2s3 U1320 ( .DIN1(n5312), .DIN2(n6714), .Q(WX6985) );
  nor2s3 U1321 ( .DIN1(n5313), .DIN2(n6714), .Q(WX6983) );
  nor2s3 U1322 ( .DIN1(n5314), .DIN2(n6714), .Q(WX6981) );
  nnd4s2 U1323 ( .DIN1(n3078), .DIN2(n3079), .DIN3(n3080), .DIN4(n3081), .Q(
        WX698) );
  nnd2s3 U1324 ( .DIN1(n3082), .DIN2(n6628), .Q(n3081) );
  nnd2s3 U1325 ( .DIN1(n6608), .DIN2(n2277), .Q(n3080) );
  nnd2s3 U1326 ( .DIN1(n6577), .DIN2(n2268), .Q(n3079) );
  nnd2s3 U1327 ( .DIN1(n6656), .DIN2(n3083), .Q(n3078) );
  nor2s3 U1328 ( .DIN1(n5315), .DIN2(n6714), .Q(WX6979) );
  nor2s3 U1329 ( .DIN1(n5316), .DIN2(n6714), .Q(WX6977) );
  nor2s3 U1330 ( .DIN1(n5317), .DIN2(n6714), .Q(WX6975) );
  nor2s3 U1331 ( .DIN1(n5318), .DIN2(n6714), .Q(WX6973) );
  nor2s3 U1332 ( .DIN1(n5319), .DIN2(n6713), .Q(WX6971) );
  nor2s3 U1333 ( .DIN1(n5320), .DIN2(n6713), .Q(WX6969) );
  nor2s3 U1334 ( .DIN1(n5321), .DIN2(n6713), .Q(WX6967) );
  nor2s3 U1335 ( .DIN1(n5322), .DIN2(n6713), .Q(WX6965) );
  nor2s3 U1336 ( .DIN1(n5323), .DIN2(n6713), .Q(WX6963) );
  nor2s3 U1337 ( .DIN1(n5324), .DIN2(n6713), .Q(WX6961) );
  nnd4s2 U1338 ( .DIN1(n3084), .DIN2(n3085), .DIN3(n3086), .DIN4(n3087), .Q(
        WX696) );
  nnd2s3 U1339 ( .DIN1(n3088), .DIN2(n6628), .Q(n3087) );
  nnd2s3 U1340 ( .DIN1(n6608), .DIN2(n2278), .Q(n3086) );
  nnd2s3 U1341 ( .DIN1(n6577), .DIN2(n2267), .Q(n3085) );
  nnd2s3 U1342 ( .DIN1(n6658), .DIN2(n3089), .Q(n3084) );
  nor2s3 U1343 ( .DIN1(n5325), .DIN2(n6713), .Q(WX6959) );
  nor2s3 U1344 ( .DIN1(n5326), .DIN2(n6713), .Q(WX6957) );
  nor2s3 U1345 ( .DIN1(n5327), .DIN2(n6713), .Q(WX6955) );
  nor2s3 U1346 ( .DIN1(n5328), .DIN2(n6713), .Q(WX6953) );
  nor2s3 U1347 ( .DIN1(n5329), .DIN2(n6713), .Q(WX6951) );
  nor2s3 U1348 ( .DIN1(n5330), .DIN2(n6713), .Q(WX6949) );
  nnd4s2 U1349 ( .DIN1(n3090), .DIN2(n3091), .DIN3(n3092), .DIN4(n3093), .Q(
        WX694) );
  nnd2s3 U1350 ( .DIN1(n3094), .DIN2(n6628), .Q(n3093) );
  nnd2s3 U1351 ( .DIN1(n6608), .DIN2(n2279), .Q(n3092) );
  nnd2s3 U1352 ( .DIN1(n6577), .DIN2(n2266), .Q(n3091) );
  nnd2s3 U1353 ( .DIN1(n6656), .DIN2(n3095), .Q(n3090) );
  nnd4s2 U1354 ( .DIN1(n3096), .DIN2(n3097), .DIN3(n3098), .DIN4(n3099), .Q(
        WX692) );
  nnd2s3 U1355 ( .DIN1(n3100), .DIN2(n6628), .Q(n3099) );
  nnd2s3 U1356 ( .DIN1(n6608), .DIN2(n2280), .Q(n3098) );
  nnd2s3 U1357 ( .DIN1(n6577), .DIN2(n2265), .Q(n3097) );
  nnd2s3 U1358 ( .DIN1(n6658), .DIN2(n3101), .Q(n3096) );
  nnd4s2 U1359 ( .DIN1(n3102), .DIN2(n3103), .DIN3(n3104), .DIN4(n3105), .Q(
        WX690) );
  nnd2s3 U1360 ( .DIN1(n3106), .DIN2(n6630), .Q(n3105) );
  nnd2s3 U1361 ( .DIN1(n6608), .DIN2(n2281), .Q(n3104) );
  nnd2s3 U1362 ( .DIN1(n6577), .DIN2(n2264), .Q(n3103) );
  nnd2s3 U1363 ( .DIN1(n6656), .DIN2(n3107), .Q(n3102) );
  nnd4s2 U1364 ( .DIN1(n3108), .DIN2(n3109), .DIN3(n3110), .DIN4(n3111), .Q(
        WX688) );
  nnd2s3 U1365 ( .DIN1(n3112), .DIN2(n6628), .Q(n3111) );
  nnd2s3 U1366 ( .DIN1(n6608), .DIN2(n2282), .Q(n3110) );
  nnd2s3 U1367 ( .DIN1(n6577), .DIN2(n2263), .Q(n3109) );
  nnd2s3 U1368 ( .DIN1(n6658), .DIN2(n3113), .Q(n3108) );
  nnd4s2 U1369 ( .DIN1(n3114), .DIN2(n3115), .DIN3(n3116), .DIN4(n3117), .Q(
        WX686) );
  nnd2s3 U1370 ( .DIN1(n3118), .DIN2(n6627), .Q(n3117) );
  nnd2s3 U1371 ( .DIN1(n6607), .DIN2(n2283), .Q(n3116) );
  nnd2s3 U1372 ( .DIN1(n6576), .DIN2(n2262), .Q(n3115) );
  nnd2s3 U1373 ( .DIN1(n6657), .DIN2(n3119), .Q(n3114) );
  nnd4s2 U1374 ( .DIN1(n3120), .DIN2(n3121), .DIN3(n3122), .DIN4(n3123), .Q(
        WX684) );
  nnd2s3 U1375 ( .DIN1(n3124), .DIN2(n6627), .Q(n3123) );
  nnd2s3 U1376 ( .DIN1(n6607), .DIN2(n2284), .Q(n3122) );
  nnd2s3 U1377 ( .DIN1(n6576), .DIN2(n2261), .Q(n3121) );
  nnd2s3 U1378 ( .DIN1(n6658), .DIN2(n3125), .Q(n3120) );
  nnd4s2 U1379 ( .DIN1(n3126), .DIN2(n3127), .DIN3(n3128), .DIN4(n3129), .Q(
        WX682) );
  nnd2s3 U1380 ( .DIN1(n3130), .DIN2(n6627), .Q(n3129) );
  nnd2s3 U1381 ( .DIN1(n6607), .DIN2(n2285), .Q(n3128) );
  nnd2s3 U1382 ( .DIN1(n6576), .DIN2(n2260), .Q(n3127) );
  nnd2s3 U1383 ( .DIN1(n6656), .DIN2(n3131), .Q(n3126) );
  nnd4s2 U1384 ( .DIN1(n3132), .DIN2(n3133), .DIN3(n3134), .DIN4(n3135), .Q(
        WX680) );
  nnd2s3 U1385 ( .DIN1(n3136), .DIN2(n6627), .Q(n3135) );
  nnd2s3 U1386 ( .DIN1(n6607), .DIN2(n2286), .Q(n3134) );
  nnd2s3 U1387 ( .DIN1(n6576), .DIN2(n2259), .Q(n3133) );
  nnd2s3 U1388 ( .DIN1(n6658), .DIN2(n3137), .Q(n3132) );
  nnd4s2 U1389 ( .DIN1(n3138), .DIN2(n3139), .DIN3(n3140), .DIN4(n3141), .Q(
        WX678) );
  nnd2s3 U1390 ( .DIN1(n3142), .DIN2(n6627), .Q(n3141) );
  nnd2s3 U1391 ( .DIN1(n6607), .DIN2(n2287), .Q(n3140) );
  nnd2s3 U1392 ( .DIN1(n6576), .DIN2(n2258), .Q(n3139) );
  nnd2s3 U1393 ( .DIN1(n6657), .DIN2(n3143), .Q(n3138) );
  nnd4s2 U1394 ( .DIN1(n3144), .DIN2(n3145), .DIN3(n3146), .DIN4(n3147), .Q(
        WX676) );
  nnd2s3 U1395 ( .DIN1(n3148), .DIN2(n6627), .Q(n3147) );
  nnd2s3 U1396 ( .DIN1(n6607), .DIN2(n2288), .Q(n3146) );
  nnd2s3 U1397 ( .DIN1(n6576), .DIN2(n2257), .Q(n3145) );
  nnd2s3 U1398 ( .DIN1(n6657), .DIN2(n3149), .Q(n3144) );
  nnd4s2 U1399 ( .DIN1(n3150), .DIN2(n3151), .DIN3(n3152), .DIN4(n3153), .Q(
        WX674) );
  nnd2s3 U1400 ( .DIN1(n3154), .DIN2(n6627), .Q(n3153) );
  nnd2s3 U1401 ( .DIN1(n6607), .DIN2(n2289), .Q(n3152) );
  nnd2s3 U1402 ( .DIN1(n6576), .DIN2(n2256), .Q(n3151) );
  nnd2s3 U1403 ( .DIN1(n6657), .DIN2(n3155), .Q(n3150) );
  nnd4s2 U1404 ( .DIN1(n3156), .DIN2(n3157), .DIN3(n3158), .DIN4(n3159), .Q(
        WX672) );
  nnd2s3 U1405 ( .DIN1(n3160), .DIN2(n6627), .Q(n3159) );
  nnd2s3 U1406 ( .DIN1(n6607), .DIN2(n2290), .Q(n3158) );
  nnd2s3 U1407 ( .DIN1(n6576), .DIN2(n2255), .Q(n3157) );
  nnd2s3 U1408 ( .DIN1(n6657), .DIN2(n3161), .Q(n3156) );
  nnd4s2 U1409 ( .DIN1(n3162), .DIN2(n3163), .DIN3(n3164), .DIN4(n3165), .Q(
        WX670) );
  nnd2s3 U1410 ( .DIN1(n3166), .DIN2(n6627), .Q(n3165) );
  nnd2s3 U1411 ( .DIN1(n6607), .DIN2(n2291), .Q(n3164) );
  nnd2s3 U1412 ( .DIN1(n6576), .DIN2(n2254), .Q(n3163) );
  nnd2s3 U1413 ( .DIN1(n6656), .DIN2(n3167), .Q(n3162) );
  nnd4s2 U1414 ( .DIN1(n3168), .DIN2(n3169), .DIN3(n3170), .DIN4(n3171), .Q(
        WX668) );
  nnd2s3 U1415 ( .DIN1(n3172), .DIN2(n6627), .Q(n3171) );
  nnd2s3 U1416 ( .DIN1(n6607), .DIN2(n2292), .Q(n3170) );
  nnd2s3 U1417 ( .DIN1(n6576), .DIN2(n2253), .Q(n3169) );
  nnd2s3 U1418 ( .DIN1(n6657), .DIN2(n3173), .Q(n3168) );
  nnd4s2 U1419 ( .DIN1(n3174), .DIN2(n3175), .DIN3(n3176), .DIN4(n3177), .Q(
        WX666) );
  nnd2s3 U1420 ( .DIN1(n3178), .DIN2(n6627), .Q(n3177) );
  nnd2s3 U1421 ( .DIN1(n6607), .DIN2(n2293), .Q(n3176) );
  nnd2s3 U1422 ( .DIN1(n6576), .DIN2(n2252), .Q(n3175) );
  nnd2s3 U1423 ( .DIN1(n6657), .DIN2(n3179), .Q(n3174) );
  nnd4s2 U1424 ( .DIN1(n3180), .DIN2(n3181), .DIN3(n3182), .DIN4(n3183), .Q(
        WX664) );
  nnd2s3 U1425 ( .DIN1(n3184), .DIN2(n6627), .Q(n3183) );
  nnd2s3 U1426 ( .DIN1(n6607), .DIN2(n2294), .Q(n3182) );
  nnd2s3 U1427 ( .DIN1(n6576), .DIN2(n2251), .Q(n3181) );
  nnd2s3 U1428 ( .DIN1(n6657), .DIN2(n3185), .Q(n3180) );
  nnd4s2 U1429 ( .DIN1(n3186), .DIN2(n3187), .DIN3(n3188), .DIN4(n3189), .Q(
        WX662) );
  nnd2s3 U1430 ( .DIN1(n3190), .DIN2(n6626), .Q(n3189) );
  nnd2s3 U1431 ( .DIN1(n6607), .DIN2(n2295), .Q(n3188) );
  nnd2s3 U1432 ( .DIN1(n6576), .DIN2(n2250), .Q(n3187) );
  nnd2s3 U1433 ( .DIN1(n6656), .DIN2(n3191), .Q(n3186) );
  nnd4s2 U1434 ( .DIN1(n3192), .DIN2(n3193), .DIN3(n3194), .DIN4(n3195), .Q(
        WX660) );
  nnd2s3 U1435 ( .DIN1(n3196), .DIN2(n6627), .Q(n3195) );
  nnd2s3 U1436 ( .DIN1(n6606), .DIN2(n2296), .Q(n3194) );
  nnd2s3 U1437 ( .DIN1(n6575), .DIN2(n2249), .Q(n3193) );
  nnd2s3 U1438 ( .DIN1(n6657), .DIN2(n3197), .Q(n3192) );
  nnd4s2 U1439 ( .DIN1(n3198), .DIN2(n3199), .DIN3(n3200), .DIN4(n3201), .Q(
        WX658) );
  nnd2s3 U1440 ( .DIN1(n3202), .DIN2(n6626), .Q(n3201) );
  nnd2s3 U1441 ( .DIN1(n6606), .DIN2(n2297), .Q(n3200) );
  nnd2s3 U1442 ( .DIN1(n6575), .DIN2(n2248), .Q(n3199) );
  nnd2s3 U1443 ( .DIN1(n6656), .DIN2(n3203), .Q(n3198) );
  nnd4s2 U1444 ( .DIN1(n3204), .DIN2(n3333), .DIN3(n3334), .DIN4(n3335), .Q(
        WX656) );
  nnd2s3 U1445 ( .DIN1(n3336), .DIN2(n6626), .Q(n3335) );
  nnd2s3 U1446 ( .DIN1(n6606), .DIN2(n2298), .Q(n3334) );
  nnd2s3 U1447 ( .DIN1(n6575), .DIN2(n2247), .Q(n3333) );
  nnd2s3 U1448 ( .DIN1(n6657), .DIN2(n3337), .Q(n3204) );
  nnd4s2 U1449 ( .DIN1(n3338), .DIN2(n3339), .DIN3(n3340), .DIN4(n3341), .Q(
        WX654) );
  nnd2s3 U1450 ( .DIN1(n3342), .DIN2(n6626), .Q(n3341) );
  nnd2s3 U1451 ( .DIN1(n6606), .DIN2(n2299), .Q(n3340) );
  nnd2s3 U1452 ( .DIN1(n6575), .DIN2(n2246), .Q(n3339) );
  nnd2s3 U1453 ( .DIN1(n6656), .DIN2(n3343), .Q(n3338) );
  nnd4s2 U1454 ( .DIN1(n3344), .DIN2(n3345), .DIN3(n3346), .DIN4(n3347), .Q(
        WX652) );
  nnd2s3 U1455 ( .DIN1(n3348), .DIN2(n6626), .Q(n3347) );
  nnd2s3 U1456 ( .DIN1(n6606), .DIN2(n2300), .Q(n3346) );
  nnd2s3 U1457 ( .DIN1(n6575), .DIN2(n2245), .Q(n3345) );
  nnd2s3 U1458 ( .DIN1(n6656), .DIN2(n3349), .Q(n3344) );
  nnd4s2 U1459 ( .DIN1(n3350), .DIN2(n3351), .DIN3(n3352), .DIN4(n3353), .Q(
        WX650) );
  nnd2s3 U1460 ( .DIN1(n3354), .DIN2(n6626), .Q(n3353) );
  nnd2s3 U1461 ( .DIN1(n6606), .DIN2(n2301), .Q(n3352) );
  nnd2s3 U1462 ( .DIN1(n6575), .DIN2(n2244), .Q(n3351) );
  nnd2s3 U1463 ( .DIN1(n6656), .DIN2(n3355), .Q(n3350) );
  nor2s3 U1464 ( .DIN1(n6796), .DIN2(n3356), .Q(WX6498) );
  xor2s3 U1465 ( .DIN1(n5469), .DIN2(n5649), .Q(n3356) );
  nor2s3 U1466 ( .DIN1(n6796), .DIN2(n3357), .Q(WX6496) );
  xor2s3 U1467 ( .DIN1(n5464), .DIN2(n5644), .Q(n3357) );
  nor2s3 U1468 ( .DIN1(n6797), .DIN2(n3358), .Q(WX6494) );
  xor2s3 U1469 ( .DIN1(n5459), .DIN2(n5639), .Q(n3358) );
  nor2s3 U1470 ( .DIN1(n6797), .DIN2(n3359), .Q(WX6492) );
  xor2s3 U1471 ( .DIN1(n5454), .DIN2(n5634), .Q(n3359) );
  nor2s3 U1472 ( .DIN1(n6798), .DIN2(n3360), .Q(WX6490) );
  xor2s3 U1473 ( .DIN1(n5449), .DIN2(n5629), .Q(n3360) );
  nor2s3 U1474 ( .DIN1(n6798), .DIN2(n3361), .Q(WX6488) );
  xor2s3 U1475 ( .DIN1(n5444), .DIN2(n5624), .Q(n3361) );
  nor2s3 U1476 ( .DIN1(n6798), .DIN2(n3362), .Q(WX6486) );
  xor2s3 U1477 ( .DIN1(n5439), .DIN2(n5619), .Q(n3362) );
  nor2s3 U1478 ( .DIN1(n6798), .DIN2(n3363), .Q(WX6484) );
  xor2s3 U1479 ( .DIN1(n5434), .DIN2(n5614), .Q(n3363) );
  nor2s3 U1480 ( .DIN1(n6798), .DIN2(n3364), .Q(WX6482) );
  xor2s3 U1481 ( .DIN1(n5429), .DIN2(n5609), .Q(n3364) );
  nor2s3 U1482 ( .DIN1(n6798), .DIN2(n3365), .Q(WX6480) );
  xor2s3 U1483 ( .DIN1(n5424), .DIN2(n5604), .Q(n3365) );
  nnd4s2 U1484 ( .DIN1(n3366), .DIN2(n3367), .DIN3(n3368), .DIN4(n3369), .Q(
        WX648) );
  nnd2s3 U1485 ( .DIN1(n3370), .DIN2(n6626), .Q(n3369) );
  nnd2s3 U1486 ( .DIN1(n6606), .DIN2(n2302), .Q(n3368) );
  nnd2s3 U1487 ( .DIN1(n6575), .DIN2(n2243), .Q(n3367) );
  nnd2s3 U1488 ( .DIN1(n6656), .DIN2(n3371), .Q(n3366) );
  nor2s3 U1489 ( .DIN1(n6799), .DIN2(n3372), .Q(WX6478) );
  xor2s3 U1490 ( .DIN1(n5419), .DIN2(n5599), .Q(n3372) );
  nor2s3 U1491 ( .DIN1(n6799), .DIN2(n3373), .Q(WX6476) );
  xor2s3 U1492 ( .DIN1(n5414), .DIN2(n5594), .Q(n3373) );
  nor2s3 U1493 ( .DIN1(n6799), .DIN2(n3374), .Q(WX6474) );
  xor2s3 U1494 ( .DIN1(n5409), .DIN2(n5589), .Q(n3374) );
  nor2s3 U1495 ( .DIN1(n6799), .DIN2(n3375), .Q(WX6472) );
  xor2s3 U1496 ( .DIN1(n5404), .DIN2(n5584), .Q(n3375) );
  nor2s3 U1497 ( .DIN1(n6799), .DIN2(n3376), .Q(WX6470) );
  xor2s3 U1498 ( .DIN1(n5399), .DIN2(n5579), .Q(n3376) );
  nor2s3 U1499 ( .DIN1(n3377), .DIN2(n6712), .Q(WX6468) );
  xnr2s3 U1500 ( .DIN1(n5574), .DIN2(n3378), .Q(n3377) );
  xor2s3 U1501 ( .DIN1(n5394), .DIN2(n5474), .Q(n3378) );
  nor2s3 U1502 ( .DIN1(n6799), .DIN2(n3379), .Q(WX6466) );
  xor2s3 U1503 ( .DIN1(n5390), .DIN2(n3268), .Q(n3379) );
  nor2s3 U1504 ( .DIN1(n6799), .DIN2(n3380), .Q(WX6464) );
  xor2s3 U1505 ( .DIN1(n5386), .DIN2(n3267), .Q(n3380) );
  nor2s3 U1506 ( .DIN1(n6799), .DIN2(n3381), .Q(WX6462) );
  xor2s3 U1507 ( .DIN1(n5382), .DIN2(n3266), .Q(n3381) );
  nor2s3 U1508 ( .DIN1(n6799), .DIN2(n3382), .Q(WX6460) );
  xor2s3 U1509 ( .DIN1(n5378), .DIN2(n3265), .Q(n3382) );
  nnd4s2 U1510 ( .DIN1(n3383), .DIN2(n3384), .DIN3(n3385), .DIN4(n3386), .Q(
        WX646) );
  nnd2s3 U1511 ( .DIN1(n3387), .DIN2(n6626), .Q(n3386) );
  nnd2s3 U1512 ( .DIN1(n6606), .DIN2(n2303), .Q(n3385) );
  nnd2s3 U1513 ( .DIN1(n6575), .DIN2(n2242), .Q(n3384) );
  nnd2s3 U1514 ( .DIN1(n6656), .DIN2(n3388), .Q(n3383) );
  nor2s3 U1515 ( .DIN1(n3389), .DIN2(n6712), .Q(WX6458) );
  xnr2s3 U1516 ( .DIN1(n3264), .DIN2(n3390), .Q(n3389) );
  xor2s3 U1517 ( .DIN1(n5374), .DIN2(n5474), .Q(n3390) );
  nor2s3 U1518 ( .DIN1(n6799), .DIN2(n3391), .Q(WX6456) );
  xor2s3 U1519 ( .DIN1(n5370), .DIN2(n3263), .Q(n3391) );
  nor2s3 U1520 ( .DIN1(n6799), .DIN2(n3392), .Q(WX6454) );
  xor2s3 U1521 ( .DIN1(n5366), .DIN2(n3262), .Q(n3392) );
  nor2s3 U1522 ( .DIN1(n6799), .DIN2(n3393), .Q(WX6452) );
  xor2s3 U1523 ( .DIN1(n5362), .DIN2(n3261), .Q(n3393) );
  nor2s3 U1524 ( .DIN1(n6799), .DIN2(n3394), .Q(WX6450) );
  xor2s3 U1525 ( .DIN1(n5358), .DIN2(n3260), .Q(n3394) );
  nor2s3 U1526 ( .DIN1(n6800), .DIN2(n3395), .Q(WX6448) );
  xor2s3 U1527 ( .DIN1(n5354), .DIN2(n3259), .Q(n3395) );
  nor2s3 U1528 ( .DIN1(n6800), .DIN2(n3396), .Q(WX6446) );
  xor2s3 U1529 ( .DIN1(n5350), .DIN2(n3258), .Q(n3396) );
  nor2s3 U1530 ( .DIN1(n3397), .DIN2(n6712), .Q(WX6444) );
  xnr2s3 U1531 ( .DIN1(n3257), .DIN2(n3398), .Q(n3397) );
  xor2s3 U1532 ( .DIN1(n5346), .DIN2(n5474), .Q(n3398) );
  nor2s3 U1533 ( .DIN1(n6800), .DIN2(n3399), .Q(WX6442) );
  xor2s3 U1534 ( .DIN1(n5342), .DIN2(n3256), .Q(n3399) );
  nor2s3 U1535 ( .DIN1(n6800), .DIN2(n3400), .Q(WX6440) );
  xor2s3 U1536 ( .DIN1(n5338), .DIN2(n3255), .Q(n3400) );
  nnd4s2 U1537 ( .DIN1(n3401), .DIN2(n3402), .DIN3(n3403), .DIN4(n3404), .Q(
        WX644) );
  nnd2s3 U1538 ( .DIN1(n3405), .DIN2(n6626), .Q(n3404) );
  nnd2s3 U1539 ( .DIN1(n6606), .DIN2(n2304), .Q(n3403) );
  nnd2s3 U1540 ( .DIN1(n6575), .DIN2(n2241), .Q(n3402) );
  nnd2s3 U1541 ( .DIN1(n6656), .DIN2(n3406), .Q(n3401) );
  nor2s3 U1542 ( .DIN1(n6800), .DIN2(n3407), .Q(WX6438) );
  xor2s3 U1543 ( .DIN1(n5334), .DIN2(n3254), .Q(n3407) );
  nor2s3 U1544 ( .DIN1(n6800), .DIN2(n3408), .Q(WX6436) );
  xor2s3 U1545 ( .DIN1(n5474), .DIN2(n3253), .Q(n3408) );
  nor2s3 U1546 ( .DIN1(n5509), .DIN2(n6712), .Q(WX6070) );
  nor2s3 U1547 ( .DIN1(n5513), .DIN2(n6712), .Q(WX6068) );
  nor2s3 U1548 ( .DIN1(n5517), .DIN2(n6712), .Q(WX6066) );
  nor2s3 U1549 ( .DIN1(n5521), .DIN2(n6712), .Q(WX6064) );
  nor2s3 U1550 ( .DIN1(n5525), .DIN2(n6712), .Q(WX6062) );
  nor2s3 U1551 ( .DIN1(n5529), .DIN2(n6712), .Q(WX6060) );
  nor2s3 U1552 ( .DIN1(n5533), .DIN2(n6712), .Q(WX6058) );
  nor2s3 U1553 ( .DIN1(n5537), .DIN2(n6712), .Q(WX6056) );
  nor2s3 U1554 ( .DIN1(n5541), .DIN2(n6717), .Q(WX6054) );
  nor2s3 U1555 ( .DIN1(n5545), .DIN2(n6734), .Q(WX6052) );
  nor2s3 U1556 ( .DIN1(n5549), .DIN2(n6733), .Q(WX6050) );
  nor2s3 U1557 ( .DIN1(n5553), .DIN2(n6733), .Q(WX6048) );
  nor2s3 U1558 ( .DIN1(n5557), .DIN2(n6733), .Q(WX6046) );
  nor2s3 U1559 ( .DIN1(n5561), .DIN2(n6733), .Q(WX6044) );
  nor2s3 U1560 ( .DIN1(n5565), .DIN2(n6733), .Q(WX6042) );
  nor2s3 U1561 ( .DIN1(n5569), .DIN2(n6733), .Q(WX6040) );
  nor2s3 U1562 ( .DIN1(n5573), .DIN2(n6733), .Q(WX6038) );
  nor2s3 U1563 ( .DIN1(n5578), .DIN2(n6733), .Q(WX6036) );
  nor2s3 U1564 ( .DIN1(n5583), .DIN2(n6733), .Q(WX6034) );
  nor2s3 U1565 ( .DIN1(n5588), .DIN2(n6733), .Q(WX6032) );
  nor2s3 U1566 ( .DIN1(n5593), .DIN2(n6733), .Q(WX6030) );
  nor2s3 U1567 ( .DIN1(n5598), .DIN2(n6733), .Q(WX6028) );
  nor2s3 U1568 ( .DIN1(n5603), .DIN2(n6732), .Q(WX6026) );
  nor2s3 U1569 ( .DIN1(n5608), .DIN2(n6732), .Q(WX6024) );
  nor2s3 U1570 ( .DIN1(n5613), .DIN2(n6732), .Q(WX6022) );
  nor2s3 U1571 ( .DIN1(n5618), .DIN2(n6732), .Q(WX6020) );
  nor2s3 U1572 ( .DIN1(n5623), .DIN2(n6732), .Q(WX6018) );
  nor2s3 U1573 ( .DIN1(n5628), .DIN2(n6732), .Q(WX6016) );
  nor2s3 U1574 ( .DIN1(n5633), .DIN2(n6732), .Q(WX6014) );
  nor2s3 U1575 ( .DIN1(n5638), .DIN2(n6732), .Q(WX6012) );
  nor2s3 U1576 ( .DIN1(n5643), .DIN2(n6732), .Q(WX6010) );
  nor2s3 U1577 ( .DIN1(n5648), .DIN2(n6732), .Q(WX6008) );
  nor2s3 U1578 ( .DIN1(n5508), .DIN2(n6732), .Q(WX6006) );
  nor2s3 U1579 ( .DIN1(n5512), .DIN2(n6732), .Q(WX6004) );
  nor2s3 U1580 ( .DIN1(n5516), .DIN2(n6731), .Q(WX6002) );
  nor2s3 U1581 ( .DIN1(n5520), .DIN2(n6731), .Q(WX6000) );
  nor2s3 U1582 ( .DIN1(n5524), .DIN2(n6731), .Q(WX5998) );
  nor2s3 U1583 ( .DIN1(n5528), .DIN2(n6731), .Q(WX5996) );
  nor2s3 U1584 ( .DIN1(n5532), .DIN2(n6731), .Q(WX5994) );
  nor2s3 U1585 ( .DIN1(n5536), .DIN2(n6731), .Q(WX5992) );
  nor2s3 U1586 ( .DIN1(n5540), .DIN2(n6731), .Q(WX5990) );
  nor2s3 U1587 ( .DIN1(n5544), .DIN2(n6731), .Q(WX5988) );
  nor2s3 U1588 ( .DIN1(n5548), .DIN2(n6731), .Q(WX5986) );
  nor2s3 U1589 ( .DIN1(n5552), .DIN2(n6731), .Q(WX5984) );
  nor2s3 U1590 ( .DIN1(n5556), .DIN2(n6731), .Q(WX5982) );
  nor2s3 U1591 ( .DIN1(n5560), .DIN2(n6731), .Q(WX5980) );
  nor2s3 U1592 ( .DIN1(n5564), .DIN2(n6730), .Q(WX5978) );
  nor2s3 U1593 ( .DIN1(n5568), .DIN2(n6730), .Q(WX5976) );
  and2s3 U1594 ( .DIN1(RESET), .DIN2(n5572), .Q(WX5974) );
  and2s3 U1595 ( .DIN1(RESET), .DIN2(n5577), .Q(WX5972) );
  and2s3 U1596 ( .DIN1(RESET), .DIN2(n5582), .Q(WX5970) );
  and2s3 U1597 ( .DIN1(RESET), .DIN2(n5587), .Q(WX5968) );
  and2s3 U1598 ( .DIN1(RESET), .DIN2(n5592), .Q(WX5966) );
  and2s3 U1599 ( .DIN1(RESET), .DIN2(n5597), .Q(WX5964) );
  and2s3 U1600 ( .DIN1(RESET), .DIN2(n5602), .Q(WX5962) );
  and2s3 U1601 ( .DIN1(RESET), .DIN2(n5607), .Q(WX5960) );
  and2s3 U1602 ( .DIN1(RESET), .DIN2(n5612), .Q(WX5958) );
  and2s3 U1603 ( .DIN1(RESET), .DIN2(n5617), .Q(WX5956) );
  and2s3 U1604 ( .DIN1(RESET), .DIN2(n5622), .Q(WX5954) );
  and2s3 U1605 ( .DIN1(RESET), .DIN2(n5627), .Q(WX5952) );
  and2s3 U1606 ( .DIN1(RESET), .DIN2(n5632), .Q(WX5950) );
  and2s3 U1607 ( .DIN1(RESET), .DIN2(n5637), .Q(WX5948) );
  and2s3 U1608 ( .DIN1(RESET), .DIN2(n5642), .Q(WX5946) );
  and2s3 U1609 ( .DIN1(RESET), .DIN2(n5647), .Q(WX5944) );
  and2s3 U1610 ( .DIN1(RESET), .DIN2(n5507), .Q(WX5942) );
  and2s3 U1611 ( .DIN1(RESET), .DIN2(n5511), .Q(WX5940) );
  and2s3 U1612 ( .DIN1(RESET), .DIN2(n5515), .Q(WX5938) );
  and2s3 U1613 ( .DIN1(RESET), .DIN2(n5519), .Q(WX5936) );
  and2s3 U1614 ( .DIN1(RESET), .DIN2(n5523), .Q(WX5934) );
  and2s3 U1615 ( .DIN1(RESET), .DIN2(n5527), .Q(WX5932) );
  and2s3 U1616 ( .DIN1(RESET), .DIN2(n5531), .Q(WX5930) );
  and2s3 U1617 ( .DIN1(RESET), .DIN2(n5535), .Q(WX5928) );
  and2s3 U1618 ( .DIN1(RESET), .DIN2(n5539), .Q(WX5926) );
  and2s3 U1619 ( .DIN1(RESET), .DIN2(n5543), .Q(WX5924) );
  and2s3 U1620 ( .DIN1(RESET), .DIN2(n5547), .Q(WX5922) );
  and2s3 U1621 ( .DIN1(RESET), .DIN2(n5551), .Q(WX5920) );
  and2s3 U1622 ( .DIN1(RESET), .DIN2(n5555), .Q(WX5918) );
  and2s3 U1623 ( .DIN1(RESET), .DIN2(n5559), .Q(WX5916) );
  and2s3 U1624 ( .DIN1(RESET), .DIN2(n5563), .Q(WX5914) );
  and2s3 U1625 ( .DIN1(RESET), .DIN2(n5567), .Q(WX5912) );
  nor2s3 U1626 ( .DIN1(n5571), .DIN2(n6730), .Q(WX5910) );
  nor2s3 U1627 ( .DIN1(n5576), .DIN2(n6730), .Q(WX5908) );
  nor2s3 U1628 ( .DIN1(n5581), .DIN2(n6730), .Q(WX5906) );
  nor2s3 U1629 ( .DIN1(n5586), .DIN2(n6730), .Q(WX5904) );
  nor2s3 U1630 ( .DIN1(n5591), .DIN2(n6730), .Q(WX5902) );
  nor2s3 U1631 ( .DIN1(n5596), .DIN2(n6730), .Q(WX5900) );
  nor2s3 U1632 ( .DIN1(n5601), .DIN2(n6730), .Q(WX5898) );
  nor2s3 U1633 ( .DIN1(n5606), .DIN2(n6730), .Q(WX5896) );
  nor2s3 U1634 ( .DIN1(n5611), .DIN2(n6730), .Q(WX5894) );
  nor2s3 U1635 ( .DIN1(n5616), .DIN2(n6730), .Q(WX5892) );
  nor2s3 U1636 ( .DIN1(n5621), .DIN2(n6729), .Q(WX5890) );
  nor2s3 U1637 ( .DIN1(n5626), .DIN2(n6729), .Q(WX5888) );
  nor2s3 U1638 ( .DIN1(n5631), .DIN2(n6729), .Q(WX5886) );
  nor2s3 U1639 ( .DIN1(n5636), .DIN2(n6729), .Q(WX5884) );
  nor2s3 U1640 ( .DIN1(n5641), .DIN2(n6729), .Q(WX5882) );
  nor2s3 U1641 ( .DIN1(n5646), .DIN2(n6729), .Q(WX5880) );
  nnd4s2 U1642 ( .DIN1(n3409), .DIN2(n3410), .DIN3(n3411), .DIN4(n3412), .Q(
        WX5878) );
  nnd2s3 U1643 ( .DIN1(n2820), .DIN2(n6626), .Q(n3412) );
  xor2s3 U1644 ( .DIN1(n3413), .DIN2(n3414), .Q(n2820) );
  xor2s3 U1645 ( .DIN1(n5331), .DIN2(n5332), .Q(n3414) );
  xnr2s3 U1646 ( .DIN1(n3237), .DIN2(n5333), .Q(n3413) );
  nnd2s3 U1647 ( .DIN1(n3415), .DIN2(n6659), .Q(n3411) );
  nnd2s3 U1648 ( .DIN1(n6606), .DIN2(n2017), .Q(n3410) );
  nnd2s3 U1649 ( .DIN1(n6575), .DIN2(n2016), .Q(n3409) );
  nnd4s2 U1650 ( .DIN1(n3416), .DIN2(n3417), .DIN3(n3418), .DIN4(n3419), .Q(
        WX5876) );
  nnd2s3 U1651 ( .DIN1(n2827), .DIN2(n6626), .Q(n3419) );
  xor2s3 U1652 ( .DIN1(n3420), .DIN2(n3421), .Q(n2827) );
  xor2s3 U1653 ( .DIN1(n5335), .DIN2(n5336), .Q(n3421) );
  xnr2s3 U1654 ( .DIN1(n3238), .DIN2(n5337), .Q(n3420) );
  nnd2s3 U1655 ( .DIN1(n3422), .DIN2(n6659), .Q(n3418) );
  nnd2s3 U1656 ( .DIN1(n6606), .DIN2(n2018), .Q(n3417) );
  nnd2s3 U1657 ( .DIN1(n6575), .DIN2(n2015), .Q(n3416) );
  nnd4s2 U1658 ( .DIN1(n3423), .DIN2(n3424), .DIN3(n3425), .DIN4(n3426), .Q(
        WX5874) );
  nnd2s3 U1659 ( .DIN1(n2834), .DIN2(n6626), .Q(n3426) );
  xor2s3 U1660 ( .DIN1(n3427), .DIN2(n3428), .Q(n2834) );
  xor2s3 U1661 ( .DIN1(n5339), .DIN2(n5340), .Q(n3428) );
  xnr2s3 U1662 ( .DIN1(n3239), .DIN2(n5341), .Q(n3427) );
  nnd2s3 U1663 ( .DIN1(n3429), .DIN2(n6659), .Q(n3425) );
  nnd2s3 U1664 ( .DIN1(n6606), .DIN2(n2019), .Q(n3424) );
  nnd2s3 U1665 ( .DIN1(n6575), .DIN2(n2014), .Q(n3423) );
  nnd4s2 U1666 ( .DIN1(n3430), .DIN2(n3431), .DIN3(n3432), .DIN4(n3433), .Q(
        WX5872) );
  nnd2s3 U1667 ( .DIN1(n2841), .DIN2(n6626), .Q(n3433) );
  xor2s3 U1668 ( .DIN1(n3434), .DIN2(n3435), .Q(n2841) );
  xor2s3 U1669 ( .DIN1(n5343), .DIN2(n5344), .Q(n3435) );
  xnr2s3 U1670 ( .DIN1(n3240), .DIN2(n5345), .Q(n3434) );
  nnd2s3 U1671 ( .DIN1(n3436), .DIN2(n6659), .Q(n3432) );
  nnd2s3 U1672 ( .DIN1(n6606), .DIN2(n2020), .Q(n3431) );
  nnd2s3 U1673 ( .DIN1(n6575), .DIN2(n2013), .Q(n3430) );
  nnd4s2 U1674 ( .DIN1(n3437), .DIN2(n3438), .DIN3(n3439), .DIN4(n3440), .Q(
        WX5870) );
  nnd2s3 U1675 ( .DIN1(n2848), .DIN2(n6625), .Q(n3440) );
  xor2s3 U1676 ( .DIN1(n3441), .DIN2(n3442), .Q(n2848) );
  xor2s3 U1677 ( .DIN1(n5347), .DIN2(n5348), .Q(n3442) );
  xnr2s3 U1678 ( .DIN1(n3241), .DIN2(n5349), .Q(n3441) );
  nnd2s3 U1679 ( .DIN1(n3443), .DIN2(n6659), .Q(n3439) );
  nnd2s3 U1680 ( .DIN1(n6605), .DIN2(n2021), .Q(n3438) );
  nnd2s3 U1681 ( .DIN1(n6574), .DIN2(n2012), .Q(n3437) );
  nnd4s2 U1682 ( .DIN1(n3444), .DIN2(n3445), .DIN3(n3446), .DIN4(n3447), .Q(
        WX5868) );
  nnd2s3 U1683 ( .DIN1(n2855), .DIN2(n6625), .Q(n3447) );
  xor2s3 U1684 ( .DIN1(n3448), .DIN2(n3449), .Q(n2855) );
  xor2s3 U1685 ( .DIN1(n5351), .DIN2(n5352), .Q(n3449) );
  xnr2s3 U1686 ( .DIN1(n3242), .DIN2(n5353), .Q(n3448) );
  nnd2s3 U1687 ( .DIN1(n3450), .DIN2(n6658), .Q(n3446) );
  nnd2s3 U1688 ( .DIN1(n6605), .DIN2(n2022), .Q(n3445) );
  nnd2s3 U1689 ( .DIN1(n6574), .DIN2(n2011), .Q(n3444) );
  nnd4s2 U1690 ( .DIN1(n3451), .DIN2(n3452), .DIN3(n3453), .DIN4(n3454), .Q(
        WX5866) );
  nnd2s3 U1691 ( .DIN1(n2862), .DIN2(n6625), .Q(n3454) );
  xor2s3 U1692 ( .DIN1(n3455), .DIN2(n3456), .Q(n2862) );
  xor2s3 U1693 ( .DIN1(n5355), .DIN2(n5356), .Q(n3456) );
  xnr2s3 U1694 ( .DIN1(n3243), .DIN2(n5357), .Q(n3455) );
  nnd2s3 U1695 ( .DIN1(n3457), .DIN2(n6659), .Q(n3453) );
  nnd2s3 U1696 ( .DIN1(n6605), .DIN2(n2023), .Q(n3452) );
  nnd2s3 U1697 ( .DIN1(n6574), .DIN2(n2010), .Q(n3451) );
  nnd4s2 U1698 ( .DIN1(n3458), .DIN2(n3459), .DIN3(n3460), .DIN4(n3461), .Q(
        WX5864) );
  nnd2s3 U1699 ( .DIN1(n2869), .DIN2(n6628), .Q(n3461) );
  xor2s3 U1700 ( .DIN1(n3462), .DIN2(n3463), .Q(n2869) );
  xor2s3 U1701 ( .DIN1(n5359), .DIN2(n5360), .Q(n3463) );
  xnr2s3 U1702 ( .DIN1(n3244), .DIN2(n5361), .Q(n3462) );
  nnd2s3 U1703 ( .DIN1(n3464), .DIN2(n6658), .Q(n3460) );
  nnd2s3 U1704 ( .DIN1(n6605), .DIN2(n2024), .Q(n3459) );
  nnd2s3 U1705 ( .DIN1(n6574), .DIN2(n2009), .Q(n3458) );
  nnd4s2 U1706 ( .DIN1(n3465), .DIN2(n3466), .DIN3(n3467), .DIN4(n3468), .Q(
        WX5862) );
  nnd2s3 U1707 ( .DIN1(n2876), .DIN2(n6625), .Q(n3468) );
  xor2s3 U1708 ( .DIN1(n3469), .DIN2(n3470), .Q(n2876) );
  xor2s3 U1709 ( .DIN1(n5363), .DIN2(n5364), .Q(n3470) );
  xnr2s3 U1710 ( .DIN1(n3245), .DIN2(n5365), .Q(n3469) );
  nnd2s3 U1711 ( .DIN1(n3471), .DIN2(n6661), .Q(n3467) );
  nnd2s3 U1712 ( .DIN1(n6605), .DIN2(n2025), .Q(n3466) );
  nnd2s3 U1713 ( .DIN1(n6574), .DIN2(n2008), .Q(n3465) );
  nnd4s2 U1714 ( .DIN1(n3472), .DIN2(n3473), .DIN3(n3474), .DIN4(n3475), .Q(
        WX5860) );
  nnd2s3 U1715 ( .DIN1(n2883), .DIN2(n6625), .Q(n3475) );
  xor2s3 U1716 ( .DIN1(n3476), .DIN2(n3477), .Q(n2883) );
  xor2s3 U1717 ( .DIN1(n5367), .DIN2(n5368), .Q(n3477) );
  xnr2s3 U1718 ( .DIN1(n3246), .DIN2(n5369), .Q(n3476) );
  nnd2s3 U1719 ( .DIN1(n3478), .DIN2(n6658), .Q(n3474) );
  nnd2s3 U1720 ( .DIN1(n6605), .DIN2(n2026), .Q(n3473) );
  nnd2s3 U1721 ( .DIN1(n6574), .DIN2(n2007), .Q(n3472) );
  nnd4s2 U1722 ( .DIN1(n3479), .DIN2(n3480), .DIN3(n3481), .DIN4(n3482), .Q(
        WX5858) );
  nnd2s3 U1723 ( .DIN1(n2890), .DIN2(n6625), .Q(n3482) );
  xor2s3 U1724 ( .DIN1(n3483), .DIN2(n3484), .Q(n2890) );
  xor2s3 U1725 ( .DIN1(n5371), .DIN2(n5372), .Q(n3484) );
  xnr2s3 U1726 ( .DIN1(n3247), .DIN2(n5373), .Q(n3483) );
  nnd2s3 U1727 ( .DIN1(n3485), .DIN2(n6659), .Q(n3481) );
  nnd2s3 U1728 ( .DIN1(n6605), .DIN2(n2027), .Q(n3480) );
  nnd2s3 U1729 ( .DIN1(n6574), .DIN2(n2006), .Q(n3479) );
  nnd4s2 U1730 ( .DIN1(n3486), .DIN2(n3487), .DIN3(n3488), .DIN4(n3489), .Q(
        WX5856) );
  nnd2s3 U1731 ( .DIN1(n2897), .DIN2(n6625), .Q(n3489) );
  xor2s3 U1732 ( .DIN1(n3490), .DIN2(n3491), .Q(n2897) );
  xor2s3 U1733 ( .DIN1(n5375), .DIN2(n5376), .Q(n3491) );
  xnr2s3 U1734 ( .DIN1(n3248), .DIN2(n5377), .Q(n3490) );
  nnd2s3 U1735 ( .DIN1(n3492), .DIN2(n6658), .Q(n3488) );
  nnd2s3 U1736 ( .DIN1(n6605), .DIN2(n2028), .Q(n3487) );
  nnd2s3 U1737 ( .DIN1(n6574), .DIN2(n2005), .Q(n3486) );
  nnd4s2 U1738 ( .DIN1(n3493), .DIN2(n3494), .DIN3(n3495), .DIN4(n3496), .Q(
        WX5854) );
  nnd2s3 U1739 ( .DIN1(n2904), .DIN2(n6625), .Q(n3496) );
  xor2s3 U1740 ( .DIN1(n3497), .DIN2(n3498), .Q(n2904) );
  xor2s3 U1741 ( .DIN1(n5379), .DIN2(n5380), .Q(n3498) );
  xnr2s3 U1742 ( .DIN1(n3249), .DIN2(n5381), .Q(n3497) );
  nnd2s3 U1743 ( .DIN1(n3499), .DIN2(n6659), .Q(n3495) );
  nnd2s3 U1744 ( .DIN1(n6605), .DIN2(n2029), .Q(n3494) );
  nnd2s3 U1745 ( .DIN1(n6574), .DIN2(n2004), .Q(n3493) );
  nnd4s2 U1746 ( .DIN1(n3500), .DIN2(n3501), .DIN3(n3502), .DIN4(n3503), .Q(
        WX5852) );
  nnd2s3 U1747 ( .DIN1(n2911), .DIN2(n6625), .Q(n3503) );
  xor2s3 U1748 ( .DIN1(n3504), .DIN2(n3505), .Q(n2911) );
  xor2s3 U1749 ( .DIN1(n5383), .DIN2(n5384), .Q(n3505) );
  xnr2s3 U1750 ( .DIN1(n3250), .DIN2(n5385), .Q(n3504) );
  nnd2s3 U1751 ( .DIN1(n3506), .DIN2(n6658), .Q(n3502) );
  nnd2s3 U1752 ( .DIN1(n6605), .DIN2(n2030), .Q(n3501) );
  nnd2s3 U1753 ( .DIN1(n6574), .DIN2(n2003), .Q(n3500) );
  nnd4s2 U1754 ( .DIN1(n3507), .DIN2(n3508), .DIN3(n3509), .DIN4(n3510), .Q(
        WX5850) );
  nnd2s3 U1755 ( .DIN1(n2918), .DIN2(n6625), .Q(n3510) );
  xor2s3 U1756 ( .DIN1(n3511), .DIN2(n3512), .Q(n2918) );
  xor2s3 U1757 ( .DIN1(n5387), .DIN2(n5388), .Q(n3512) );
  xnr2s3 U1758 ( .DIN1(n3251), .DIN2(n5389), .Q(n3511) );
  nnd2s3 U1759 ( .DIN1(n3513), .DIN2(n6659), .Q(n3509) );
  nnd2s3 U1760 ( .DIN1(n6605), .DIN2(n2031), .Q(n3508) );
  nnd2s3 U1761 ( .DIN1(n6574), .DIN2(n2002), .Q(n3507) );
  nnd4s2 U1762 ( .DIN1(n3514), .DIN2(n3515), .DIN3(n3516), .DIN4(n3517), .Q(
        WX5848) );
  nnd2s3 U1763 ( .DIN1(n2925), .DIN2(n6630), .Q(n3517) );
  xor2s3 U1764 ( .DIN1(n3518), .DIN2(n3519), .Q(n2925) );
  xor2s3 U1765 ( .DIN1(n5391), .DIN2(n5392), .Q(n3519) );
  xnr2s3 U1766 ( .DIN1(n3252), .DIN2(n5393), .Q(n3518) );
  nnd2s3 U1767 ( .DIN1(n3520), .DIN2(n6658), .Q(n3516) );
  nnd2s3 U1768 ( .DIN1(n6605), .DIN2(n2032), .Q(n3515) );
  nnd2s3 U1769 ( .DIN1(n6574), .DIN2(n2001), .Q(n3514) );
  nnd4s2 U1770 ( .DIN1(n3521), .DIN2(n3522), .DIN3(n3523), .DIN4(n3524), .Q(
        WX5846) );
  nnd2s3 U1771 ( .DIN1(n2933), .DIN2(n6647), .Q(n3524) );
  xor2s3 U1772 ( .DIN1(n3525), .DIN2(n3526), .Q(n2933) );
  xor2s3 U1773 ( .DIN1(n5397), .DIN2(n3527), .Q(n3526) );
  xor2s3 U1774 ( .DIN1(n5395), .DIN2(n5396), .Q(n3527) );
  xor2s3 U1775 ( .DIN1(n5398), .DIN2(n6689), .Q(n3525) );
  nnd2s3 U1776 ( .DIN1(n3528), .DIN2(n6678), .Q(n3523) );
  nnd2s3 U1777 ( .DIN1(n6605), .DIN2(n2033), .Q(n3522) );
  nnd2s3 U1778 ( .DIN1(n6574), .DIN2(n2000), .Q(n3521) );
  nnd4s2 U1779 ( .DIN1(n3529), .DIN2(n3530), .DIN3(n3531), .DIN4(n3532), .Q(
        WX5844) );
  nnd2s3 U1780 ( .DIN1(n2941), .DIN2(n6647), .Q(n3532) );
  xor2s3 U1781 ( .DIN1(n3533), .DIN2(n3534), .Q(n2941) );
  xor2s3 U1782 ( .DIN1(n5402), .DIN2(n3535), .Q(n3534) );
  xor2s3 U1783 ( .DIN1(n5400), .DIN2(n5401), .Q(n3535) );
  xor2s3 U1784 ( .DIN1(n5403), .DIN2(n6689), .Q(n3533) );
  nnd2s3 U1785 ( .DIN1(n3536), .DIN2(n6678), .Q(n3531) );
  nnd2s3 U1786 ( .DIN1(n6604), .DIN2(n2034), .Q(n3530) );
  nnd2s3 U1787 ( .DIN1(n6573), .DIN2(n1999), .Q(n3529) );
  nnd4s2 U1788 ( .DIN1(n3537), .DIN2(n3538), .DIN3(n3539), .DIN4(n3540), .Q(
        WX5842) );
  nnd2s3 U1789 ( .DIN1(n2949), .DIN2(n6646), .Q(n3540) );
  xor2s3 U1790 ( .DIN1(n3541), .DIN2(n3542), .Q(n2949) );
  xor2s3 U1791 ( .DIN1(n5407), .DIN2(n3543), .Q(n3542) );
  xor2s3 U1792 ( .DIN1(n5405), .DIN2(n5406), .Q(n3543) );
  xor2s3 U1793 ( .DIN1(n5408), .DIN2(n6689), .Q(n3541) );
  nnd2s3 U1794 ( .DIN1(n3544), .DIN2(n6677), .Q(n3539) );
  nnd2s3 U1795 ( .DIN1(n6604), .DIN2(n2035), .Q(n3538) );
  nnd2s3 U1796 ( .DIN1(n6573), .DIN2(n1998), .Q(n3537) );
  nnd4s2 U1797 ( .DIN1(n3545), .DIN2(n3546), .DIN3(n3547), .DIN4(n3548), .Q(
        WX5840) );
  nnd2s3 U1798 ( .DIN1(n2957), .DIN2(n6646), .Q(n3548) );
  xor2s3 U1799 ( .DIN1(n3549), .DIN2(n3550), .Q(n2957) );
  xor2s3 U1800 ( .DIN1(n5412), .DIN2(n3551), .Q(n3550) );
  xor2s3 U1801 ( .DIN1(n5410), .DIN2(n5411), .Q(n3551) );
  xor2s3 U1802 ( .DIN1(n5413), .DIN2(n6689), .Q(n3549) );
  nnd2s3 U1803 ( .DIN1(n3552), .DIN2(n6677), .Q(n3547) );
  nnd2s3 U1804 ( .DIN1(n6604), .DIN2(n2036), .Q(n3546) );
  nnd2s3 U1805 ( .DIN1(n6573), .DIN2(n1997), .Q(n3545) );
  nnd4s2 U1806 ( .DIN1(n3553), .DIN2(n3554), .DIN3(n3555), .DIN4(n3556), .Q(
        WX5838) );
  nnd2s3 U1807 ( .DIN1(n2965), .DIN2(n6646), .Q(n3556) );
  xor2s3 U1808 ( .DIN1(n3557), .DIN2(n3558), .Q(n2965) );
  xor2s3 U1809 ( .DIN1(n5417), .DIN2(n3559), .Q(n3558) );
  xor2s3 U1810 ( .DIN1(n5415), .DIN2(n5416), .Q(n3559) );
  xor2s3 U1811 ( .DIN1(n5418), .DIN2(n6689), .Q(n3557) );
  nnd2s3 U1812 ( .DIN1(n3560), .DIN2(n6677), .Q(n3555) );
  nnd2s3 U1813 ( .DIN1(n6604), .DIN2(n2037), .Q(n3554) );
  nnd2s3 U1814 ( .DIN1(n6573), .DIN2(n1996), .Q(n3553) );
  nnd4s2 U1815 ( .DIN1(n3561), .DIN2(n3562), .DIN3(n3563), .DIN4(n3564), .Q(
        WX5836) );
  nnd2s3 U1816 ( .DIN1(n2973), .DIN2(n6646), .Q(n3564) );
  xor2s3 U1817 ( .DIN1(n3565), .DIN2(n3566), .Q(n2973) );
  xor2s3 U1818 ( .DIN1(n5422), .DIN2(n3567), .Q(n3566) );
  xor2s3 U1819 ( .DIN1(n5420), .DIN2(n5421), .Q(n3567) );
  xor2s3 U1820 ( .DIN1(n5423), .DIN2(n6689), .Q(n3565) );
  nnd2s3 U1821 ( .DIN1(n3568), .DIN2(n6677), .Q(n3563) );
  nnd2s3 U1822 ( .DIN1(n6604), .DIN2(n2038), .Q(n3562) );
  nnd2s3 U1823 ( .DIN1(n6573), .DIN2(n1995), .Q(n3561) );
  nnd4s2 U1824 ( .DIN1(n3569), .DIN2(n3570), .DIN3(n3571), .DIN4(n3572), .Q(
        WX5834) );
  nnd2s3 U1825 ( .DIN1(n2981), .DIN2(n6646), .Q(n3572) );
  xor2s3 U1826 ( .DIN1(n3573), .DIN2(n3574), .Q(n2981) );
  xor2s3 U1827 ( .DIN1(n5427), .DIN2(n3575), .Q(n3574) );
  xor2s3 U1828 ( .DIN1(n5425), .DIN2(n5426), .Q(n3575) );
  xor2s3 U1829 ( .DIN1(n5428), .DIN2(n6689), .Q(n3573) );
  nnd2s3 U1830 ( .DIN1(n3576), .DIN2(n6677), .Q(n3571) );
  nnd2s3 U1831 ( .DIN1(n6604), .DIN2(n2039), .Q(n3570) );
  nnd2s3 U1832 ( .DIN1(n6573), .DIN2(n1994), .Q(n3569) );
  nnd4s2 U1833 ( .DIN1(n3577), .DIN2(n3578), .DIN3(n3579), .DIN4(n3580), .Q(
        WX5832) );
  nnd2s3 U1834 ( .DIN1(n2989), .DIN2(n6646), .Q(n3580) );
  xor2s3 U1835 ( .DIN1(n3581), .DIN2(n3582), .Q(n2989) );
  xor2s3 U1836 ( .DIN1(n5432), .DIN2(n3583), .Q(n3582) );
  xor2s3 U1837 ( .DIN1(n5430), .DIN2(n5431), .Q(n3583) );
  xor2s3 U1838 ( .DIN1(n5433), .DIN2(n6690), .Q(n3581) );
  nnd2s3 U1839 ( .DIN1(n3584), .DIN2(n6677), .Q(n3579) );
  nnd2s3 U1840 ( .DIN1(n6604), .DIN2(n2040), .Q(n3578) );
  nnd2s3 U1841 ( .DIN1(n6573), .DIN2(n1993), .Q(n3577) );
  nnd4s2 U1842 ( .DIN1(n3585), .DIN2(n3586), .DIN3(n3587), .DIN4(n3588), .Q(
        WX5830) );
  nnd2s3 U1843 ( .DIN1(n2997), .DIN2(n6646), .Q(n3588) );
  xor2s3 U1844 ( .DIN1(n3589), .DIN2(n3590), .Q(n2997) );
  xor2s3 U1845 ( .DIN1(n5437), .DIN2(n3591), .Q(n3590) );
  xor2s3 U1846 ( .DIN1(n5435), .DIN2(n5436), .Q(n3591) );
  xor2s3 U1847 ( .DIN1(n5438), .DIN2(n6690), .Q(n3589) );
  nnd2s3 U1848 ( .DIN1(n3592), .DIN2(n6677), .Q(n3587) );
  nnd2s3 U1849 ( .DIN1(n6604), .DIN2(n2041), .Q(n3586) );
  nnd2s3 U1850 ( .DIN1(n6573), .DIN2(n1992), .Q(n3585) );
  nnd4s2 U1851 ( .DIN1(n3593), .DIN2(n3594), .DIN3(n3595), .DIN4(n3596), .Q(
        WX5828) );
  nnd2s3 U1852 ( .DIN1(n3005), .DIN2(n6646), .Q(n3596) );
  xor2s3 U1853 ( .DIN1(n3597), .DIN2(n3598), .Q(n3005) );
  xor2s3 U1854 ( .DIN1(n5442), .DIN2(n3599), .Q(n3598) );
  xor2s3 U1855 ( .DIN1(n5440), .DIN2(n5441), .Q(n3599) );
  xor2s3 U1856 ( .DIN1(n5443), .DIN2(n6690), .Q(n3597) );
  nnd2s3 U1857 ( .DIN1(n3600), .DIN2(n6677), .Q(n3595) );
  nnd2s3 U1858 ( .DIN1(n6604), .DIN2(n2042), .Q(n3594) );
  nnd2s3 U1859 ( .DIN1(n6573), .DIN2(n1991), .Q(n3593) );
  nnd4s2 U1860 ( .DIN1(n3601), .DIN2(n3602), .DIN3(n3603), .DIN4(n3604), .Q(
        WX5826) );
  nnd2s3 U1861 ( .DIN1(n3013), .DIN2(n6646), .Q(n3604) );
  xor2s3 U1862 ( .DIN1(n3605), .DIN2(n3606), .Q(n3013) );
  xor2s3 U1863 ( .DIN1(n5447), .DIN2(n3607), .Q(n3606) );
  xor2s3 U1864 ( .DIN1(n5445), .DIN2(n5446), .Q(n3607) );
  xor2s3 U1865 ( .DIN1(n5448), .DIN2(n6690), .Q(n3605) );
  nnd2s3 U1866 ( .DIN1(n3608), .DIN2(n6677), .Q(n3603) );
  nnd2s3 U1867 ( .DIN1(n6604), .DIN2(n2043), .Q(n3602) );
  nnd2s3 U1868 ( .DIN1(n6573), .DIN2(n1990), .Q(n3601) );
  nnd4s2 U1869 ( .DIN1(n3609), .DIN2(n3610), .DIN3(n3611), .DIN4(n3612), .Q(
        WX5824) );
  nnd2s3 U1870 ( .DIN1(n3021), .DIN2(n6646), .Q(n3612) );
  xor2s3 U1871 ( .DIN1(n3613), .DIN2(n3614), .Q(n3021) );
  xor2s3 U1872 ( .DIN1(n5452), .DIN2(n3615), .Q(n3614) );
  xor2s3 U1873 ( .DIN1(n5450), .DIN2(n5451), .Q(n3615) );
  xor2s3 U1874 ( .DIN1(n5453), .DIN2(n6690), .Q(n3613) );
  nnd2s3 U1875 ( .DIN1(n3616), .DIN2(n6677), .Q(n3611) );
  nnd2s3 U1876 ( .DIN1(n6604), .DIN2(n2044), .Q(n3610) );
  nnd2s3 U1877 ( .DIN1(n6573), .DIN2(n1989), .Q(n3609) );
  nnd4s2 U1878 ( .DIN1(n3617), .DIN2(n3618), .DIN3(n3619), .DIN4(n3620), .Q(
        WX5822) );
  nnd2s3 U1879 ( .DIN1(n3029), .DIN2(n6646), .Q(n3620) );
  xor2s3 U1880 ( .DIN1(n3621), .DIN2(n3622), .Q(n3029) );
  xor2s3 U1881 ( .DIN1(n5457), .DIN2(n3623), .Q(n3622) );
  xor2s3 U1882 ( .DIN1(n5455), .DIN2(n5456), .Q(n3623) );
  xor2s3 U1883 ( .DIN1(n5458), .DIN2(n6690), .Q(n3621) );
  nnd2s3 U1884 ( .DIN1(n3624), .DIN2(n6677), .Q(n3619) );
  nnd2s3 U1885 ( .DIN1(n6604), .DIN2(n2045), .Q(n3618) );
  nnd2s3 U1886 ( .DIN1(n6573), .DIN2(n1988), .Q(n3617) );
  nnd4s2 U1887 ( .DIN1(n3625), .DIN2(n3626), .DIN3(n3627), .DIN4(n3628), .Q(
        WX5820) );
  nnd2s3 U1888 ( .DIN1(n3037), .DIN2(n6646), .Q(n3628) );
  xor2s3 U1889 ( .DIN1(n3629), .DIN2(n3630), .Q(n3037) );
  xor2s3 U1890 ( .DIN1(n5462), .DIN2(n3631), .Q(n3630) );
  xor2s3 U1891 ( .DIN1(n5460), .DIN2(n5461), .Q(n3631) );
  xor2s3 U1892 ( .DIN1(n5463), .DIN2(n6690), .Q(n3629) );
  nnd2s3 U1893 ( .DIN1(n3632), .DIN2(n6677), .Q(n3627) );
  nnd2s3 U1894 ( .DIN1(n6604), .DIN2(n2046), .Q(n3626) );
  nnd2s3 U1895 ( .DIN1(n6573), .DIN2(n1987), .Q(n3625) );
  nnd4s2 U1896 ( .DIN1(n3633), .DIN2(n3634), .DIN3(n3635), .DIN4(n3636), .Q(
        WX5818) );
  nnd2s3 U1897 ( .DIN1(n3045), .DIN2(n6646), .Q(n3636) );
  xor2s3 U1898 ( .DIN1(n3637), .DIN2(n3638), .Q(n3045) );
  xor2s3 U1899 ( .DIN1(n5467), .DIN2(n3639), .Q(n3638) );
  xor2s3 U1900 ( .DIN1(n5465), .DIN2(n5466), .Q(n3639) );
  xor2s3 U1901 ( .DIN1(n5468), .DIN2(n6690), .Q(n3637) );
  nnd2s3 U1902 ( .DIN1(n3640), .DIN2(n6677), .Q(n3635) );
  nnd2s3 U1903 ( .DIN1(n6603), .DIN2(n2047), .Q(n3634) );
  nnd2s3 U1904 ( .DIN1(n6572), .DIN2(n1986), .Q(n3633) );
  nnd4s2 U1905 ( .DIN1(n3641), .DIN2(n3642), .DIN3(n3643), .DIN4(n3644), .Q(
        WX5816) );
  nnd2s3 U1906 ( .DIN1(n3053), .DIN2(n6645), .Q(n3644) );
  xor2s3 U1907 ( .DIN1(n3645), .DIN2(n3646), .Q(n3053) );
  xor2s3 U1908 ( .DIN1(n5472), .DIN2(n3647), .Q(n3646) );
  xor2s3 U1909 ( .DIN1(n5470), .DIN2(n5471), .Q(n3647) );
  xor2s3 U1910 ( .DIN1(n5473), .DIN2(n6690), .Q(n3645) );
  nnd2s3 U1911 ( .DIN1(n3648), .DIN2(n6676), .Q(n3643) );
  nnd2s3 U1912 ( .DIN1(n6603), .DIN2(n2048), .Q(n3642) );
  nnd2s3 U1913 ( .DIN1(n6572), .DIN2(n1985), .Q(n3641) );
  nor2s3 U1914 ( .DIN1(n6805), .DIN2(n2048), .Q(WX5718) );
  nor2s3 U1915 ( .DIN1(n5476), .DIN2(n6729), .Q(WX5716) );
  nor2s3 U1916 ( .DIN1(n5477), .DIN2(n6729), .Q(WX5714) );
  nor2s3 U1917 ( .DIN1(n5478), .DIN2(n6729), .Q(WX5712) );
  nor2s3 U1918 ( .DIN1(n5479), .DIN2(n6729), .Q(WX5710) );
  nor2s3 U1919 ( .DIN1(n5480), .DIN2(n6729), .Q(WX5708) );
  nor2s3 U1920 ( .DIN1(n5481), .DIN2(n6729), .Q(WX5706) );
  nor2s3 U1921 ( .DIN1(n5482), .DIN2(n6728), .Q(WX5704) );
  nor2s3 U1922 ( .DIN1(n5483), .DIN2(n6728), .Q(WX5702) );
  nor2s3 U1923 ( .DIN1(n5484), .DIN2(n6728), .Q(WX5700) );
  nor2s3 U1924 ( .DIN1(n5485), .DIN2(n6728), .Q(WX5698) );
  nor2s3 U1925 ( .DIN1(n5486), .DIN2(n6728), .Q(WX5696) );
  nor2s3 U1926 ( .DIN1(n5487), .DIN2(n6728), .Q(WX5694) );
  nor2s3 U1927 ( .DIN1(n5488), .DIN2(n6728), .Q(WX5692) );
  nor2s3 U1928 ( .DIN1(n5489), .DIN2(n6728), .Q(WX5690) );
  nor2s3 U1929 ( .DIN1(n5490), .DIN2(n6728), .Q(WX5688) );
  nor2s3 U1930 ( .DIN1(n5491), .DIN2(n6728), .Q(WX5686) );
  nor2s3 U1931 ( .DIN1(n5492), .DIN2(n6728), .Q(WX5684) );
  nor2s3 U1932 ( .DIN1(n5493), .DIN2(n6727), .Q(WX5682) );
  nor2s3 U1933 ( .DIN1(n5494), .DIN2(n6727), .Q(WX5680) );
  nor2s3 U1934 ( .DIN1(n5495), .DIN2(n6727), .Q(WX5678) );
  nor2s3 U1935 ( .DIN1(n5496), .DIN2(n6727), .Q(WX5676) );
  nor2s3 U1936 ( .DIN1(n5497), .DIN2(n6727), .Q(WX5674) );
  nor2s3 U1937 ( .DIN1(n5498), .DIN2(n6727), .Q(WX5672) );
  nor2s3 U1938 ( .DIN1(n5499), .DIN2(n6727), .Q(WX5670) );
  nor2s3 U1939 ( .DIN1(n5500), .DIN2(n6727), .Q(WX5668) );
  nor2s3 U1940 ( .DIN1(n5501), .DIN2(n6727), .Q(WX5666) );
  nor2s3 U1941 ( .DIN1(n5502), .DIN2(n6727), .Q(WX5664) );
  nor2s3 U1942 ( .DIN1(n5503), .DIN2(n6727), .Q(WX5662) );
  nor2s3 U1943 ( .DIN1(n5504), .DIN2(n6727), .Q(WX5660) );
  nor2s3 U1944 ( .DIN1(n5505), .DIN2(n6726), .Q(WX5658) );
  nor2s3 U1945 ( .DIN1(n5506), .DIN2(n6726), .Q(WX5656) );
  nor2s3 U1946 ( .DIN1(n6790), .DIN2(n2304), .Q(WX546) );
  nor2s3 U1947 ( .DIN1(n6179), .DIN2(n6726), .Q(WX544) );
  nor2s3 U1948 ( .DIN1(n6180), .DIN2(n6726), .Q(WX542) );
  nor2s3 U1949 ( .DIN1(n6181), .DIN2(n6726), .Q(WX540) );
  nor2s3 U1950 ( .DIN1(n6182), .DIN2(n6726), .Q(WX538) );
  nor2s3 U1951 ( .DIN1(n6183), .DIN2(n6726), .Q(WX536) );
  nor2s3 U1952 ( .DIN1(n6184), .DIN2(n6726), .Q(WX534) );
  nor2s3 U1953 ( .DIN1(n6185), .DIN2(n6726), .Q(WX532) );
  nor2s3 U1954 ( .DIN1(n6186), .DIN2(n6726), .Q(WX530) );
  nor2s3 U1955 ( .DIN1(n6187), .DIN2(n6726), .Q(WX528) );
  nor2s3 U1956 ( .DIN1(n6188), .DIN2(n6726), .Q(WX526) );
  nor2s3 U1957 ( .DIN1(n6189), .DIN2(n6725), .Q(WX524) );
  nor2s3 U1958 ( .DIN1(n6190), .DIN2(n6725), .Q(WX522) );
  nor2s3 U1959 ( .DIN1(n6794), .DIN2(n3649), .Q(WX5205) );
  xor2s3 U1960 ( .DIN1(n5645), .DIN2(n5825), .Q(n3649) );
  nor2s3 U1961 ( .DIN1(n6794), .DIN2(n3650), .Q(WX5203) );
  xor2s3 U1962 ( .DIN1(n5640), .DIN2(n5820), .Q(n3650) );
  nor2s3 U1963 ( .DIN1(n6794), .DIN2(n3651), .Q(WX5201) );
  xor2s3 U1964 ( .DIN1(n5635), .DIN2(n5815), .Q(n3651) );
  nor2s3 U1965 ( .DIN1(n6191), .DIN2(n6756), .Q(WX520) );
  nor2s3 U1966 ( .DIN1(n6794), .DIN2(n3652), .Q(WX5199) );
  xor2s3 U1967 ( .DIN1(n5630), .DIN2(n5810), .Q(n3652) );
  nor2s3 U1968 ( .DIN1(n6795), .DIN2(n3653), .Q(WX5197) );
  xor2s3 U1969 ( .DIN1(n5625), .DIN2(n5805), .Q(n3653) );
  nor2s3 U1970 ( .DIN1(n6795), .DIN2(n3654), .Q(WX5195) );
  xor2s3 U1971 ( .DIN1(n5620), .DIN2(n5800), .Q(n3654) );
  nor2s3 U1972 ( .DIN1(n6788), .DIN2(n3655), .Q(WX5193) );
  xor2s3 U1973 ( .DIN1(n5615), .DIN2(n5795), .Q(n3655) );
  nor2s3 U1974 ( .DIN1(n6795), .DIN2(n3656), .Q(WX5191) );
  xor2s3 U1975 ( .DIN1(n5610), .DIN2(n5790), .Q(n3656) );
  nor2s3 U1976 ( .DIN1(n6795), .DIN2(n3657), .Q(WX5189) );
  xor2s3 U1977 ( .DIN1(n5605), .DIN2(n5785), .Q(n3657) );
  nor2s3 U1978 ( .DIN1(n6795), .DIN2(n3658), .Q(WX5187) );
  xor2s3 U1979 ( .DIN1(n5600), .DIN2(n5780), .Q(n3658) );
  nor2s3 U1980 ( .DIN1(n6795), .DIN2(n3659), .Q(WX5185) );
  xor2s3 U1981 ( .DIN1(n5595), .DIN2(n5775), .Q(n3659) );
  nor2s3 U1982 ( .DIN1(n6795), .DIN2(n3660), .Q(WX5183) );
  xor2s3 U1983 ( .DIN1(n5590), .DIN2(n5770), .Q(n3660) );
  nor2s3 U1984 ( .DIN1(n6795), .DIN2(n3661), .Q(WX5181) );
  xor2s3 U1985 ( .DIN1(n5585), .DIN2(n5765), .Q(n3661) );
  nor2s3 U1986 ( .DIN1(n6192), .DIN2(n6725), .Q(WX518) );
  nor2s3 U1987 ( .DIN1(n6791), .DIN2(n3662), .Q(WX5179) );
  xor2s3 U1988 ( .DIN1(n5580), .DIN2(n5760), .Q(n3662) );
  nor2s3 U1989 ( .DIN1(n6791), .DIN2(n3663), .Q(WX5177) );
  xor2s3 U1990 ( .DIN1(n5575), .DIN2(n5755), .Q(n3663) );
  nor2s3 U1991 ( .DIN1(n3664), .DIN2(n6725), .Q(WX5175) );
  xnr2s3 U1992 ( .DIN1(n5750), .DIN2(n3665), .Q(n3664) );
  xor2s3 U1993 ( .DIN1(n5570), .DIN2(n5650), .Q(n3665) );
  nor2s3 U1994 ( .DIN1(n6790), .DIN2(n3666), .Q(WX5173) );
  xor2s3 U1995 ( .DIN1(n5566), .DIN2(n3284), .Q(n3666) );
  nor2s3 U1996 ( .DIN1(n6790), .DIN2(n3667), .Q(WX5171) );
  xor2s3 U1997 ( .DIN1(n5562), .DIN2(n3283), .Q(n3667) );
  nor2s3 U1998 ( .DIN1(n6790), .DIN2(n3668), .Q(WX5169) );
  xor2s3 U1999 ( .DIN1(n5558), .DIN2(n3282), .Q(n3668) );
  nor2s3 U2000 ( .DIN1(n6789), .DIN2(n3669), .Q(WX5167) );
  xor2s3 U2001 ( .DIN1(n5554), .DIN2(n3281), .Q(n3669) );
  nor2s3 U2002 ( .DIN1(n3670), .DIN2(n6725), .Q(WX5165) );
  xnr2s3 U2003 ( .DIN1(n3280), .DIN2(n3671), .Q(n3670) );
  xor2s3 U2004 ( .DIN1(n5550), .DIN2(n5650), .Q(n3671) );
  nor2s3 U2005 ( .DIN1(n6789), .DIN2(n3672), .Q(WX5163) );
  xor2s3 U2006 ( .DIN1(n5546), .DIN2(n3279), .Q(n3672) );
  nor2s3 U2007 ( .DIN1(n6789), .DIN2(n3673), .Q(WX5161) );
  xor2s3 U2008 ( .DIN1(n5542), .DIN2(n3278), .Q(n3673) );
  nor2s3 U2009 ( .DIN1(n6193), .DIN2(n6725), .Q(WX516) );
  nor2s3 U2010 ( .DIN1(n6789), .DIN2(n3674), .Q(WX5159) );
  xor2s3 U2011 ( .DIN1(n5538), .DIN2(n3277), .Q(n3674) );
  nor2s3 U2012 ( .DIN1(n6791), .DIN2(n3675), .Q(WX5157) );
  xor2s3 U2013 ( .DIN1(n5534), .DIN2(n3276), .Q(n3675) );
  nor2s3 U2014 ( .DIN1(n6790), .DIN2(n3676), .Q(WX5155) );
  xor2s3 U2015 ( .DIN1(n5530), .DIN2(n3275), .Q(n3676) );
  nor2s3 U2016 ( .DIN1(n6788), .DIN2(n3677), .Q(WX5153) );
  xor2s3 U2017 ( .DIN1(n5526), .DIN2(n3274), .Q(n3677) );
  nor2s3 U2018 ( .DIN1(n3678), .DIN2(n6725), .Q(WX5151) );
  xnr2s3 U2019 ( .DIN1(n3273), .DIN2(n3679), .Q(n3678) );
  xor2s3 U2020 ( .DIN1(n5522), .DIN2(n5650), .Q(n3679) );
  nor2s3 U2021 ( .DIN1(n6788), .DIN2(n3680), .Q(WX5149) );
  xor2s3 U2022 ( .DIN1(n5518), .DIN2(n3272), .Q(n3680) );
  nor2s3 U2023 ( .DIN1(n6789), .DIN2(n3681), .Q(WX5147) );
  xor2s3 U2024 ( .DIN1(n5514), .DIN2(n3271), .Q(n3681) );
  nor2s3 U2025 ( .DIN1(n6788), .DIN2(n3682), .Q(WX5145) );
  xor2s3 U2026 ( .DIN1(n5510), .DIN2(n3270), .Q(n3682) );
  nor2s3 U2027 ( .DIN1(n6789), .DIN2(n3683), .Q(WX5143) );
  xor2s3 U2028 ( .DIN1(n5650), .DIN2(n3269), .Q(n3683) );
  nor2s3 U2029 ( .DIN1(n6194), .DIN2(n6725), .Q(WX514) );
  nor2s3 U2030 ( .DIN1(n6195), .DIN2(n6725), .Q(WX512) );
  nor2s3 U2031 ( .DIN1(n6196), .DIN2(n6725), .Q(WX510) );
  nor2s3 U2032 ( .DIN1(n6286), .DIN2(n6725), .Q(WX508) );
  nor2s3 U2033 ( .DIN1(n6342), .DIN2(n6724), .Q(WX506) );
  nor2s3 U2034 ( .DIN1(n6354), .DIN2(n6724), .Q(WX504) );
  nor2s3 U2035 ( .DIN1(n6376), .DIN2(n6724), .Q(WX502) );
  nor2s3 U2036 ( .DIN1(n6377), .DIN2(n6724), .Q(WX500) );
  nor2s3 U2037 ( .DIN1(n6378), .DIN2(n6724), .Q(WX498) );
  nor2s3 U2038 ( .DIN1(n6379), .DIN2(n6724), .Q(WX496) );
  nor2s3 U2039 ( .DIN1(n6380), .DIN2(n6724), .Q(WX494) );
  nor2s3 U2040 ( .DIN1(n6381), .DIN2(n6724), .Q(WX492) );
  nor2s3 U2041 ( .DIN1(n6382), .DIN2(n6724), .Q(WX490) );
  nor2s3 U2042 ( .DIN1(n6431), .DIN2(n6724), .Q(WX488) );
  nor2s3 U2043 ( .DIN1(n6432), .DIN2(n6724), .Q(WX486) );
  nor2s3 U2044 ( .DIN1(n6433), .DIN2(n6724), .Q(WX484) );
  nor2s3 U2045 ( .DIN1(n5685), .DIN2(n6723), .Q(WX4777) );
  nor2s3 U2046 ( .DIN1(n5689), .DIN2(n6723), .Q(WX4775) );
  nor2s3 U2047 ( .DIN1(n5693), .DIN2(n6723), .Q(WX4773) );
  nor2s3 U2048 ( .DIN1(n5697), .DIN2(n6723), .Q(WX4771) );
  nor2s3 U2049 ( .DIN1(n5701), .DIN2(n6723), .Q(WX4769) );
  nor2s3 U2050 ( .DIN1(n5705), .DIN2(n6723), .Q(WX4767) );
  nor2s3 U2051 ( .DIN1(n5709), .DIN2(n6723), .Q(WX4765) );
  nor2s3 U2052 ( .DIN1(n5713), .DIN2(n6723), .Q(WX4763) );
  nor2s3 U2053 ( .DIN1(n5717), .DIN2(n6723), .Q(WX4761) );
  nor2s3 U2054 ( .DIN1(n5721), .DIN2(n6723), .Q(WX4759) );
  nor2s3 U2055 ( .DIN1(n5725), .DIN2(n6723), .Q(WX4757) );
  nor2s3 U2056 ( .DIN1(n5729), .DIN2(n6728), .Q(WX4755) );
  nor2s3 U2057 ( .DIN1(n5733), .DIN2(n6734), .Q(WX4753) );
  nor2s3 U2058 ( .DIN1(n5737), .DIN2(n6782), .Q(WX4751) );
  nor2s3 U2059 ( .DIN1(n5741), .DIN2(n6785), .Q(WX4749) );
  nor2s3 U2060 ( .DIN1(n5745), .DIN2(n6785), .Q(WX4747) );
  nor2s3 U2061 ( .DIN1(n5749), .DIN2(n6786), .Q(WX4745) );
  nor2s3 U2062 ( .DIN1(n5754), .DIN2(n6786), .Q(WX4743) );
  nor2s3 U2063 ( .DIN1(n5759), .DIN2(n6786), .Q(WX4741) );
  nor2s3 U2064 ( .DIN1(n5764), .DIN2(n6786), .Q(WX4739) );
  nor2s3 U2065 ( .DIN1(n5769), .DIN2(n6786), .Q(WX4737) );
  nor2s3 U2066 ( .DIN1(n5774), .DIN2(n6786), .Q(WX4735) );
  nor2s3 U2067 ( .DIN1(n5779), .DIN2(n6786), .Q(WX4733) );
  nor2s3 U2068 ( .DIN1(n5784), .DIN2(n6786), .Q(WX4731) );
  nor2s3 U2069 ( .DIN1(n5789), .DIN2(n6787), .Q(WX4729) );
  nor2s3 U2070 ( .DIN1(n5794), .DIN2(n6786), .Q(WX4727) );
  nor2s3 U2071 ( .DIN1(n5799), .DIN2(n6788), .Q(WX4725) );
  nor2s3 U2072 ( .DIN1(n5804), .DIN2(n6787), .Q(WX4723) );
  nor2s3 U2073 ( .DIN1(n5809), .DIN2(n6787), .Q(WX4721) );
  nor2s3 U2074 ( .DIN1(n5814), .DIN2(n6787), .Q(WX4719) );
  nor2s3 U2075 ( .DIN1(n5819), .DIN2(n6787), .Q(WX4717) );
  nor2s3 U2076 ( .DIN1(n5824), .DIN2(n6787), .Q(WX4715) );
  nor2s3 U2077 ( .DIN1(n5684), .DIN2(n6787), .Q(WX4713) );
  nor2s3 U2078 ( .DIN1(n5688), .DIN2(n6787), .Q(WX4711) );
  nor2s3 U2079 ( .DIN1(n5692), .DIN2(n6787), .Q(WX4709) );
  nor2s3 U2080 ( .DIN1(n5696), .DIN2(n6786), .Q(WX4707) );
  nor2s3 U2081 ( .DIN1(n5700), .DIN2(n6787), .Q(WX4705) );
  nor2s3 U2082 ( .DIN1(n5704), .DIN2(n6786), .Q(WX4703) );
  nor2s3 U2083 ( .DIN1(n5708), .DIN2(n6788), .Q(WX4701) );
  nor2s3 U2084 ( .DIN1(n5712), .DIN2(n6783), .Q(WX4699) );
  nor2s3 U2085 ( .DIN1(n5716), .DIN2(n6783), .Q(WX4697) );
  nor2s3 U2086 ( .DIN1(n5720), .DIN2(n6782), .Q(WX4695) );
  nor2s3 U2087 ( .DIN1(n5724), .DIN2(n6782), .Q(WX4693) );
  nor2s3 U2088 ( .DIN1(n5728), .DIN2(n6782), .Q(WX4691) );
  nor2s3 U2089 ( .DIN1(n5732), .DIN2(n6782), .Q(WX4689) );
  nor2s3 U2090 ( .DIN1(n5736), .DIN2(n6781), .Q(WX4687) );
  nor2s3 U2091 ( .DIN1(n5740), .DIN2(n6780), .Q(WX4685) );
  nor2s3 U2092 ( .DIN1(n5744), .DIN2(n6780), .Q(WX4683) );
  and2s3 U2093 ( .DIN1(RESET), .DIN2(n5748), .Q(WX4681) );
  and2s3 U2094 ( .DIN1(RESET), .DIN2(n5753), .Q(WX4679) );
  and2s3 U2095 ( .DIN1(RESET), .DIN2(n5758), .Q(WX4677) );
  and2s3 U2096 ( .DIN1(RESET), .DIN2(n5763), .Q(WX4675) );
  and2s3 U2097 ( .DIN1(RESET), .DIN2(n5768), .Q(WX4673) );
  and2s3 U2098 ( .DIN1(RESET), .DIN2(n5773), .Q(WX4671) );
  and2s3 U2099 ( .DIN1(RESET), .DIN2(n5778), .Q(WX4669) );
  and2s3 U2100 ( .DIN1(RESET), .DIN2(n5783), .Q(WX4667) );
  and2s3 U2101 ( .DIN1(RESET), .DIN2(n5788), .Q(WX4665) );
  and2s3 U2102 ( .DIN1(RESET), .DIN2(n5793), .Q(WX4663) );
  and2s3 U2103 ( .DIN1(RESET), .DIN2(n5798), .Q(WX4661) );
  and2s3 U2104 ( .DIN1(RESET), .DIN2(n5803), .Q(WX4659) );
  and2s3 U2105 ( .DIN1(RESET), .DIN2(n5808), .Q(WX4657) );
  and2s3 U2106 ( .DIN1(RESET), .DIN2(n5813), .Q(WX4655) );
  and2s3 U2107 ( .DIN1(RESET), .DIN2(n5818), .Q(WX4653) );
  and2s3 U2108 ( .DIN1(RESET), .DIN2(n5823), .Q(WX4651) );
  and2s3 U2109 ( .DIN1(RESET), .DIN2(n5683), .Q(WX4649) );
  and2s3 U2110 ( .DIN1(RESET), .DIN2(n5687), .Q(WX4647) );
  and2s3 U2111 ( .DIN1(RESET), .DIN2(n5691), .Q(WX4645) );
  and2s3 U2112 ( .DIN1(RESET), .DIN2(n5695), .Q(WX4643) );
  and2s3 U2113 ( .DIN1(RESET), .DIN2(n5699), .Q(WX4641) );
  and2s3 U2114 ( .DIN1(RESET), .DIN2(n5703), .Q(WX4639) );
  and2s3 U2115 ( .DIN1(RESET), .DIN2(n5707), .Q(WX4637) );
  and2s3 U2116 ( .DIN1(RESET), .DIN2(n5711), .Q(WX4635) );
  and2s3 U2117 ( .DIN1(RESET), .DIN2(n5715), .Q(WX4633) );
  and2s3 U2118 ( .DIN1(RESET), .DIN2(n5719), .Q(WX4631) );
  and2s3 U2119 ( .DIN1(RESET), .DIN2(n5723), .Q(WX4629) );
  and2s3 U2120 ( .DIN1(RESET), .DIN2(n5727), .Q(WX4627) );
  and2s3 U2121 ( .DIN1(RESET), .DIN2(n5731), .Q(WX4625) );
  and2s3 U2122 ( .DIN1(RESET), .DIN2(n5735), .Q(WX4623) );
  and2s3 U2123 ( .DIN1(RESET), .DIN2(n5739), .Q(WX4621) );
  and2s3 U2124 ( .DIN1(RESET), .DIN2(n5743), .Q(WX4619) );
  nor2s3 U2125 ( .DIN1(n5747), .DIN2(n6780), .Q(WX4617) );
  nor2s3 U2126 ( .DIN1(n5752), .DIN2(n6779), .Q(WX4615) );
  nor2s3 U2127 ( .DIN1(n5757), .DIN2(n6779), .Q(WX4613) );
  nor2s3 U2128 ( .DIN1(n5762), .DIN2(n6779), .Q(WX4611) );
  nor2s3 U2129 ( .DIN1(n5767), .DIN2(n6778), .Q(WX4609) );
  nor2s3 U2130 ( .DIN1(n5772), .DIN2(n6778), .Q(WX4607) );
  nor2s3 U2131 ( .DIN1(n5777), .DIN2(n6778), .Q(WX4605) );
  nor2s3 U2132 ( .DIN1(n5782), .DIN2(n6778), .Q(WX4603) );
  nor2s3 U2133 ( .DIN1(n5787), .DIN2(n6778), .Q(WX4601) );
  nor2s3 U2134 ( .DIN1(n5792), .DIN2(n6778), .Q(WX4599) );
  nor2s3 U2135 ( .DIN1(n5797), .DIN2(n6778), .Q(WX4597) );
  nor2s3 U2136 ( .DIN1(n5802), .DIN2(n6778), .Q(WX4595) );
  nor2s3 U2137 ( .DIN1(n5807), .DIN2(n6778), .Q(WX4593) );
  nor2s3 U2138 ( .DIN1(n5812), .DIN2(n6777), .Q(WX4591) );
  nor2s3 U2139 ( .DIN1(n5817), .DIN2(n6777), .Q(WX4589) );
  nor2s3 U2140 ( .DIN1(n5822), .DIN2(n6777), .Q(WX4587) );
  nnd4s2 U2141 ( .DIN1(n3684), .DIN2(n3685), .DIN3(n3686), .DIN4(n3687), .Q(
        WX4585) );
  nnd2s3 U2142 ( .DIN1(n3415), .DIN2(n6645), .Q(n3687) );
  xor2s3 U2143 ( .DIN1(n3688), .DIN2(n3689), .Q(n3415) );
  xor2s3 U2144 ( .DIN1(n5507), .DIN2(n5508), .Q(n3689) );
  xnr2s3 U2145 ( .DIN1(n3253), .DIN2(n5509), .Q(n3688) );
  nnd2s3 U2146 ( .DIN1(n3690), .DIN2(n6676), .Q(n3686) );
  nnd2s3 U2147 ( .DIN1(n6603), .DIN2(n2081), .Q(n3685) );
  nnd2s3 U2148 ( .DIN1(n6572), .DIN2(n2080), .Q(n3684) );
  nnd4s2 U2149 ( .DIN1(n3691), .DIN2(n3692), .DIN3(n3693), .DIN4(n3694), .Q(
        WX4583) );
  nnd2s3 U2150 ( .DIN1(n3422), .DIN2(n6645), .Q(n3694) );
  xor2s3 U2151 ( .DIN1(n3695), .DIN2(n3696), .Q(n3422) );
  xor2s3 U2152 ( .DIN1(n5511), .DIN2(n5512), .Q(n3696) );
  xnr2s3 U2153 ( .DIN1(n3254), .DIN2(n5513), .Q(n3695) );
  nnd2s3 U2154 ( .DIN1(n3697), .DIN2(n6676), .Q(n3693) );
  nnd2s3 U2155 ( .DIN1(n6603), .DIN2(n2082), .Q(n3692) );
  nnd2s3 U2156 ( .DIN1(n6572), .DIN2(n2079), .Q(n3691) );
  nnd4s2 U2157 ( .DIN1(n3698), .DIN2(n3699), .DIN3(n3700), .DIN4(n3701), .Q(
        WX4581) );
  nnd2s3 U2158 ( .DIN1(n3429), .DIN2(n6645), .Q(n3701) );
  xor2s3 U2159 ( .DIN1(n3702), .DIN2(n3703), .Q(n3429) );
  xor2s3 U2160 ( .DIN1(n5515), .DIN2(n5516), .Q(n3703) );
  xnr2s3 U2161 ( .DIN1(n3255), .DIN2(n5517), .Q(n3702) );
  nnd2s3 U2162 ( .DIN1(n3704), .DIN2(n6676), .Q(n3700) );
  nnd2s3 U2163 ( .DIN1(n6603), .DIN2(n2083), .Q(n3699) );
  nnd2s3 U2164 ( .DIN1(n6572), .DIN2(n2078), .Q(n3698) );
  nnd4s2 U2165 ( .DIN1(n3705), .DIN2(n3706), .DIN3(n3707), .DIN4(n3708), .Q(
        WX4579) );
  nnd2s3 U2166 ( .DIN1(n3436), .DIN2(n6645), .Q(n3708) );
  xor2s3 U2167 ( .DIN1(n3709), .DIN2(n3710), .Q(n3436) );
  xor2s3 U2168 ( .DIN1(n5519), .DIN2(n5520), .Q(n3710) );
  xnr2s3 U2169 ( .DIN1(n3256), .DIN2(n5521), .Q(n3709) );
  nnd2s3 U2170 ( .DIN1(n3711), .DIN2(n6676), .Q(n3707) );
  nnd2s3 U2171 ( .DIN1(n6603), .DIN2(n2084), .Q(n3706) );
  nnd2s3 U2172 ( .DIN1(n6572), .DIN2(n2077), .Q(n3705) );
  nnd4s2 U2173 ( .DIN1(n3712), .DIN2(n3713), .DIN3(n3714), .DIN4(n3715), .Q(
        WX4577) );
  nnd2s3 U2174 ( .DIN1(n3443), .DIN2(n6645), .Q(n3715) );
  xor2s3 U2175 ( .DIN1(n3716), .DIN2(n3717), .Q(n3443) );
  xor2s3 U2176 ( .DIN1(n5523), .DIN2(n5524), .Q(n3717) );
  xnr2s3 U2177 ( .DIN1(n3257), .DIN2(n5525), .Q(n3716) );
  nnd2s3 U2178 ( .DIN1(n3718), .DIN2(n6676), .Q(n3714) );
  nnd2s3 U2179 ( .DIN1(n6603), .DIN2(n2085), .Q(n3713) );
  nnd2s3 U2180 ( .DIN1(n6572), .DIN2(n2076), .Q(n3712) );
  nnd4s2 U2181 ( .DIN1(n3719), .DIN2(n3720), .DIN3(n3721), .DIN4(n3722), .Q(
        WX4575) );
  nnd2s3 U2182 ( .DIN1(n3450), .DIN2(n6645), .Q(n3722) );
  xor2s3 U2183 ( .DIN1(n3723), .DIN2(n3724), .Q(n3450) );
  xor2s3 U2184 ( .DIN1(n5527), .DIN2(n5528), .Q(n3724) );
  xnr2s3 U2185 ( .DIN1(n3258), .DIN2(n5529), .Q(n3723) );
  nnd2s3 U2186 ( .DIN1(n3725), .DIN2(n6676), .Q(n3721) );
  nnd2s3 U2187 ( .DIN1(n6603), .DIN2(n2086), .Q(n3720) );
  nnd2s3 U2188 ( .DIN1(n6572), .DIN2(n2075), .Q(n3719) );
  nnd4s2 U2189 ( .DIN1(n3726), .DIN2(n3727), .DIN3(n3728), .DIN4(n3729), .Q(
        WX4573) );
  nnd2s3 U2190 ( .DIN1(n3457), .DIN2(n6645), .Q(n3729) );
  xor2s3 U2191 ( .DIN1(n3730), .DIN2(n3731), .Q(n3457) );
  xor2s3 U2192 ( .DIN1(n5531), .DIN2(n5532), .Q(n3731) );
  xnr2s3 U2193 ( .DIN1(n3259), .DIN2(n5533), .Q(n3730) );
  nnd2s3 U2194 ( .DIN1(n3732), .DIN2(n6676), .Q(n3728) );
  nnd2s3 U2195 ( .DIN1(n6603), .DIN2(n2087), .Q(n3727) );
  nnd2s3 U2196 ( .DIN1(n6572), .DIN2(n2074), .Q(n3726) );
  nnd4s2 U2197 ( .DIN1(n3733), .DIN2(n3734), .DIN3(n3735), .DIN4(n3736), .Q(
        WX4571) );
  nnd2s3 U2198 ( .DIN1(n3464), .DIN2(n6645), .Q(n3736) );
  xor2s3 U2199 ( .DIN1(n3737), .DIN2(n3738), .Q(n3464) );
  xor2s3 U2200 ( .DIN1(n5535), .DIN2(n5536), .Q(n3738) );
  xnr2s3 U2201 ( .DIN1(n3260), .DIN2(n5537), .Q(n3737) );
  nnd2s3 U2202 ( .DIN1(n3739), .DIN2(n6676), .Q(n3735) );
  nnd2s3 U2203 ( .DIN1(n6603), .DIN2(n2088), .Q(n3734) );
  nnd2s3 U2204 ( .DIN1(n6572), .DIN2(n2073), .Q(n3733) );
  nnd4s2 U2205 ( .DIN1(n3740), .DIN2(n3741), .DIN3(n3742), .DIN4(n3743), .Q(
        WX4569) );
  nnd2s3 U2206 ( .DIN1(n3471), .DIN2(n6645), .Q(n3743) );
  xor2s3 U2207 ( .DIN1(n3744), .DIN2(n3745), .Q(n3471) );
  xor2s3 U2208 ( .DIN1(n5539), .DIN2(n5540), .Q(n3745) );
  xnr2s3 U2209 ( .DIN1(n3261), .DIN2(n5541), .Q(n3744) );
  nnd2s3 U2210 ( .DIN1(n3746), .DIN2(n6676), .Q(n3742) );
  nnd2s3 U2211 ( .DIN1(n6603), .DIN2(n2089), .Q(n3741) );
  nnd2s3 U2212 ( .DIN1(n6572), .DIN2(n2072), .Q(n3740) );
  nnd4s2 U2213 ( .DIN1(n3747), .DIN2(n3748), .DIN3(n3749), .DIN4(n3750), .Q(
tempWX4567) );
  nnd2s3 U2214 ( .DIN1(n3478), .DIN2(n6645), .Q(n3750) );
  xor2s3 U2215 ( .DIN1(n3751), .DIN2(n3752), .Q(n3478) );
  xor2s3 U2216 ( .DIN1(n5543), .DIN2(n5544), .Q(n3752) );
  xnr2s3 U2217 ( .DIN1(n3262), .DIN2(n5545), .Q(n3751) );
  nnd2s3 U2218 ( .DIN1(n3753), .DIN2(n6676), .Q(n3749) );
  nnd2s3 U2219 ( .DIN1(n6603), .DIN2(n2090), .Q(n3748) );
  nnd2s3 U2220 ( .DIN1(n6572), .DIN2(n2071), .Q(n3747) );
  nnd4s2 U2221 ( .DIN1(n3754), .DIN2(n3755), .DIN3(n3756), .DIN4(n3757), .Q(
        WX4565) );
  nnd2s3 U2222 ( .DIN1(n3485), .DIN2(n6645), .Q(n3757) );
  xor2s3 U2223 ( .DIN1(n3758), .DIN2(n3759), .Q(n3485) );
  xor2s3 U2224 ( .DIN1(n5547), .DIN2(n5548), .Q(n3759) );
  xnr2s3 U2225 ( .DIN1(n3263), .DIN2(n5549), .Q(n3758) );
  nnd2s3 U2226 ( .DIN1(n3760), .DIN2(n6676), .Q(n3756) );
  nnd2s3 U2227 ( .DIN1(n6603), .DIN2(n2091), .Q(n3755) );
  nnd2s3 U2228 ( .DIN1(n6572), .DIN2(n2070), .Q(n3754) );
  nnd4s2 U2229 ( .DIN1(n3761), .DIN2(n3762), .DIN3(n3763), .DIN4(n3764), .Q(
        WX4563) );
  nnd2s3 U2230 ( .DIN1(n3492), .DIN2(n6645), .Q(n3764) );
  xor2s3 U2231 ( .DIN1(n3765), .DIN2(n3766), .Q(n3492) );
  xor2s3 U2232 ( .DIN1(n5551), .DIN2(n5552), .Q(n3766) );
  xnr2s3 U2233 ( .DIN1(n3264), .DIN2(n5553), .Q(n3765) );
  nnd2s3 U2234 ( .DIN1(n3767), .DIN2(n6676), .Q(n3763) );
  nnd2s3 U2235 ( .DIN1(n6602), .DIN2(n2092), .Q(n3762) );
  nnd2s3 U2236 ( .DIN1(n6571), .DIN2(n2069), .Q(n3761) );
  nnd4s2 U2237 ( .DIN1(n3768), .DIN2(n3769), .DIN3(n3770), .DIN4(n3771), .Q(
        WX4561) );
  nnd2s3 U2238 ( .DIN1(n3499), .DIN2(n6644), .Q(n3771) );
  xor2s3 U2239 ( .DIN1(n3772), .DIN2(n3773), .Q(n3499) );
  xor2s3 U2240 ( .DIN1(n5555), .DIN2(n5556), .Q(n3773) );
  xnr2s3 U2241 ( .DIN1(n3265), .DIN2(n5557), .Q(n3772) );
  nnd2s3 U2242 ( .DIN1(n3774), .DIN2(n6675), .Q(n3770) );
  nnd2s3 U2243 ( .DIN1(n6602), .DIN2(n2093), .Q(n3769) );
  nnd2s3 U2244 ( .DIN1(n6571), .DIN2(n2068), .Q(n3768) );
  nnd4s2 U2245 ( .DIN1(n3775), .DIN2(n3776), .DIN3(n3777), .DIN4(n3778), .Q(
        WX4559) );
  nnd2s3 U2246 ( .DIN1(n3506), .DIN2(n6644), .Q(n3778) );
  xor2s3 U2247 ( .DIN1(n3779), .DIN2(n3780), .Q(n3506) );
  xor2s3 U2248 ( .DIN1(n5559), .DIN2(n5560), .Q(n3780) );
  xnr2s3 U2249 ( .DIN1(n3266), .DIN2(n5561), .Q(n3779) );
  nnd2s3 U2250 ( .DIN1(n3781), .DIN2(n6675), .Q(n3777) );
  nnd2s3 U2251 ( .DIN1(n6602), .DIN2(n2094), .Q(n3776) );
  nnd2s3 U2252 ( .DIN1(n6571), .DIN2(n2067), .Q(n3775) );
  nnd4s2 U2253 ( .DIN1(n3782), .DIN2(n3783), .DIN3(n3784), .DIN4(n3785), .Q(
        WX4557) );
  nnd2s3 U2254 ( .DIN1(n3513), .DIN2(n6644), .Q(n3785) );
  xor2s3 U2255 ( .DIN1(n3786), .DIN2(n3787), .Q(n3513) );
  xor2s3 U2256 ( .DIN1(n5563), .DIN2(n5564), .Q(n3787) );
  xnr2s3 U2257 ( .DIN1(n3267), .DIN2(n5565), .Q(n3786) );
  nnd2s3 U2258 ( .DIN1(n3788), .DIN2(n6675), .Q(n3784) );
  nnd2s3 U2259 ( .DIN1(n6602), .DIN2(n2095), .Q(n3783) );
  nnd2s3 U2260 ( .DIN1(n6571), .DIN2(n2066), .Q(n3782) );
  nnd4s2 U2261 ( .DIN1(n3789), .DIN2(n3790), .DIN3(n3791), .DIN4(n3792), .Q(
        WX4555) );
  nnd2s3 U2262 ( .DIN1(n3520), .DIN2(n6644), .Q(n3792) );
  xor2s3 U2263 ( .DIN1(n3793), .DIN2(n3794), .Q(n3520) );
  xor2s3 U2264 ( .DIN1(n5567), .DIN2(n5568), .Q(n3794) );
  xnr2s3 U2265 ( .DIN1(n3268), .DIN2(n5569), .Q(n3793) );
  nnd2s3 U2266 ( .DIN1(n3795), .DIN2(n6675), .Q(n3791) );
  nnd2s3 U2267 ( .DIN1(n6602), .DIN2(n2096), .Q(n3790) );
  nnd2s3 U2268 ( .DIN1(n6571), .DIN2(n2065), .Q(n3789) );
  nnd4s2 U2269 ( .DIN1(n3796), .DIN2(n3797), .DIN3(n3798), .DIN4(n3799), .Q(
        WX4553) );
  nnd2s3 U2270 ( .DIN1(n3528), .DIN2(n6644), .Q(n3799) );
  xor2s3 U2271 ( .DIN1(n3800), .DIN2(n3801), .Q(n3528) );
  xor2s3 U2272 ( .DIN1(n5573), .DIN2(n3802), .Q(n3801) );
  xor2s3 U2273 ( .DIN1(n5571), .DIN2(n5572), .Q(n3802) );
  xor2s3 U2274 ( .DIN1(n5574), .DIN2(n6690), .Q(n3800) );
  nnd2s3 U2275 ( .DIN1(n3803), .DIN2(n6675), .Q(n3798) );
  nnd2s3 U2276 ( .DIN1(n6602), .DIN2(n2097), .Q(n3797) );
  nnd2s3 U2277 ( .DIN1(n6571), .DIN2(n2064), .Q(n3796) );
  nnd4s2 U2278 ( .DIN1(n3804), .DIN2(n3805), .DIN3(n3806), .DIN4(n3807), .Q(
        WX4551) );
  nnd2s3 U2279 ( .DIN1(n3536), .DIN2(n6644), .Q(n3807) );
  xor2s3 U2280 ( .DIN1(n3808), .DIN2(n3809), .Q(n3536) );
  xor2s3 U2281 ( .DIN1(n5578), .DIN2(n3810), .Q(n3809) );
  xor2s3 U2282 ( .DIN1(n5576), .DIN2(n5577), .Q(n3810) );
  xor2s3 U2283 ( .DIN1(n5579), .DIN2(n6690), .Q(n3808) );
  nnd2s3 U2284 ( .DIN1(n3811), .DIN2(n6675), .Q(n3806) );
  nnd2s3 U2285 ( .DIN1(n6602), .DIN2(n2098), .Q(n3805) );
  nnd2s3 U2286 ( .DIN1(n6571), .DIN2(n2063), .Q(n3804) );
  nnd4s2 U2287 ( .DIN1(n3812), .DIN2(n3813), .DIN3(n3814), .DIN4(n3815), .Q(
        WX4549) );
  nnd2s3 U2288 ( .DIN1(n3544), .DIN2(n6644), .Q(n3815) );
  xor2s3 U2289 ( .DIN1(n3816), .DIN2(n3817), .Q(n3544) );
  xor2s3 U2290 ( .DIN1(n5583), .DIN2(n3818), .Q(n3817) );
  xor2s3 U2291 ( .DIN1(n5581), .DIN2(n5582), .Q(n3818) );
  xor2s3 U2292 ( .DIN1(n5584), .DIN2(n6690), .Q(n3816) );
  nnd2s3 U2293 ( .DIN1(n3819), .DIN2(n6675), .Q(n3814) );
  nnd2s3 U2294 ( .DIN1(n6602), .DIN2(n2099), .Q(n3813) );
  nnd2s3 U2295 ( .DIN1(n6571), .DIN2(n2062), .Q(n3812) );
  nnd4s2 U2296 ( .DIN1(n3820), .DIN2(n3821), .DIN3(n3822), .DIN4(n3823), .Q(
        WX4547) );
  nnd2s3 U2297 ( .DIN1(n3552), .DIN2(n6644), .Q(n3823) );
  xor2s3 U2298 ( .DIN1(n3824), .DIN2(n3825), .Q(n3552) );
  xor2s3 U2299 ( .DIN1(n5588), .DIN2(n3826), .Q(n3825) );
  xor2s3 U2300 ( .DIN1(n5586), .DIN2(n5587), .Q(n3826) );
  xor2s3 U2301 ( .DIN1(n5589), .DIN2(n6690), .Q(n3824) );
  nnd2s3 U2302 ( .DIN1(n3827), .DIN2(n6675), .Q(n3822) );
  nnd2s3 U2303 ( .DIN1(n6602), .DIN2(n2100), .Q(n3821) );
  nnd2s3 U2304 ( .DIN1(n6571), .DIN2(n2061), .Q(n3820) );
  nnd4s2 U2305 ( .DIN1(n3828), .DIN2(n3829), .DIN3(n3830), .DIN4(n3831), .Q(
        WX4545) );
  nnd2s3 U2306 ( .DIN1(n3560), .DIN2(n6644), .Q(n3831) );
  xor2s3 U2307 ( .DIN1(n3832), .DIN2(n3833), .Q(n3560) );
  xor2s3 U2308 ( .DIN1(n5593), .DIN2(n3834), .Q(n3833) );
  xor2s3 U2309 ( .DIN1(n5591), .DIN2(n5592), .Q(n3834) );
  xor2s3 U2310 ( .DIN1(n5594), .DIN2(n6691), .Q(n3832) );
  nnd2s3 U2311 ( .DIN1(n3835), .DIN2(n6675), .Q(n3830) );
  nnd2s3 U2312 ( .DIN1(n6602), .DIN2(n2101), .Q(n3829) );
  nnd2s3 U2313 ( .DIN1(n6571), .DIN2(n2060), .Q(n3828) );
  nnd4s2 U2314 ( .DIN1(n3836), .DIN2(n3837), .DIN3(n3838), .DIN4(n3839), .Q(
        WX4543) );
  nnd2s3 U2315 ( .DIN1(n3568), .DIN2(n6644), .Q(n3839) );
  xor2s3 U2316 ( .DIN1(n3840), .DIN2(n3841), .Q(n3568) );
  xor2s3 U2317 ( .DIN1(n5598), .DIN2(n3842), .Q(n3841) );
  xor2s3 U2318 ( .DIN1(n5596), .DIN2(n5597), .Q(n3842) );
  xor2s3 U2319 ( .DIN1(n5599), .DIN2(n6691), .Q(n3840) );
  nnd2s3 U2320 ( .DIN1(n3843), .DIN2(n6675), .Q(n3838) );
  nnd2s3 U2321 ( .DIN1(n6602), .DIN2(n2102), .Q(n3837) );
  nnd2s3 U2322 ( .DIN1(n6571), .DIN2(n2059), .Q(n3836) );
  nnd4s2 U2323 ( .DIN1(n3844), .DIN2(n3845), .DIN3(n3846), .DIN4(n3847), .Q(
        WX4541) );
  nnd2s3 U2324 ( .DIN1(n3576), .DIN2(n6644), .Q(n3847) );
  xor2s3 U2325 ( .DIN1(n3848), .DIN2(n3849), .Q(n3576) );
  xor2s3 U2326 ( .DIN1(n5603), .DIN2(n3850), .Q(n3849) );
  xor2s3 U2327 ( .DIN1(n5601), .DIN2(n5602), .Q(n3850) );
  xor2s3 U2328 ( .DIN1(n5604), .DIN2(n6691), .Q(n3848) );
  nnd2s3 U2329 ( .DIN1(n3851), .DIN2(n6675), .Q(n3846) );
  nnd2s3 U2330 ( .DIN1(n6602), .DIN2(n2103), .Q(n3845) );
  nnd2s3 U2331 ( .DIN1(n6571), .DIN2(n2058), .Q(n3844) );
  nnd4s2 U2332 ( .DIN1(n3852), .DIN2(n3853), .DIN3(n3854), .DIN4(n3855), .Q(
        WX4539) );
  nnd2s3 U2333 ( .DIN1(n3584), .DIN2(n6644), .Q(n3855) );
  xor2s3 U2334 ( .DIN1(n3856), .DIN2(n3857), .Q(n3584) );
  xor2s3 U2335 ( .DIN1(n5608), .DIN2(n3858), .Q(n3857) );
  xor2s3 U2336 ( .DIN1(n5606), .DIN2(n5607), .Q(n3858) );
  xor2s3 U2337 ( .DIN1(n5609), .DIN2(n6691), .Q(n3856) );
  nnd2s3 U2338 ( .DIN1(n3859), .DIN2(n6675), .Q(n3854) );
  nnd2s3 U2339 ( .DIN1(n6602), .DIN2(n2104), .Q(n3853) );
  nnd2s3 U2340 ( .DIN1(n6571), .DIN2(n2057), .Q(n3852) );
  nnd4s2 U2341 ( .DIN1(n3860), .DIN2(n3861), .DIN3(n3862), .DIN4(n3863), .Q(
        WX4537) );
  nnd2s3 U2342 ( .DIN1(n3592), .DIN2(n6644), .Q(n3863) );
  xor2s3 U2343 ( .DIN1(n3864), .DIN2(n3865), .Q(n3592) );
  xor2s3 U2344 ( .DIN1(n5613), .DIN2(n3866), .Q(n3865) );
  xor2s3 U2345 ( .DIN1(n5611), .DIN2(n5612), .Q(n3866) );
  xor2s3 U2346 ( .DIN1(n5614), .DIN2(n6691), .Q(n3864) );
  nnd2s3 U2347 ( .DIN1(n3867), .DIN2(n6675), .Q(n3862) );
  nnd2s3 U2348 ( .DIN1(n6601), .DIN2(n2105), .Q(n3861) );
  nnd2s3 U2349 ( .DIN1(n6570), .DIN2(n2056), .Q(n3860) );
  nnd4s2 U2350 ( .DIN1(n3868), .DIN2(n3869), .DIN3(n3870), .DIN4(n3871), .Q(
        WX4535) );
  nnd2s3 U2351 ( .DIN1(n3600), .DIN2(n6643), .Q(n3871) );
  xor2s3 U2352 ( .DIN1(n3872), .DIN2(n3873), .Q(n3600) );
  xor2s3 U2353 ( .DIN1(n5618), .DIN2(n3874), .Q(n3873) );
  xor2s3 U2354 ( .DIN1(n5616), .DIN2(n5617), .Q(n3874) );
  xor2s3 U2355 ( .DIN1(n5619), .DIN2(n6691), .Q(n3872) );
  nnd2s3 U2356 ( .DIN1(n3875), .DIN2(n6674), .Q(n3870) );
  nnd2s3 U2357 ( .DIN1(n6601), .DIN2(n2106), .Q(n3869) );
  nnd2s3 U2358 ( .DIN1(n6570), .DIN2(n2055), .Q(n3868) );
  nnd4s2 U2359 ( .DIN1(n3876), .DIN2(n3877), .DIN3(n3878), .DIN4(n3879), .Q(
        WX4533) );
  nnd2s3 U2360 ( .DIN1(n3608), .DIN2(n6643), .Q(n3879) );
  xor2s3 U2361 ( .DIN1(n3880), .DIN2(n3881), .Q(n3608) );
  xor2s3 U2362 ( .DIN1(n5623), .DIN2(n3882), .Q(n3881) );
  xor2s3 U2363 ( .DIN1(n5621), .DIN2(n5622), .Q(n3882) );
  xor2s3 U2364 ( .DIN1(n5624), .DIN2(n6691), .Q(n3880) );
  nnd2s3 U2365 ( .DIN1(n3883), .DIN2(n6674), .Q(n3878) );
  nnd2s3 U2366 ( .DIN1(n6601), .DIN2(n2107), .Q(n3877) );
  nnd2s3 U2367 ( .DIN1(n6570), .DIN2(n2054), .Q(n3876) );
  nnd4s2 U2368 ( .DIN1(n3884), .DIN2(n3885), .DIN3(n3886), .DIN4(n3887), .Q(
        WX4531) );
  nnd2s3 U2369 ( .DIN1(n3616), .DIN2(n6643), .Q(n3887) );
  xor2s3 U2370 ( .DIN1(n3888), .DIN2(n3889), .Q(n3616) );
  xor2s3 U2371 ( .DIN1(n5628), .DIN2(n3890), .Q(n3889) );
  xor2s3 U2372 ( .DIN1(n5626), .DIN2(n5627), .Q(n3890) );
  xor2s3 U2373 ( .DIN1(n5629), .DIN2(n6691), .Q(n3888) );
  nnd2s3 U2374 ( .DIN1(n3891), .DIN2(n6674), .Q(n3886) );
  nnd2s3 U2375 ( .DIN1(n6601), .DIN2(n2108), .Q(n3885) );
  nnd2s3 U2376 ( .DIN1(n6570), .DIN2(n2053), .Q(n3884) );
  nnd4s2 U2377 ( .DIN1(n3892), .DIN2(n3893), .DIN3(n3894), .DIN4(n3895), .Q(
        WX4529) );
  nnd2s3 U2378 ( .DIN1(n3624), .DIN2(n6643), .Q(n3895) );
  xor2s3 U2379 ( .DIN1(n3896), .DIN2(n3897), .Q(n3624) );
  xor2s3 U2380 ( .DIN1(n5633), .DIN2(n3898), .Q(n3897) );
  xor2s3 U2381 ( .DIN1(n5631), .DIN2(n5632), .Q(n3898) );
  xor2s3 U2382 ( .DIN1(n5634), .DIN2(n6691), .Q(n3896) );
  nnd2s3 U2383 ( .DIN1(n3899), .DIN2(n6674), .Q(n3894) );
  nnd2s3 U2384 ( .DIN1(n6601), .DIN2(n2109), .Q(n3893) );
  nnd2s3 U2385 ( .DIN1(n6570), .DIN2(n2052), .Q(n3892) );
  nnd4s2 U2386 ( .DIN1(n3900), .DIN2(n3901), .DIN3(n3902), .DIN4(n3903), .Q(
        WX4527) );
  nnd2s3 U2387 ( .DIN1(n3632), .DIN2(n6643), .Q(n3903) );
  xor2s3 U2388 ( .DIN1(n3904), .DIN2(n3905), .Q(n3632) );
  xor2s3 U2389 ( .DIN1(n5638), .DIN2(n3906), .Q(n3905) );
  xor2s3 U2390 ( .DIN1(n5636), .DIN2(n5637), .Q(n3906) );
  xor2s3 U2391 ( .DIN1(n5639), .DIN2(n6691), .Q(n3904) );
  nnd2s3 U2392 ( .DIN1(n3907), .DIN2(n6674), .Q(n3902) );
  nnd2s3 U2393 ( .DIN1(n6601), .DIN2(n2110), .Q(n3901) );
  nnd2s3 U2394 ( .DIN1(n6570), .DIN2(n2051), .Q(n3900) );
  nnd4s2 U2395 ( .DIN1(n3908), .DIN2(n3909), .DIN3(n3910), .DIN4(n3911), .Q(
        WX4525) );
  nnd2s3 U2396 ( .DIN1(n3640), .DIN2(n6643), .Q(n3911) );
  xor2s3 U2397 ( .DIN1(n3912), .DIN2(n3913), .Q(n3640) );
  xor2s3 U2398 ( .DIN1(n5643), .DIN2(n3914), .Q(n3913) );
  xor2s3 U2399 ( .DIN1(n5641), .DIN2(n5642), .Q(n3914) );
  xor2s3 U2400 ( .DIN1(n5644), .DIN2(n6691), .Q(n3912) );
  nnd2s3 U2401 ( .DIN1(n3915), .DIN2(n6674), .Q(n3910) );
  nnd2s3 U2402 ( .DIN1(n6601), .DIN2(n2111), .Q(n3909) );
  nnd2s3 U2403 ( .DIN1(n6570), .DIN2(n2050), .Q(n3908) );
  nnd4s2 U2404 ( .DIN1(n3916), .DIN2(n3917), .DIN3(n3918), .DIN4(n3919), .Q(
        WX4523) );
  nnd2s3 U2405 ( .DIN1(n3648), .DIN2(n6643), .Q(n3919) );
  xor2s3 U2406 ( .DIN1(n3920), .DIN2(n3921), .Q(n3648) );
  xor2s3 U2407 ( .DIN1(n5648), .DIN2(n3922), .Q(n3921) );
  xor2s3 U2408 ( .DIN1(n5646), .DIN2(n5647), .Q(n3922) );
  xor2s3 U2409 ( .DIN1(n5649), .DIN2(n6691), .Q(n3920) );
  nnd2s3 U2410 ( .DIN1(n3923), .DIN2(n6674), .Q(n3918) );
  nnd2s3 U2411 ( .DIN1(n6601), .DIN2(n2112), .Q(n3917) );
  nnd2s3 U2412 ( .DIN1(n6570), .DIN2(n2049), .Q(n3916) );
  nor2s3 U2413 ( .DIN1(n6789), .DIN2(n2112), .Q(WX4425) );
  nor2s3 U2414 ( .DIN1(n5652), .DIN2(n6777), .Q(WX4423) );
  nor2s3 U2415 ( .DIN1(n5653), .DIN2(n6777), .Q(WX4421) );
  nor2s3 U2416 ( .DIN1(n5654), .DIN2(n6777), .Q(WX4419) );
  nor2s3 U2417 ( .DIN1(n5655), .DIN2(n6777), .Q(WX4417) );
  nor2s3 U2418 ( .DIN1(n5656), .DIN2(n6777), .Q(WX4415) );
  nor2s3 U2419 ( .DIN1(n5657), .DIN2(n6777), .Q(WX4413) );
  nor2s3 U2420 ( .DIN1(n5658), .DIN2(n6777), .Q(WX4411) );
  nor2s3 U2421 ( .DIN1(n5659), .DIN2(n6776), .Q(WX4409) );
  nor2s3 U2422 ( .DIN1(n5660), .DIN2(n6776), .Q(WX4407) );
  nor2s3 U2423 ( .DIN1(n5661), .DIN2(n6776), .Q(WX4405) );
  nor2s3 U2424 ( .DIN1(n5662), .DIN2(n6776), .Q(WX4403) );
  nor2s3 U2425 ( .DIN1(n5663), .DIN2(n6776), .Q(WX4401) );
  nor2s3 U2426 ( .DIN1(n5664), .DIN2(n6776), .Q(WX4399) );
  nor2s3 U2427 ( .DIN1(n5665), .DIN2(n6776), .Q(WX4397) );
  nor2s3 U2428 ( .DIN1(n5666), .DIN2(n6776), .Q(WX4395) );
  nor2s3 U2429 ( .DIN1(n5667), .DIN2(n6776), .Q(WX4393) );
  nor2s3 U2430 ( .DIN1(n5668), .DIN2(n6776), .Q(WX4391) );
  nor2s3 U2431 ( .DIN1(n5669), .DIN2(n6783), .Q(WX4389) );
  nor2s3 U2432 ( .DIN1(n5670), .DIN2(n6776), .Q(WX4387) );
  nor2s3 U2433 ( .DIN1(n5671), .DIN2(n6777), .Q(WX4385) );
  nor2s3 U2434 ( .DIN1(n5672), .DIN2(n6777), .Q(WX4383) );
  nor2s3 U2435 ( .DIN1(n5673), .DIN2(n6778), .Q(WX4381) );
  nor2s3 U2436 ( .DIN1(n5674), .DIN2(n6778), .Q(WX4379) );
  nor2s3 U2437 ( .DIN1(n5675), .DIN2(n6778), .Q(WX4377) );
  nor2s3 U2438 ( .DIN1(n5676), .DIN2(n6779), .Q(WX4375) );
  nor2s3 U2439 ( .DIN1(n5677), .DIN2(n6779), .Q(WX4373) );
  nor2s3 U2440 ( .DIN1(n5678), .DIN2(n6779), .Q(WX4371) );
  nor2s3 U2441 ( .DIN1(n5679), .DIN2(n6779), .Q(WX4369) );
  nor2s3 U2442 ( .DIN1(n5680), .DIN2(n6779), .Q(WX4367) );
  nor2s3 U2443 ( .DIN1(n5681), .DIN2(n6779), .Q(WX4365) );
  nor2s3 U2444 ( .DIN1(n5682), .DIN2(n6779), .Q(WX4363) );
  nor2s3 U2445 ( .DIN1(n6804), .DIN2(n3924), .Q(WX3912) );
  xor2s3 U2446 ( .DIN1(n5821), .DIN2(n6109), .Q(n3924) );
  nor2s3 U2447 ( .DIN1(n6804), .DIN2(n3925), .Q(WX3910) );
  xor2s3 U2448 ( .DIN1(n5816), .DIN2(n6100), .Q(n3925) );
  nor2s3 U2449 ( .DIN1(n6804), .DIN2(n3926), .Q(WX3908) );
  xor2s3 U2450 ( .DIN1(n5811), .DIN2(n6091), .Q(n3926) );
  nor2s3 U2451 ( .DIN1(n6804), .DIN2(n3927), .Q(WX3906) );
  xor2s3 U2452 ( .DIN1(n5806), .DIN2(n6082), .Q(n3927) );
  nor2s3 U2453 ( .DIN1(n6804), .DIN2(n3928), .Q(WX3904) );
  xor2s3 U2454 ( .DIN1(n5801), .DIN2(n6073), .Q(n3928) );
  nor2s3 U2455 ( .DIN1(n6804), .DIN2(n3929), .Q(WX3902) );
  xor2s3 U2456 ( .DIN1(n5796), .DIN2(n6064), .Q(n3929) );
  nor2s3 U2457 ( .DIN1(n6804), .DIN2(n3930), .Q(WX3900) );
  xor2s3 U2458 ( .DIN1(n5791), .DIN2(n6055), .Q(n3930) );
  nor2s3 U2459 ( .DIN1(n6804), .DIN2(n3931), .Q(WX3898) );
  xor2s3 U2460 ( .DIN1(n5786), .DIN2(n6046), .Q(n3931) );
  nor2s3 U2461 ( .DIN1(n6804), .DIN2(n3932), .Q(WX3896) );
  xor2s3 U2462 ( .DIN1(n5781), .DIN2(n6037), .Q(n3932) );
  nor2s3 U2463 ( .DIN1(n6804), .DIN2(n3933), .Q(WX3894) );
  xor2s3 U2464 ( .DIN1(n5776), .DIN2(n6028), .Q(n3933) );
  nor2s3 U2465 ( .DIN1(n6804), .DIN2(n3934), .Q(WX3892) );
  xor2s3 U2466 ( .DIN1(n5771), .DIN2(n6019), .Q(n3934) );
  nor2s3 U2467 ( .DIN1(n6804), .DIN2(n3935), .Q(WX3890) );
  xor2s3 U2468 ( .DIN1(n5766), .DIN2(n6010), .Q(n3935) );
  nor2s3 U2469 ( .DIN1(n6804), .DIN2(n3936), .Q(WX3888) );
  xor2s3 U2470 ( .DIN1(n5761), .DIN2(n6001), .Q(n3936) );
  nor2s3 U2471 ( .DIN1(n6803), .DIN2(n3937), .Q(WX3886) );
  xor2s3 U2472 ( .DIN1(n5756), .DIN2(n5992), .Q(n3937) );
  nor2s3 U2473 ( .DIN1(n6803), .DIN2(n3938), .Q(WX3884) );
  xor2s3 U2474 ( .DIN1(n5751), .DIN2(n5983), .Q(n3938) );
  nor2s3 U2475 ( .DIN1(n3939), .DIN2(n6779), .Q(WX3882) );
  xnr2s3 U2476 ( .DIN1(n5974), .DIN2(n3940), .Q(n3939) );
  xor2s3 U2477 ( .DIN1(n5746), .DIN2(n5826), .Q(n3940) );
  nor2s3 U2478 ( .DIN1(n6803), .DIN2(n3941), .Q(WX3880) );
  xor2s3 U2479 ( .DIN1(n5742), .DIN2(n3315), .Q(n3941) );
  nor2s3 U2480 ( .DIN1(n6803), .DIN2(n3942), .Q(WX3878) );
  xor2s3 U2481 ( .DIN1(n5738), .DIN2(n3313), .Q(n3942) );
  nor2s3 U2482 ( .DIN1(n6803), .DIN2(n3943), .Q(WX3876) );
  xor2s3 U2483 ( .DIN1(n5734), .DIN2(n3311), .Q(n3943) );
  nor2s3 U2484 ( .DIN1(n6803), .DIN2(n3944), .Q(WX3874) );
  xor2s3 U2485 ( .DIN1(n5730), .DIN2(n3309), .Q(n3944) );
  nor2s3 U2486 ( .DIN1(n3945), .DIN2(n6779), .Q(WX3872) );
  xnr2s3 U2487 ( .DIN1(n3307), .DIN2(n3946), .Q(n3945) );
  xor2s3 U2488 ( .DIN1(n5726), .DIN2(n5826), .Q(n3946) );
  nor2s3 U2489 ( .DIN1(n6803), .DIN2(n3947), .Q(WX3870) );
  xor2s3 U2490 ( .DIN1(n5722), .DIN2(n3305), .Q(n3947) );
  nor2s3 U2491 ( .DIN1(n6803), .DIN2(n3948), .Q(WX3868) );
  xor2s3 U2492 ( .DIN1(n5718), .DIN2(n3303), .Q(n3948) );
  nor2s3 U2493 ( .DIN1(n6803), .DIN2(n3949), .Q(WX3866) );
  xor2s3 U2494 ( .DIN1(n5714), .DIN2(n3301), .Q(n3949) );
  nor2s3 U2495 ( .DIN1(n6803), .DIN2(n3950), .Q(WX3864) );
  xor2s3 U2496 ( .DIN1(n5710), .DIN2(n3299), .Q(n3950) );
  nor2s3 U2497 ( .DIN1(n6803), .DIN2(n3951), .Q(WX3862) );
  xor2s3 U2498 ( .DIN1(n5706), .DIN2(n3297), .Q(n3951) );
  nor2s3 U2499 ( .DIN1(n6803), .DIN2(n3952), .Q(WX3860) );
  xor2s3 U2500 ( .DIN1(n5702), .DIN2(n3295), .Q(n3952) );
  nor2s3 U2501 ( .DIN1(n3953), .DIN2(n6780), .Q(WX3858) );
  xnr2s3 U2502 ( .DIN1(n3293), .DIN2(n3954), .Q(n3953) );
  xor2s3 U2503 ( .DIN1(n5698), .DIN2(n5826), .Q(n3954) );
  nor2s3 U2504 ( .DIN1(n6802), .DIN2(n3955), .Q(WX3856) );
  xor2s3 U2505 ( .DIN1(n5694), .DIN2(n3291), .Q(n3955) );
  nor2s3 U2506 ( .DIN1(n6802), .DIN2(n3956), .Q(WX3854) );
  xor2s3 U2507 ( .DIN1(n5690), .DIN2(n3289), .Q(n3956) );
  nor2s3 U2508 ( .DIN1(n6802), .DIN2(n3957), .Q(WX3852) );
  xor2s3 U2509 ( .DIN1(n5686), .DIN2(n3287), .Q(n3957) );
  nor2s3 U2510 ( .DIN1(n6802), .DIN2(n3958), .Q(WX3850) );
  xor2s3 U2511 ( .DIN1(n5826), .DIN2(n3285), .Q(n3958) );
  nor2s3 U2512 ( .DIN1(n5861), .DIN2(n6780), .Q(WX3484) );
  nor2s3 U2513 ( .DIN1(n5868), .DIN2(n6780), .Q(WX3482) );
  nor2s3 U2514 ( .DIN1(n5875), .DIN2(n6780), .Q(WX3480) );
  nor2s3 U2515 ( .DIN1(n5882), .DIN2(n6780), .Q(WX3478) );
  nor2s3 U2516 ( .DIN1(n5889), .DIN2(n6780), .Q(WX3476) );
  nor2s3 U2517 ( .DIN1(n5896), .DIN2(n6780), .Q(WX3474) );
  nor2s3 U2518 ( .DIN1(n5903), .DIN2(n6780), .Q(WX3472) );
  nor2s3 U2519 ( .DIN1(n5910), .DIN2(n6780), .Q(WX3470) );
  nor2s3 U2520 ( .DIN1(n5917), .DIN2(n6781), .Q(WX3468) );
  nor2s3 U2521 ( .DIN1(n5924), .DIN2(n6781), .Q(WX3466) );
  nor2s3 U2522 ( .DIN1(n5931), .DIN2(n6781), .Q(WX3464) );
  nor2s3 U2523 ( .DIN1(n5938), .DIN2(n6781), .Q(WX3462) );
  nor2s3 U2524 ( .DIN1(n5945), .DIN2(n6781), .Q(WX3460) );
  nor2s3 U2525 ( .DIN1(n5952), .DIN2(n6781), .Q(WX3458) );
  nor2s3 U2526 ( .DIN1(n5959), .DIN2(n6781), .Q(WX3456) );
  nor2s3 U2527 ( .DIN1(n5966), .DIN2(n6781), .Q(WX3454) );
  nor2s3 U2528 ( .DIN1(n5973), .DIN2(n6781), .Q(WX3452) );
  nor2s3 U2529 ( .DIN1(n5982), .DIN2(n6781), .Q(WX3450) );
  nor2s3 U2530 ( .DIN1(n5991), .DIN2(n6781), .Q(WX3448) );
  nor2s3 U2531 ( .DIN1(n6000), .DIN2(n6782), .Q(WX3446) );
  nor2s3 U2532 ( .DIN1(n6009), .DIN2(n6782), .Q(WX3444) );
  nor2s3 U2533 ( .DIN1(n6018), .DIN2(n6782), .Q(WX3442) );
  nor2s3 U2534 ( .DIN1(n6027), .DIN2(n6782), .Q(WX3440) );
  nor2s3 U2535 ( .DIN1(n6036), .DIN2(n6782), .Q(WX3438) );
  nor2s3 U2536 ( .DIN1(n6045), .DIN2(n6782), .Q(WX3436) );
  nor2s3 U2537 ( .DIN1(n6054), .DIN2(n6782), .Q(WX3434) );
  nor2s3 U2538 ( .DIN1(n6063), .DIN2(n6783), .Q(WX3432) );
  nor2s3 U2539 ( .DIN1(n6072), .DIN2(n6787), .Q(WX3430) );
  nor2s3 U2540 ( .DIN1(n6081), .DIN2(n6787), .Q(WX3428) );
  nor2s3 U2541 ( .DIN1(n6090), .DIN2(n6785), .Q(WX3426) );
  nor2s3 U2542 ( .DIN1(n6099), .DIN2(n6785), .Q(WX3424) );
  nor2s3 U2543 ( .DIN1(n6108), .DIN2(n6785), .Q(WX3422) );
  nor2s3 U2544 ( .DIN1(n5860), .DIN2(n6785), .Q(WX3420) );
  nor2s3 U2545 ( .DIN1(n5867), .DIN2(n6786), .Q(WX3418) );
  nor2s3 U2546 ( .DIN1(n5874), .DIN2(n6785), .Q(WX3416) );
  nor2s3 U2547 ( .DIN1(n5881), .DIN2(n6785), .Q(WX3414) );
  nor2s3 U2548 ( .DIN1(n5888), .DIN2(n6785), .Q(WX3412) );
  nor2s3 U2549 ( .DIN1(n5895), .DIN2(n6785), .Q(WX3410) );
  nor2s3 U2550 ( .DIN1(n5902), .DIN2(n6785), .Q(WX3408) );
  nor2s3 U2551 ( .DIN1(n5909), .DIN2(n6785), .Q(WX3406) );
  nor2s3 U2552 ( .DIN1(n5916), .DIN2(n6784), .Q(WX3404) );
  nor2s3 U2553 ( .DIN1(n5923), .DIN2(n6784), .Q(WX3402) );
  nor2s3 U2554 ( .DIN1(n5930), .DIN2(n6784), .Q(WX3400) );
  nor2s3 U2555 ( .DIN1(n5937), .DIN2(n6784), .Q(WX3398) );
  nor2s3 U2556 ( .DIN1(n5944), .DIN2(n6784), .Q(WX3396) );
  nor2s3 U2557 ( .DIN1(n5951), .DIN2(n6784), .Q(WX3394) );
  nor2s3 U2558 ( .DIN1(n5958), .DIN2(n6784), .Q(WX3392) );
  nor2s3 U2559 ( .DIN1(n5965), .DIN2(n6784), .Q(WX3390) );
  and2s3 U2560 ( .DIN1(RESET), .DIN2(n5972), .Q(WX3388) );
  and2s3 U2561 ( .DIN1(RESET), .DIN2(n5981), .Q(WX3386) );
  and2s3 U2562 ( .DIN1(RESET), .DIN2(n5990), .Q(WX3384) );
  and2s3 U2563 ( .DIN1(RESET), .DIN2(n5999), .Q(WX3382) );
  and2s3 U2564 ( .DIN1(RESET), .DIN2(n6008), .Q(WX3380) );
  and2s3 U2565 ( .DIN1(RESET), .DIN2(n6017), .Q(WX3378) );
  and2s3 U2566 ( .DIN1(RESET), .DIN2(n6026), .Q(WX3376) );
  and2s3 U2567 ( .DIN1(RESET), .DIN2(n6035), .Q(WX3374) );
  and2s3 U2568 ( .DIN1(RESET), .DIN2(n6044), .Q(WX3372) );
  and2s3 U2569 ( .DIN1(RESET), .DIN2(n6053), .Q(WX3370) );
  and2s3 U2570 ( .DIN1(RESET), .DIN2(n6062), .Q(WX3368) );
  and2s3 U2571 ( .DIN1(RESET), .DIN2(n6071), .Q(WX3366) );
  and2s3 U2572 ( .DIN1(RESET), .DIN2(n6080), .Q(WX3364) );
  and2s3 U2573 ( .DIN1(RESET), .DIN2(n6089), .Q(WX3362) );
  and2s3 U2574 ( .DIN1(RESET), .DIN2(n6098), .Q(WX3360) );
  and2s3 U2575 ( .DIN1(RESET), .DIN2(n6107), .Q(WX3358) );
  and2s3 U2576 ( .DIN1(RESET), .DIN2(n5859), .Q(WX3356) );
  and2s3 U2577 ( .DIN1(RESET), .DIN2(n5866), .Q(WX3354) );
  and2s3 U2578 ( .DIN1(RESET), .DIN2(n5873), .Q(WX3352) );
  and2s3 U2579 ( .DIN1(RESET), .DIN2(n5880), .Q(WX3350) );
  and2s3 U2580 ( .DIN1(RESET), .DIN2(n5887), .Q(WX3348) );
  and2s3 U2581 ( .DIN1(RESET), .DIN2(n5894), .Q(WX3346) );
  and2s3 U2582 ( .DIN1(RESET), .DIN2(n5901), .Q(WX3344) );
  and2s3 U2583 ( .DIN1(RESET), .DIN2(n5908), .Q(WX3342) );
  and2s3 U2584 ( .DIN1(RESET), .DIN2(n5915), .Q(WX3340) );
  and2s3 U2585 ( .DIN1(RESET), .DIN2(n5922), .Q(WX3338) );
  and2s3 U2586 ( .DIN1(RESET), .DIN2(n5929), .Q(WX3336) );
  and2s3 U2587 ( .DIN1(RESET), .DIN2(n5936), .Q(WX3334) );
  and2s3 U2588 ( .DIN1(RESET), .DIN2(n5943), .Q(WX3332) );
  and2s3 U2589 ( .DIN1(RESET), .DIN2(n5950), .Q(WX3330) );
  and2s3 U2590 ( .DIN1(RESET), .DIN2(n5957), .Q(WX3328) );
  and2s3 U2591 ( .DIN1(RESET), .DIN2(n5964), .Q(WX3326) );
  nor2s3 U2592 ( .DIN1(n5971), .DIN2(n6784), .Q(WX3324) );
  nor2s3 U2593 ( .DIN1(n5980), .DIN2(n6784), .Q(WX3322) );
  nor2s3 U2594 ( .DIN1(n5989), .DIN2(n6784), .Q(WX3320) );
  nor2s3 U2595 ( .DIN1(n5998), .DIN2(n6784), .Q(WX3318) );
  nor2s3 U2596 ( .DIN1(n6007), .DIN2(n6783), .Q(WX3316) );
  nor2s3 U2597 ( .DIN1(n6016), .DIN2(n6783), .Q(WX3314) );
  nor2s3 U2598 ( .DIN1(n6025), .DIN2(n6783), .Q(WX3312) );
  nor2s3 U2599 ( .DIN1(n6034), .DIN2(n6783), .Q(WX3310) );
  nor2s3 U2600 ( .DIN1(n6043), .DIN2(n6783), .Q(WX3308) );
  nor2s3 U2601 ( .DIN1(n6052), .DIN2(n6783), .Q(WX3306) );
  nor2s3 U2602 ( .DIN1(n6061), .DIN2(n6783), .Q(WX3304) );
  nor2s3 U2603 ( .DIN1(n6070), .DIN2(n6783), .Q(WX3302) );
  nor2s3 U2604 ( .DIN1(n6079), .DIN2(n6766), .Q(WX3300) );
  nor2s3 U2605 ( .DIN1(n6088), .DIN2(n6766), .Q(WX3298) );
  nor2s3 U2606 ( .DIN1(n6097), .DIN2(n6765), .Q(WX3296) );
  nor2s3 U2607 ( .DIN1(n6106), .DIN2(n6765), .Q(WX3294) );
  nnd4s2 U2608 ( .DIN1(n3959), .DIN2(n3960), .DIN3(n3961), .DIN4(n3962), .Q(
        WX3292) );
  nnd2s3 U2609 ( .DIN1(n3690), .DIN2(n6643), .Q(n3962) );
  xor2s3 U2610 ( .DIN1(n3963), .DIN2(n3964), .Q(n3690) );
  xor2s3 U2611 ( .DIN1(n5683), .DIN2(n5684), .Q(n3964) );
  xnr2s3 U2612 ( .DIN1(n3269), .DIN2(n5685), .Q(n3963) );
  nnd2s3 U2613 ( .DIN1(n3965), .DIN2(n6674), .Q(n3961) );
  nnd2s3 U2614 ( .DIN1(n6601), .DIN2(n2145), .Q(n3960) );
  nnd2s3 U2615 ( .DIN1(n6570), .DIN2(n2144), .Q(n3959) );
  nnd4s2 U2616 ( .DIN1(n3966), .DIN2(n3967), .DIN3(n3968), .DIN4(n3969), .Q(
        WX3290) );
  nnd2s3 U2617 ( .DIN1(n3697), .DIN2(n6643), .Q(n3969) );
  xor2s3 U2618 ( .DIN1(n3970), .DIN2(n3971), .Q(n3697) );
  xor2s3 U2619 ( .DIN1(n5687), .DIN2(n5688), .Q(n3971) );
  xnr2s3 U2620 ( .DIN1(n3270), .DIN2(n5689), .Q(n3970) );
  nnd2s3 U2621 ( .DIN1(n3972), .DIN2(n6674), .Q(n3968) );
  nnd2s3 U2622 ( .DIN1(n6601), .DIN2(n2146), .Q(n3967) );
  nnd2s3 U2623 ( .DIN1(n6570), .DIN2(n2143), .Q(n3966) );
  nnd4s2 U2624 ( .DIN1(n3973), .DIN2(n3974), .DIN3(n3975), .DIN4(n3976), .Q(
        WX3288) );
  nnd2s3 U2625 ( .DIN1(n3704), .DIN2(n6643), .Q(n3976) );
  xor2s3 U2626 ( .DIN1(n3977), .DIN2(n3978), .Q(n3704) );
  xor2s3 U2627 ( .DIN1(n5691), .DIN2(n5692), .Q(n3978) );
  xnr2s3 U2628 ( .DIN1(n3271), .DIN2(n5693), .Q(n3977) );
  nnd2s3 U2629 ( .DIN1(n3979), .DIN2(n6674), .Q(n3975) );
  nnd2s3 U2630 ( .DIN1(n6601), .DIN2(n2147), .Q(n3974) );
  nnd2s3 U2631 ( .DIN1(n6570), .DIN2(n2142), .Q(n3973) );
  nnd4s2 U2632 ( .DIN1(n3980), .DIN2(n3981), .DIN3(n3982), .DIN4(n3983), .Q(
        WX3286) );
  nnd2s3 U2633 ( .DIN1(n3711), .DIN2(n6643), .Q(n3983) );
  xor2s3 U2634 ( .DIN1(n3984), .DIN2(n3985), .Q(n3711) );
  xor2s3 U2635 ( .DIN1(n5695), .DIN2(n5696), .Q(n3985) );
  xnr2s3 U2636 ( .DIN1(n3272), .DIN2(n5697), .Q(n3984) );
  nnd2s3 U2637 ( .DIN1(n3986), .DIN2(n6674), .Q(n3982) );
  nnd2s3 U2638 ( .DIN1(n6601), .DIN2(n2148), .Q(n3981) );
  nnd2s3 U2639 ( .DIN1(n6570), .DIN2(n2141), .Q(n3980) );
  nnd4s2 U2640 ( .DIN1(n3987), .DIN2(n3988), .DIN3(n3989), .DIN4(n3990), .Q(
        WX3284) );
  nnd2s3 U2641 ( .DIN1(n3718), .DIN2(n6643), .Q(n3990) );
  xor2s3 U2642 ( .DIN1(n3991), .DIN2(n3992), .Q(n3718) );
  xor2s3 U2643 ( .DIN1(n5699), .DIN2(n5700), .Q(n3992) );
  xnr2s3 U2644 ( .DIN1(n3273), .DIN2(n5701), .Q(n3991) );
  nnd2s3 U2645 ( .DIN1(n3993), .DIN2(n6674), .Q(n3989) );
  nnd2s3 U2646 ( .DIN1(n6601), .DIN2(n2149), .Q(n3988) );
  nnd2s3 U2647 ( .DIN1(n6570), .DIN2(n2140), .Q(n3987) );
  nnd4s2 U2648 ( .DIN1(n3994), .DIN2(n3995), .DIN3(n3996), .DIN4(n3997), .Q(
        WX3282) );
  nnd2s3 U2649 ( .DIN1(n3725), .DIN2(n6643), .Q(n3997) );
  xor2s3 U2650 ( .DIN1(n3998), .DIN2(n3999), .Q(n3725) );
  xor2s3 U2651 ( .DIN1(n5703), .DIN2(n5704), .Q(n3999) );
  xnr2s3 U2652 ( .DIN1(n3274), .DIN2(n5705), .Q(n3998) );
  nnd2s3 U2653 ( .DIN1(n4000), .DIN2(n6674), .Q(n3996) );
  nnd2s3 U2654 ( .DIN1(n6600), .DIN2(n2150), .Q(n3995) );
  nnd2s3 U2655 ( .DIN1(n6569), .DIN2(n2139), .Q(n3994) );
  nnd4s2 U2656 ( .DIN1(n4001), .DIN2(n4002), .DIN3(n4003), .DIN4(n4004), .Q(
        WX3280) );
  nnd2s3 U2657 ( .DIN1(n3732), .DIN2(n6642), .Q(n4004) );
  xor2s3 U2658 ( .DIN1(n4005), .DIN2(n4006), .Q(n3732) );
  xor2s3 U2659 ( .DIN1(n5707), .DIN2(n5708), .Q(n4006) );
  xnr2s3 U2660 ( .DIN1(n3275), .DIN2(n5709), .Q(n4005) );
  nnd2s3 U2661 ( .DIN1(n4007), .DIN2(n6673), .Q(n4003) );
  nnd2s3 U2662 ( .DIN1(n6600), .DIN2(n2151), .Q(n4002) );
  nnd2s3 U2663 ( .DIN1(n6569), .DIN2(n2138), .Q(n4001) );
  nnd4s2 U2664 ( .DIN1(n4008), .DIN2(n4009), .DIN3(n4010), .DIN4(n4011), .Q(
        WX3278) );
  nnd2s3 U2665 ( .DIN1(n3739), .DIN2(n6642), .Q(n4011) );
  xor2s3 U2666 ( .DIN1(n4012), .DIN2(n4013), .Q(n3739) );
  xor2s3 U2667 ( .DIN1(n5711), .DIN2(n5712), .Q(n4013) );
  xnr2s3 U2668 ( .DIN1(n3276), .DIN2(n5713), .Q(n4012) );
  nnd2s3 U2669 ( .DIN1(n4014), .DIN2(n6673), .Q(n4010) );
  nnd2s3 U2670 ( .DIN1(n6600), .DIN2(n2152), .Q(n4009) );
  nnd2s3 U2671 ( .DIN1(n6569), .DIN2(n2137), .Q(n4008) );
  nnd4s2 U2672 ( .DIN1(n4015), .DIN2(n4016), .DIN3(n4017), .DIN4(n4018), .Q(
        WX3276) );
  nnd2s3 U2673 ( .DIN1(n3746), .DIN2(n6642), .Q(n4018) );
  xor2s3 U2674 ( .DIN1(n4019), .DIN2(n4020), .Q(n3746) );
  xor2s3 U2675 ( .DIN1(n5715), .DIN2(n5716), .Q(n4020) );
  xnr2s3 U2676 ( .DIN1(n3277), .DIN2(n5717), .Q(n4019) );
  nnd2s3 U2677 ( .DIN1(n4021), .DIN2(n6673), .Q(n4017) );
  nnd2s3 U2678 ( .DIN1(n6600), .DIN2(n2153), .Q(n4016) );
  nnd2s3 U2679 ( .DIN1(n6569), .DIN2(n2136), .Q(n4015) );
  nnd4s2 U2680 ( .DIN1(n4022), .DIN2(n4023), .DIN3(n4024), .DIN4(n4025), .Q(
        WX3274) );
  nnd2s3 U2681 ( .DIN1(n3753), .DIN2(n6642), .Q(n4025) );
  xor2s3 U2682 ( .DIN1(n4026), .DIN2(n4027), .Q(n3753) );
  xor2s3 U2683 ( .DIN1(n5719), .DIN2(n5720), .Q(n4027) );
  xnr2s3 U2684 ( .DIN1(n3278), .DIN2(n5721), .Q(n4026) );
  nnd2s3 U2685 ( .DIN1(n4028), .DIN2(n6673), .Q(n4024) );
  nnd2s3 U2686 ( .DIN1(n6600), .DIN2(n2154), .Q(n4023) );
  nnd2s3 U2687 ( .DIN1(n6569), .DIN2(n2135), .Q(n4022) );
  nnd4s2 U2688 ( .DIN1(n4029), .DIN2(n4030), .DIN3(n4031), .DIN4(n4032), .Q(
        WX3272) );
  nnd2s3 U2689 ( .DIN1(n3760), .DIN2(n6642), .Q(n4032) );
  xor2s3 U2690 ( .DIN1(n4033), .DIN2(n4034), .Q(n3760) );
  xor2s3 U2691 ( .DIN1(n5723), .DIN2(n5724), .Q(n4034) );
  xnr2s3 U2692 ( .DIN1(n3279), .DIN2(n5725), .Q(n4033) );
  nnd2s3 U2693 ( .DIN1(n4035), .DIN2(n6673), .Q(n4031) );
  nnd2s3 U2694 ( .DIN1(n6600), .DIN2(n2155), .Q(n4030) );
  nnd2s3 U2695 ( .DIN1(n6569), .DIN2(n2134), .Q(n4029) );
  nnd4s2 U2696 ( .DIN1(n4036), .DIN2(n4037), .DIN3(n4038), .DIN4(n4039), .Q(
        WX3270) );
  nnd2s3 U2697 ( .DIN1(n3767), .DIN2(n6642), .Q(n4039) );
  xor2s3 U2698 ( .DIN1(n4040), .DIN2(n4041), .Q(n3767) );
  xor2s3 U2699 ( .DIN1(n5727), .DIN2(n5728), .Q(n4041) );
  xnr2s3 U2700 ( .DIN1(n3280), .DIN2(n5729), .Q(n4040) );
  nnd2s3 U2701 ( .DIN1(n4042), .DIN2(n6673), .Q(n4038) );
  nnd2s3 U2702 ( .DIN1(n6600), .DIN2(n2156), .Q(n4037) );
  nnd2s3 U2703 ( .DIN1(n6569), .DIN2(n2133), .Q(n4036) );
  nnd4s2 U2704 ( .DIN1(n4043), .DIN2(n4044), .DIN3(n4045), .DIN4(n4046), .Q(
        WX3268) );
  nnd2s3 U2705 ( .DIN1(n3774), .DIN2(n6642), .Q(n4046) );
  xor2s3 U2706 ( .DIN1(n4047), .DIN2(n4048), .Q(n3774) );
  xor2s3 U2707 ( .DIN1(n5731), .DIN2(n5732), .Q(n4048) );
  xnr2s3 U2708 ( .DIN1(n3281), .DIN2(n5733), .Q(n4047) );
  nnd2s3 U2709 ( .DIN1(n4049), .DIN2(n6673), .Q(n4045) );
  nnd2s3 U2710 ( .DIN1(n6600), .DIN2(n2157), .Q(n4044) );
  nnd2s3 U2711 ( .DIN1(n6569), .DIN2(n2132), .Q(n4043) );
  nnd4s2 U2712 ( .DIN1(n4050), .DIN2(n4051), .DIN3(n4052), .DIN4(n4053), .Q(
        WX3266) );
  nnd2s3 U2713 ( .DIN1(n3781), .DIN2(n6642), .Q(n4053) );
  xor2s3 U2714 ( .DIN1(n4054), .DIN2(n4055), .Q(n3781) );
  xor2s3 U2715 ( .DIN1(n5735), .DIN2(n5736), .Q(n4055) );
  xnr2s3 U2716 ( .DIN1(n3282), .DIN2(n5737), .Q(n4054) );
  nnd2s3 U2717 ( .DIN1(n4056), .DIN2(n6673), .Q(n4052) );
  nnd2s3 U2718 ( .DIN1(n6600), .DIN2(n2158), .Q(n4051) );
  nnd2s3 U2719 ( .DIN1(n6569), .DIN2(n2131), .Q(n4050) );
  nnd4s2 U2720 ( .DIN1(n4057), .DIN2(n4058), .DIN3(n4059), .DIN4(n4060), .Q(
        WX3264) );
  nnd2s3 U2721 ( .DIN1(n3788), .DIN2(n6642), .Q(n4060) );
  xor2s3 U2722 ( .DIN1(n4061), .DIN2(n4062), .Q(n3788) );
  xor2s3 U2723 ( .DIN1(n5739), .DIN2(n5740), .Q(n4062) );
  xnr2s3 U2724 ( .DIN1(n3283), .DIN2(n5741), .Q(n4061) );
  nnd2s3 U2725 ( .DIN1(n4063), .DIN2(n6673), .Q(n4059) );
  nnd2s3 U2726 ( .DIN1(n6600), .DIN2(n2159), .Q(n4058) );
  nnd2s3 U2727 ( .DIN1(n6569), .DIN2(n2130), .Q(n4057) );
  nnd4s2 U2728 ( .DIN1(n4064), .DIN2(n4065), .DIN3(n4066), .DIN4(n4067), .Q(
        WX3262) );
  nnd2s3 U2729 ( .DIN1(n3795), .DIN2(n6642), .Q(n4067) );
  xor2s3 U2730 ( .DIN1(n4068), .DIN2(n4069), .Q(n3795) );
  xor2s3 U2731 ( .DIN1(n5743), .DIN2(n5744), .Q(n4069) );
  xnr2s3 U2732 ( .DIN1(n3284), .DIN2(n5745), .Q(n4068) );
  nnd2s3 U2733 ( .DIN1(n4070), .DIN2(n6673), .Q(n4066) );
  nnd2s3 U2734 ( .DIN1(n6600), .DIN2(n2160), .Q(n4065) );
  nnd2s3 U2735 ( .DIN1(n6569), .DIN2(n2129), .Q(n4064) );
  nnd4s2 U2736 ( .DIN1(n4071), .DIN2(n4072), .DIN3(n4073), .DIN4(n4074), .Q(
        WX3260) );
  nnd2s3 U2737 ( .DIN1(n3803), .DIN2(n6642), .Q(n4074) );
  xor2s3 U2738 ( .DIN1(n4075), .DIN2(n4076), .Q(n3803) );
  xor2s3 U2739 ( .DIN1(n5749), .DIN2(n4077), .Q(n4076) );
  xor2s3 U2740 ( .DIN1(n5747), .DIN2(n5748), .Q(n4077) );
  xor2s3 U2741 ( .DIN1(n5750), .DIN2(n6691), .Q(n4075) );
  nnd2s3 U2742 ( .DIN1(n4078), .DIN2(n6673), .Q(n4073) );
  nnd2s3 U2743 ( .DIN1(n6600), .DIN2(n2161), .Q(n4072) );
  nnd2s3 U2744 ( .DIN1(n6569), .DIN2(n2128), .Q(n4071) );
  nnd4s2 U2745 ( .DIN1(n4079), .DIN2(n4080), .DIN3(n4081), .DIN4(n4082), .Q(
        WX3258) );
  nnd2s3 U2746 ( .DIN1(n3811), .DIN2(n6642), .Q(n4082) );
  xor2s3 U2747 ( .DIN1(n4083), .DIN2(n4084), .Q(n3811) );
  xor2s3 U2748 ( .DIN1(n5754), .DIN2(n4085), .Q(n4084) );
  xor2s3 U2749 ( .DIN1(n5752), .DIN2(n5753), .Q(n4085) );
  xor2s3 U2750 ( .DIN1(n5755), .DIN2(n6692), .Q(n4083) );
  nnd2s3 U2751 ( .DIN1(n4086), .DIN2(n6673), .Q(n4081) );
  nnd2s3 U2752 ( .DIN1(n6600), .DIN2(n2162), .Q(n4080) );
  nnd2s3 U2753 ( .DIN1(n6569), .DIN2(n2127), .Q(n4079) );
  nnd4s2 U2754 ( .DIN1(n4087), .DIN2(n4088), .DIN3(n4089), .DIN4(n4090), .Q(
        WX3256) );
  nnd2s3 U2755 ( .DIN1(n3819), .DIN2(n6642), .Q(n4090) );
  xor2s3 U2756 ( .DIN1(n4091), .DIN2(n4092), .Q(n3819) );
  xor2s3 U2757 ( .DIN1(n5759), .DIN2(n4093), .Q(n4092) );
  xor2s3 U2758 ( .DIN1(n5757), .DIN2(n5758), .Q(n4093) );
  xor2s3 U2759 ( .DIN1(n5760), .DIN2(n6692), .Q(n4091) );
  nnd2s3 U2760 ( .DIN1(n4094), .DIN2(n6673), .Q(n4089) );
  nnd2s3 U2761 ( .DIN1(n6599), .DIN2(n2163), .Q(n4088) );
  nnd2s3 U2762 ( .DIN1(n6568), .DIN2(n2126), .Q(n4087) );
  nnd4s2 U2763 ( .DIN1(n4095), .DIN2(n4096), .DIN3(n4097), .DIN4(n4098), .Q(
        WX3254) );
  nnd2s3 U2764 ( .DIN1(n3827), .DIN2(n6641), .Q(n4098) );
  xor2s3 U2765 ( .DIN1(n4099), .DIN2(n4100), .Q(n3827) );
  xor2s3 U2766 ( .DIN1(n5764), .DIN2(n4101), .Q(n4100) );
  xor2s3 U2767 ( .DIN1(n5762), .DIN2(n5763), .Q(n4101) );
  xor2s3 U2768 ( .DIN1(n5765), .DIN2(n6692), .Q(n4099) );
  nnd2s3 U2769 ( .DIN1(n4102), .DIN2(n6672), .Q(n4097) );
  nnd2s3 U2770 ( .DIN1(n6599), .DIN2(n2164), .Q(n4096) );
  nnd2s3 U2771 ( .DIN1(n6568), .DIN2(n2125), .Q(n4095) );
  nnd4s2 U2772 ( .DIN1(n4103), .DIN2(n4104), .DIN3(n4105), .DIN4(n4106), .Q(
        WX3252) );
  nnd2s3 U2773 ( .DIN1(n3835), .DIN2(n6641), .Q(n4106) );
  xor2s3 U2774 ( .DIN1(n4107), .DIN2(n4108), .Q(n3835) );
  xor2s3 U2775 ( .DIN1(n5769), .DIN2(n4109), .Q(n4108) );
  xor2s3 U2776 ( .DIN1(n5767), .DIN2(n5768), .Q(n4109) );
  xor2s3 U2777 ( .DIN1(n5770), .DIN2(n6692), .Q(n4107) );
  nnd2s3 U2778 ( .DIN1(n4110), .DIN2(n6672), .Q(n4105) );
  nnd2s3 U2779 ( .DIN1(n6599), .DIN2(n2165), .Q(n4104) );
  nnd2s3 U2780 ( .DIN1(n6568), .DIN2(n2124), .Q(n4103) );
  nnd4s2 U2781 ( .DIN1(n4111), .DIN2(n4112), .DIN3(n4113), .DIN4(n4114), .Q(
        WX3250) );
  nnd2s3 U2782 ( .DIN1(n3843), .DIN2(n6641), .Q(n4114) );
  xor2s3 U2783 ( .DIN1(n4115), .DIN2(n4116), .Q(n3843) );
  xor2s3 U2784 ( .DIN1(n5774), .DIN2(n4117), .Q(n4116) );
  xor2s3 U2785 ( .DIN1(n5772), .DIN2(n5773), .Q(n4117) );
  xor2s3 U2786 ( .DIN1(n5775), .DIN2(n6692), .Q(n4115) );
  nnd2s3 U2787 ( .DIN1(n4118), .DIN2(n6672), .Q(n4113) );
  nnd2s3 U2788 ( .DIN1(n6599), .DIN2(n2166), .Q(n4112) );
  nnd2s3 U2789 ( .DIN1(n6568), .DIN2(n2123), .Q(n4111) );
  nnd4s2 U2790 ( .DIN1(n4119), .DIN2(n4120), .DIN3(n4121), .DIN4(n4122), .Q(
        WX3248) );
  nnd2s3 U2791 ( .DIN1(n3851), .DIN2(n6641), .Q(n4122) );
  xor2s3 U2792 ( .DIN1(n4123), .DIN2(n4124), .Q(n3851) );
  xor2s3 U2793 ( .DIN1(n5779), .DIN2(n4125), .Q(n4124) );
  xor2s3 U2794 ( .DIN1(n5777), .DIN2(n5778), .Q(n4125) );
  xor2s3 U2795 ( .DIN1(n5780), .DIN2(n6692), .Q(n4123) );
  nnd2s3 U2796 ( .DIN1(n4126), .DIN2(n6672), .Q(n4121) );
  nnd2s3 U2797 ( .DIN1(n6599), .DIN2(n2167), .Q(n4120) );
  nnd2s3 U2798 ( .DIN1(n6568), .DIN2(n2122), .Q(n4119) );
  nnd4s2 U2799 ( .DIN1(n4127), .DIN2(n4128), .DIN3(n4129), .DIN4(n4130), .Q(
        WX3246) );
  nnd2s3 U2800 ( .DIN1(n3859), .DIN2(n6641), .Q(n4130) );
  xor2s3 U2801 ( .DIN1(n4131), .DIN2(n4132), .Q(n3859) );
  xor2s3 U2802 ( .DIN1(n5784), .DIN2(n4133), .Q(n4132) );
  xor2s3 U2803 ( .DIN1(n5782), .DIN2(n5783), .Q(n4133) );
  xor2s3 U2804 ( .DIN1(n5785), .DIN2(n6692), .Q(n4131) );
  nnd2s3 U2805 ( .DIN1(n4134), .DIN2(n6672), .Q(n4129) );
  nnd2s3 U2806 ( .DIN1(n6599), .DIN2(n2168), .Q(n4128) );
  nnd2s3 U2807 ( .DIN1(n6568), .DIN2(n2121), .Q(n4127) );
  nnd4s2 U2808 ( .DIN1(n4135), .DIN2(n4136), .DIN3(n4137), .DIN4(n4138), .Q(
        WX3244) );
  nnd2s3 U2809 ( .DIN1(n3867), .DIN2(n6641), .Q(n4138) );
  xor2s3 U2810 ( .DIN1(n4139), .DIN2(n4140), .Q(n3867) );
  xor2s3 U2811 ( .DIN1(n5789), .DIN2(n4141), .Q(n4140) );
  xor2s3 U2812 ( .DIN1(n5787), .DIN2(n5788), .Q(n4141) );
  xor2s3 U2813 ( .DIN1(n5790), .DIN2(n6692), .Q(n4139) );
  nnd2s3 U2814 ( .DIN1(n4142), .DIN2(n6672), .Q(n4137) );
  nnd2s3 U2815 ( .DIN1(n6599), .DIN2(n2169), .Q(n4136) );
  nnd2s3 U2816 ( .DIN1(n6568), .DIN2(n2120), .Q(n4135) );
  nnd4s2 U2817 ( .DIN1(n4143), .DIN2(n4144), .DIN3(n4145), .DIN4(n4146), .Q(
        WX3242) );
  nnd2s3 U2818 ( .DIN1(n3875), .DIN2(n6641), .Q(n4146) );
  xor2s3 U2819 ( .DIN1(n4147), .DIN2(n4148), .Q(n3875) );
  xor2s3 U2820 ( .DIN1(n5794), .DIN2(n4149), .Q(n4148) );
  xor2s3 U2821 ( .DIN1(n5792), .DIN2(n5793), .Q(n4149) );
  xor2s3 U2822 ( .DIN1(n5795), .DIN2(n6692), .Q(n4147) );
  nnd2s3 U2823 ( .DIN1(n4150), .DIN2(n6672), .Q(n4145) );
  nnd2s3 U2824 ( .DIN1(n6599), .DIN2(n2170), .Q(n4144) );
  nnd2s3 U2825 ( .DIN1(n6568), .DIN2(n2119), .Q(n4143) );
  nnd4s2 U2826 ( .DIN1(n4151), .DIN2(n4152), .DIN3(n4153), .DIN4(n4154), .Q(
        WX3240) );
  nnd2s3 U2827 ( .DIN1(n3883), .DIN2(n6641), .Q(n4154) );
  xor2s3 U2828 ( .DIN1(n4155), .DIN2(n4156), .Q(n3883) );
  xor2s3 U2829 ( .DIN1(n5799), .DIN2(n4157), .Q(n4156) );
  xor2s3 U2830 ( .DIN1(n5797), .DIN2(n5798), .Q(n4157) );
  xor2s3 U2831 ( .DIN1(n5800), .DIN2(n6692), .Q(n4155) );
  nnd2s3 U2832 ( .DIN1(n4158), .DIN2(n6672), .Q(n4153) );
  nnd2s3 U2833 ( .DIN1(n6599), .DIN2(n2171), .Q(n4152) );
  nnd2s3 U2834 ( .DIN1(n6568), .DIN2(n2118), .Q(n4151) );
  nnd4s2 U2835 ( .DIN1(n4159), .DIN2(n4160), .DIN3(n4161), .DIN4(n4162), .Q(
        WX3238) );
  nnd2s3 U2836 ( .DIN1(n3891), .DIN2(n6641), .Q(n4162) );
  xor2s3 U2837 ( .DIN1(n4163), .DIN2(n4164), .Q(n3891) );
  xor2s3 U2838 ( .DIN1(n5804), .DIN2(n4165), .Q(n4164) );
  xor2s3 U2839 ( .DIN1(n5802), .DIN2(n5803), .Q(n4165) );
  xor2s3 U2840 ( .DIN1(n5805), .DIN2(n6692), .Q(n4163) );
  nnd2s3 U2841 ( .DIN1(n4166), .DIN2(n6672), .Q(n4161) );
  nnd2s3 U2842 ( .DIN1(n6599), .DIN2(n2172), .Q(n4160) );
  nnd2s3 U2843 ( .DIN1(n6568), .DIN2(n2117), .Q(n4159) );
  nnd4s2 U2844 ( .DIN1(n4167), .DIN2(n4168), .DIN3(n4169), .DIN4(n4170), .Q(
        WX3236) );
  nnd2s3 U2845 ( .DIN1(n3899), .DIN2(n6641), .Q(n4170) );
  xor2s3 U2846 ( .DIN1(n4171), .DIN2(n4172), .Q(n3899) );
  xor2s3 U2847 ( .DIN1(n5809), .DIN2(n4173), .Q(n4172) );
  xor2s3 U2848 ( .DIN1(n5807), .DIN2(n5808), .Q(n4173) );
  xor2s3 U2849 ( .DIN1(n5810), .DIN2(n6692), .Q(n4171) );
  nnd2s3 U2850 ( .DIN1(n4174), .DIN2(n6672), .Q(n4169) );
  nnd2s3 U2851 ( .DIN1(n6599), .DIN2(n2173), .Q(n4168) );
  nnd2s3 U2852 ( .DIN1(n6568), .DIN2(n2116), .Q(n4167) );
  nnd4s2 U2853 ( .DIN1(n4175), .DIN2(n4176), .DIN3(n4177), .DIN4(n4178), .Q(
        WX3234) );
  nnd2s3 U2854 ( .DIN1(n3907), .DIN2(n6641), .Q(n4178) );
  xor2s3 U2855 ( .DIN1(n4179), .DIN2(n4180), .Q(n3907) );
  xor2s3 U2856 ( .DIN1(n5814), .DIN2(n4181), .Q(n4180) );
  xor2s3 U2857 ( .DIN1(n5812), .DIN2(n5813), .Q(n4181) );
  xor2s3 U2858 ( .DIN1(n5815), .DIN2(n6693), .Q(n4179) );
  nnd2s3 U2859 ( .DIN1(n4182), .DIN2(n6672), .Q(n4177) );
  nnd2s3 U2860 ( .DIN1(n6599), .DIN2(n2174), .Q(n4176) );
  nnd2s3 U2861 ( .DIN1(n6568), .DIN2(n2115), .Q(n4175) );
  nnd4s2 U2862 ( .DIN1(n4183), .DIN2(n4184), .DIN3(n4185), .DIN4(n4186), .Q(
        WX3232) );
  nnd2s3 U2863 ( .DIN1(n3915), .DIN2(n6641), .Q(n4186) );
  xor2s3 U2864 ( .DIN1(n4187), .DIN2(n4188), .Q(n3915) );
  xor2s3 U2865 ( .DIN1(n5819), .DIN2(n4189), .Q(n4188) );
  xor2s3 U2866 ( .DIN1(n5817), .DIN2(n5818), .Q(n4189) );
  xor2s3 U2867 ( .DIN1(n5820), .DIN2(n6693), .Q(n4187) );
  nnd2s3 U2868 ( .DIN1(n4190), .DIN2(n6672), .Q(n4185) );
  nnd2s3 U2869 ( .DIN1(n6599), .DIN2(n2175), .Q(n4184) );
  nnd2s3 U2870 ( .DIN1(n6568), .DIN2(n2114), .Q(n4183) );
  nnd4s2 U2871 ( .DIN1(n4191), .DIN2(n4192), .DIN3(n4193), .DIN4(n4194), .Q(
        WX3230) );
  nnd2s3 U2872 ( .DIN1(n3923), .DIN2(n6640), .Q(n4194) );
  xor2s3 U2873 ( .DIN1(n4195), .DIN2(n4196), .Q(n3923) );
  xor2s3 U2874 ( .DIN1(n5824), .DIN2(n4197), .Q(n4196) );
  xor2s3 U2875 ( .DIN1(n5822), .DIN2(n5823), .Q(n4197) );
  xor2s3 U2876 ( .DIN1(n5825), .DIN2(n6693), .Q(n4195) );
  nnd2s3 U2877 ( .DIN1(n4198), .DIN2(n6671), .Q(n4193) );
  nnd2s3 U2878 ( .DIN1(n6598), .DIN2(n2176), .Q(n4192) );
  nnd2s3 U2879 ( .DIN1(n6567), .DIN2(n2113), .Q(n4191) );
  nor2s3 U2880 ( .DIN1(n6802), .DIN2(n2176), .Q(WX3132) );
  nor2s3 U2881 ( .DIN1(n5828), .DIN2(n6765), .Q(WX3130) );
  nor2s3 U2882 ( .DIN1(n5829), .DIN2(n6765), .Q(WX3128) );
  nor2s3 U2883 ( .DIN1(n5830), .DIN2(n6765), .Q(WX3126) );
  nor2s3 U2884 ( .DIN1(n5831), .DIN2(n6765), .Q(WX3124) );
  nor2s3 U2885 ( .DIN1(n5832), .DIN2(n6765), .Q(WX3122) );
  nor2s3 U2886 ( .DIN1(n5833), .DIN2(n6765), .Q(WX3120) );
  nor2s3 U2887 ( .DIN1(n5834), .DIN2(n6765), .Q(WX3118) );
  nor2s3 U2888 ( .DIN1(n5835), .DIN2(n6765), .Q(WX3116) );
  nor2s3 U2889 ( .DIN1(n5836), .DIN2(n6765), .Q(WX3114) );
  nor2s3 U2890 ( .DIN1(n5837), .DIN2(n6765), .Q(WX3112) );
  nor2s3 U2891 ( .DIN1(n5838), .DIN2(n6764), .Q(WX3110) );
  nor2s3 U2892 ( .DIN1(n5839), .DIN2(n6764), .Q(WX3108) );
  nor2s3 U2893 ( .DIN1(n5840), .DIN2(n6764), .Q(WX3106) );
  nor2s3 U2894 ( .DIN1(n5841), .DIN2(n6764), .Q(WX3104) );
  nor2s3 U2895 ( .DIN1(n5842), .DIN2(n6764), .Q(WX3102) );
  nor2s3 U2896 ( .DIN1(n5843), .DIN2(n6764), .Q(WX3100) );
  nor2s3 U2897 ( .DIN1(n5844), .DIN2(n6764), .Q(WX3098) );
  nor2s3 U2898 ( .DIN1(n5845), .DIN2(n6764), .Q(WX3096) );
  nor2s3 U2899 ( .DIN1(n5846), .DIN2(n6764), .Q(WX3094) );
  nor2s3 U2900 ( .DIN1(n5847), .DIN2(n6764), .Q(WX3092) );
  nor2s3 U2901 ( .DIN1(n5848), .DIN2(n6764), .Q(WX3090) );
  nor2s3 U2902 ( .DIN1(n5849), .DIN2(n6764), .Q(WX3088) );
  nor2s3 U2903 ( .DIN1(n5850), .DIN2(n6763), .Q(WX3086) );
  nor2s3 U2904 ( .DIN1(n5851), .DIN2(n6763), .Q(WX3084) );
  nor2s3 U2905 ( .DIN1(n5852), .DIN2(n6763), .Q(WX3082) );
  nor2s3 U2906 ( .DIN1(n5853), .DIN2(n6763), .Q(WX3080) );
  nor2s3 U2907 ( .DIN1(n5854), .DIN2(n6763), .Q(WX3078) );
  nor2s3 U2908 ( .DIN1(n5855), .DIN2(n6763), .Q(WX3076) );
  nor2s3 U2909 ( .DIN1(n5856), .DIN2(n6763), .Q(WX3074) );
  nor2s3 U2910 ( .DIN1(n5857), .DIN2(n6763), .Q(WX3072) );
  nor2s3 U2911 ( .DIN1(n5858), .DIN2(n6763), .Q(WX3070) );
  nor2s3 U2912 ( .DIN1(n6796), .DIN2(n4199), .Q(WX2619) );
  xor2s3 U2913 ( .DIN1(n6105), .DIN2(n6113), .Q(n4199) );
  nor2s3 U2914 ( .DIN1(n6796), .DIN2(n4200), .Q(WX2617) );
  xor2s3 U2915 ( .DIN1(n6096), .DIN2(n6104), .Q(n4200) );
  nor2s3 U2916 ( .DIN1(n6796), .DIN2(n4201), .Q(WX2615) );
  xor2s3 U2917 ( .DIN1(n6087), .DIN2(n6095), .Q(n4201) );
  nor2s3 U2918 ( .DIN1(n6796), .DIN2(n4202), .Q(WX2613) );
  xor2s3 U2919 ( .DIN1(n6078), .DIN2(n6086), .Q(n4202) );
  nor2s3 U2920 ( .DIN1(n6796), .DIN2(n4203), .Q(WX2611) );
  xor2s3 U2921 ( .DIN1(n6069), .DIN2(n6077), .Q(n4203) );
  nor2s3 U2922 ( .DIN1(n6796), .DIN2(n4204), .Q(WX2609) );
  xor2s3 U2923 ( .DIN1(n6060), .DIN2(n6068), .Q(n4204) );
  nor2s3 U2924 ( .DIN1(n6796), .DIN2(n4205), .Q(WX2607) );
  xor2s3 U2925 ( .DIN1(n6051), .DIN2(n6059), .Q(n4205) );
  nor2s3 U2926 ( .DIN1(n6796), .DIN2(n4206), .Q(WX2605) );
  xor2s3 U2927 ( .DIN1(n6042), .DIN2(n6050), .Q(n4206) );
  nor2s3 U2928 ( .DIN1(n6796), .DIN2(n4207), .Q(WX2603) );
  xor2s3 U2929 ( .DIN1(n6033), .DIN2(n6041), .Q(n4207) );
  nor2s3 U2930 ( .DIN1(n6796), .DIN2(n4208), .Q(WX2601) );
  xor2s3 U2931 ( .DIN1(n6024), .DIN2(n6032), .Q(n4208) );
  nor2s3 U2932 ( .DIN1(n6796), .DIN2(n4209), .Q(WX2599) );
  xor2s3 U2933 ( .DIN1(n6015), .DIN2(n6023), .Q(n4209) );
  nor2s3 U2934 ( .DIN1(n6797), .DIN2(n4210), .Q(WX2597) );
  xor2s3 U2935 ( .DIN1(n6006), .DIN2(n6014), .Q(n4210) );
  nor2s3 U2936 ( .DIN1(n6797), .DIN2(n4211), .Q(WX2595) );
  xor2s3 U2937 ( .DIN1(n5997), .DIN2(n6005), .Q(n4211) );
  nor2s3 U2938 ( .DIN1(n6797), .DIN2(n4212), .Q(WX2593) );
  xor2s3 U2939 ( .DIN1(n5988), .DIN2(n5996), .Q(n4212) );
  nor2s3 U2940 ( .DIN1(n6797), .DIN2(n4213), .Q(WX2591) );
  xor2s3 U2941 ( .DIN1(n5979), .DIN2(n5987), .Q(n4213) );
  nor2s3 U2942 ( .DIN1(n4214), .DIN2(n6763), .Q(WX2589) );
  xor2s3 U2943 ( .DIN1(n2177), .DIN2(n4215), .Q(n4214) );
  xor2s3 U2944 ( .DIN1(n5970), .DIN2(n5978), .Q(n4215) );
  nor2s3 U2945 ( .DIN1(n6797), .DIN2(n4216), .Q(WX2587) );
  xor2s3 U2946 ( .DIN1(n5963), .DIN2(n3316), .Q(n4216) );
  nor2s3 U2947 ( .DIN1(n6797), .DIN2(n4217), .Q(WX2585) );
  xor2s3 U2948 ( .DIN1(n5956), .DIN2(n3314), .Q(n4217) );
  nor2s3 U2949 ( .DIN1(n6797), .DIN2(n4218), .Q(WX2583) );
  xor2s3 U2950 ( .DIN1(n5949), .DIN2(n3312), .Q(n4218) );
  nor2s3 U2951 ( .DIN1(n6797), .DIN2(n4219), .Q(WX2581) );
  xor2s3 U2952 ( .DIN1(n5942), .DIN2(n3310), .Q(n4219) );
  nor2s3 U2953 ( .DIN1(n4220), .DIN2(n6763), .Q(WX2579) );
  xnr2s3 U2954 ( .DIN1(n3308), .DIN2(n4221), .Q(n4220) );
  xor2s3 U2955 ( .DIN1(n5935), .DIN2(n6114), .Q(n4221) );
  nor2s3 U2956 ( .DIN1(n6797), .DIN2(n4222), .Q(WX2577) );
  xor2s3 U2957 ( .DIN1(n5928), .DIN2(n3306), .Q(n4222) );
  nor2s3 U2958 ( .DIN1(n6797), .DIN2(n4223), .Q(WX2575) );
  xor2s3 U2959 ( .DIN1(n5921), .DIN2(n3304), .Q(n4223) );
  nor2s3 U2960 ( .DIN1(n6797), .DIN2(n4224), .Q(WX2573) );
  xor2s3 U2961 ( .DIN1(n5914), .DIN2(n3302), .Q(n4224) );
  nor2s3 U2962 ( .DIN1(n6798), .DIN2(n4225), .Q(WX2571) );
  xor2s3 U2963 ( .DIN1(n5907), .DIN2(n3300), .Q(n4225) );
  nor2s3 U2964 ( .DIN1(n6798), .DIN2(n4226), .Q(WX2569) );
  xor2s3 U2965 ( .DIN1(n5900), .DIN2(n3298), .Q(n4226) );
  nor2s3 U2966 ( .DIN1(n6798), .DIN2(n4227), .Q(WX2567) );
  xor2s3 U2967 ( .DIN1(n5893), .DIN2(n3296), .Q(n4227) );
  nor2s3 U2968 ( .DIN1(n4228), .DIN2(n6763), .Q(WX2565) );
  xnr2s3 U2969 ( .DIN1(n3294), .DIN2(n4229), .Q(n4228) );
  xor2s3 U2970 ( .DIN1(n5886), .DIN2(n6114), .Q(n4229) );
  nor2s3 U2971 ( .DIN1(n6798), .DIN2(n4230), .Q(WX2563) );
  xor2s3 U2972 ( .DIN1(n5879), .DIN2(n3292), .Q(n4230) );
  nor2s3 U2973 ( .DIN1(n6798), .DIN2(n4231), .Q(WX2561) );
  xor2s3 U2974 ( .DIN1(n5872), .DIN2(n3290), .Q(n4231) );
  nor2s3 U2975 ( .DIN1(n6798), .DIN2(n4232), .Q(WX2559) );
  xor2s3 U2976 ( .DIN1(n5865), .DIN2(n3288), .Q(n4232) );
  nor2s3 U2977 ( .DIN1(n6798), .DIN2(n4233), .Q(WX2557) );
  xor2s3 U2978 ( .DIN1(n6114), .DIN2(n3286), .Q(n4233) );
  nor2s3 U2979 ( .DIN1(n5864), .DIN2(n6762), .Q(WX2191) );
  nor2s3 U2980 ( .DIN1(n5871), .DIN2(n6762), .Q(WX2189) );
  nor2s3 U2981 ( .DIN1(n5878), .DIN2(n6762), .Q(WX2187) );
  nor2s3 U2982 ( .DIN1(n5885), .DIN2(n6762), .Q(WX2185) );
  nor2s3 U2983 ( .DIN1(n5892), .DIN2(n6762), .Q(WX2183) );
  nor2s3 U2984 ( .DIN1(n5899), .DIN2(n6762), .Q(WX2181) );
  nor2s3 U2985 ( .DIN1(n5906), .DIN2(n6762), .Q(WX2179) );
  nor2s3 U2986 ( .DIN1(n5913), .DIN2(n6762), .Q(WX2177) );
  nor2s3 U2987 ( .DIN1(n5920), .DIN2(n6762), .Q(WX2175) );
  nor2s3 U2988 ( .DIN1(n5927), .DIN2(n6762), .Q(WX2173) );
  nor2s3 U2989 ( .DIN1(n5934), .DIN2(n6762), .Q(WX2171) );
  nor2s3 U2990 ( .DIN1(n5941), .DIN2(n6762), .Q(WX2169) );
  nor2s3 U2991 ( .DIN1(n5948), .DIN2(n6761), .Q(WX2167) );
  nor2s3 U2992 ( .DIN1(n5955), .DIN2(n6761), .Q(WX2165) );
  nor2s3 U2993 ( .DIN1(n5962), .DIN2(n6761), .Q(WX2163) );
  nor2s3 U2994 ( .DIN1(n5969), .DIN2(n6761), .Q(WX2161) );
  nor2s3 U2995 ( .DIN1(n5977), .DIN2(n6761), .Q(WX2159) );
  nor2s3 U2996 ( .DIN1(n5986), .DIN2(n6761), .Q(WX2157) );
  nor2s3 U2997 ( .DIN1(n5995), .DIN2(n6761), .Q(WX2155) );
  nor2s3 U2998 ( .DIN1(n6004), .DIN2(n6761), .Q(WX2153) );
  nor2s3 U2999 ( .DIN1(n6013), .DIN2(n6761), .Q(WX2151) );
  nor2s3 U3000 ( .DIN1(n6022), .DIN2(n6761), .Q(WX2149) );
  nor2s3 U3001 ( .DIN1(n6031), .DIN2(n6761), .Q(WX2147) );
  nor2s3 U3002 ( .DIN1(n6040), .DIN2(n6760), .Q(WX2145) );
  nor2s3 U3003 ( .DIN1(n6049), .DIN2(n6760), .Q(WX2143) );
  nor2s3 U3004 ( .DIN1(n6058), .DIN2(n6760), .Q(WX2141) );
  nor2s3 U3005 ( .DIN1(n6067), .DIN2(n6760), .Q(WX2139) );
  nor2s3 U3006 ( .DIN1(n6076), .DIN2(n6760), .Q(WX2137) );
  nor2s3 U3007 ( .DIN1(n6085), .DIN2(n6760), .Q(WX2135) );
  nor2s3 U3008 ( .DIN1(n6094), .DIN2(n6760), .Q(WX2133) );
  nor2s3 U3009 ( .DIN1(n6103), .DIN2(n6760), .Q(WX2131) );
  nor2s3 U3010 ( .DIN1(n6112), .DIN2(n6760), .Q(WX2129) );
  and2s3 U3011 ( .DIN1(RESET), .DIN2(n5863), .Q(WX2127) );
  and2s3 U3012 ( .DIN1(RESET), .DIN2(n5870), .Q(WX2125) );
  and2s3 U3013 ( .DIN1(RESET), .DIN2(n5877), .Q(WX2123) );
  and2s3 U3014 ( .DIN1(RESET), .DIN2(n5884), .Q(WX2121) );
  and2s3 U3015 ( .DIN1(RESET), .DIN2(n5891), .Q(WX2119) );
  and2s3 U3016 ( .DIN1(RESET), .DIN2(n5898), .Q(WX2117) );
  and2s3 U3017 ( .DIN1(RESET), .DIN2(n5905), .Q(WX2115) );
  and2s3 U3018 ( .DIN1(RESET), .DIN2(n5912), .Q(WX2113) );
  and2s3 U3019 ( .DIN1(RESET), .DIN2(n5919), .Q(WX2111) );
  and2s3 U3020 ( .DIN1(RESET), .DIN2(n5926), .Q(WX2109) );
  and2s3 U3021 ( .DIN1(RESET), .DIN2(n5933), .Q(WX2107) );
  and2s3 U3022 ( .DIN1(RESET), .DIN2(n5940), .Q(WX2105) );
  and2s3 U3023 ( .DIN1(RESET), .DIN2(n5947), .Q(WX2103) );
  and2s3 U3024 ( .DIN1(RESET), .DIN2(n5954), .Q(WX2101) );
  and2s3 U3025 ( .DIN1(RESET), .DIN2(n5961), .Q(WX2099) );
  and2s3 U3026 ( .DIN1(RESET), .DIN2(n5968), .Q(WX2097) );
  and2s3 U3027 ( .DIN1(RESET), .DIN2(n5976), .Q(WX2095) );
  and2s3 U3028 ( .DIN1(RESET), .DIN2(n5985), .Q(WX2093) );
  and2s3 U3029 ( .DIN1(RESET), .DIN2(n5994), .Q(WX2091) );
  and2s3 U3030 ( .DIN1(RESET), .DIN2(n6003), .Q(WX2089) );
  and2s3 U3031 ( .DIN1(RESET), .DIN2(n6012), .Q(WX2087) );
  and2s3 U3032 ( .DIN1(RESET), .DIN2(n6021), .Q(WX2085) );
  and2s3 U3033 ( .DIN1(RESET), .DIN2(n6030), .Q(WX2083) );
  and2s3 U3034 ( .DIN1(RESET), .DIN2(n6039), .Q(WX2081) );
  and2s3 U3035 ( .DIN1(RESET), .DIN2(n6048), .Q(WX2079) );
  and2s3 U3036 ( .DIN1(RESET), .DIN2(n6057), .Q(WX2077) );
  and2s3 U3037 ( .DIN1(RESET), .DIN2(n6066), .Q(WX2075) );
  and2s3 U3038 ( .DIN1(RESET), .DIN2(n6075), .Q(WX2073) );
  and2s3 U3039 ( .DIN1(RESET), .DIN2(n6084), .Q(WX2071) );
  and2s3 U3040 ( .DIN1(RESET), .DIN2(n6093), .Q(WX2069) );
  and2s3 U3041 ( .DIN1(RESET), .DIN2(n6102), .Q(WX2067) );
  and2s3 U3042 ( .DIN1(RESET), .DIN2(n6111), .Q(WX2065) );
  nor2s3 U3043 ( .DIN1(n5862), .DIN2(n6760), .Q(WX2063) );
  nor2s3 U3044 ( .DIN1(n5869), .DIN2(n6760), .Q(WX2061) );
  nor2s3 U3045 ( .DIN1(n5876), .DIN2(n6760), .Q(WX2059) );
  nor2s3 U3046 ( .DIN1(n5883), .DIN2(n6759), .Q(WX2057) );
  nor2s3 U3047 ( .DIN1(n5890), .DIN2(n6759), .Q(WX2055) );
  nor2s3 U3048 ( .DIN1(n5897), .DIN2(n6759), .Q(WX2053) );
  nor2s3 U3049 ( .DIN1(n5904), .DIN2(n6759), .Q(WX2051) );
  nor2s3 U3050 ( .DIN1(n5911), .DIN2(n6759), .Q(WX2049) );
  nor2s3 U3051 ( .DIN1(n5918), .DIN2(n6759), .Q(WX2047) );
  nor2s3 U3052 ( .DIN1(n5925), .DIN2(n6759), .Q(WX2045) );
  nor2s3 U3053 ( .DIN1(n5932), .DIN2(n6759), .Q(WX2043) );
  nor2s3 U3054 ( .DIN1(n5939), .DIN2(n6759), .Q(WX2041) );
  nor2s3 U3055 ( .DIN1(n5946), .DIN2(n6759), .Q(WX2039) );
  nor2s3 U3056 ( .DIN1(n5953), .DIN2(n6759), .Q(WX2037) );
  nor2s3 U3057 ( .DIN1(n5960), .DIN2(n6759), .Q(WX2035) );
  nor2s3 U3058 ( .DIN1(n5967), .DIN2(n6758), .Q(WX2033) );
  nor2s3 U3059 ( .DIN1(n5975), .DIN2(n6758), .Q(WX2031) );
  nor2s3 U3060 ( .DIN1(n5984), .DIN2(n6758), .Q(WX2029) );
  nor2s3 U3061 ( .DIN1(n5993), .DIN2(n6758), .Q(WX2027) );
  nor2s3 U3062 ( .DIN1(n6002), .DIN2(n6758), .Q(WX2025) );
  nor2s3 U3063 ( .DIN1(n6011), .DIN2(n6758), .Q(WX2023) );
  nor2s3 U3064 ( .DIN1(n6020), .DIN2(n6758), .Q(WX2021) );
  nor2s3 U3065 ( .DIN1(n6029), .DIN2(n6758), .Q(WX2019) );
  nor2s3 U3066 ( .DIN1(n6038), .DIN2(n6758), .Q(WX2017) );
  nor2s3 U3067 ( .DIN1(n6047), .DIN2(n6758), .Q(WX2015) );
  nor2s3 U3068 ( .DIN1(n6056), .DIN2(n6758), .Q(WX2013) );
  nor2s3 U3069 ( .DIN1(n6065), .DIN2(n6758), .Q(WX2011) );
  nor2s3 U3070 ( .DIN1(n6074), .DIN2(n6757), .Q(WX2009) );
  nor2s3 U3071 ( .DIN1(n6083), .DIN2(n6757), .Q(WX2007) );
  nor2s3 U3072 ( .DIN1(n6092), .DIN2(n6757), .Q(WX2005) );
  nor2s3 U3073 ( .DIN1(n6101), .DIN2(n6757), .Q(WX2003) );
  nor2s3 U3074 ( .DIN1(n6110), .DIN2(n6757), .Q(WX2001) );
  nnd4s2 U3075 ( .DIN1(n4234), .DIN2(n4235), .DIN3(n4236), .DIN4(n4237), .Q(
        WX1999) );
  nnd2s3 U3076 ( .DIN1(n3965), .DIN2(n6640), .Q(n4237) );
  xor2s3 U3077 ( .DIN1(n4238), .DIN2(n4239), .Q(n3965) );
  xor2s3 U3078 ( .DIN1(n5859), .DIN2(n5860), .Q(n4239) );
  xnr2s3 U3079 ( .DIN1(n3285), .DIN2(n5861), .Q(n4238) );
  nnd2s3 U3080 ( .DIN1(n3058), .DIN2(n6671), .Q(n4236) );
  xor2s3 U3081 ( .DIN1(n4240), .DIN2(n4241), .Q(n3058) );
  xor2s3 U3082 ( .DIN1(n5862), .DIN2(n5863), .Q(n4241) );
  xnr2s3 U3083 ( .DIN1(n3286), .DIN2(n5864), .Q(n4240) );
  nnd2s3 U3084 ( .DIN1(n6598), .DIN2(n2209), .Q(n4235) );
  nnd2s3 U3085 ( .DIN1(n6567), .DIN2(n2208), .Q(n4234) );
  nnd4s2 U3086 ( .DIN1(n4242), .DIN2(n4243), .DIN3(n4244), .DIN4(n4245), .Q(
        WX1997) );
  nnd2s3 U3087 ( .DIN1(n3972), .DIN2(n6640), .Q(n4245) );
  xor2s3 U3088 ( .DIN1(n4246), .DIN2(n4247), .Q(n3972) );
  xor2s3 U3089 ( .DIN1(n5866), .DIN2(n5867), .Q(n4247) );
  xnr2s3 U3090 ( .DIN1(n3287), .DIN2(n5868), .Q(n4246) );
  nnd2s3 U3091 ( .DIN1(n3064), .DIN2(n6671), .Q(n4244) );
  xor2s3 U3092 ( .DIN1(n4248), .DIN2(n4249), .Q(n3064) );
  xor2s3 U3093 ( .DIN1(n5869), .DIN2(n5870), .Q(n4249) );
  xnr2s3 U3094 ( .DIN1(n3288), .DIN2(n5871), .Q(n4248) );
  nnd2s3 U3095 ( .DIN1(n6598), .DIN2(n2210), .Q(n4243) );
  nnd2s3 U3096 ( .DIN1(n6567), .DIN2(n2207), .Q(n4242) );
  nnd4s2 U3097 ( .DIN1(n4250), .DIN2(n4251), .DIN3(n4252), .DIN4(n4253), .Q(
        WX1995) );
  nnd2s3 U3098 ( .DIN1(n3979), .DIN2(n6640), .Q(n4253) );
  xor2s3 U3099 ( .DIN1(n4254), .DIN2(n4255), .Q(n3979) );
  xor2s3 U3100 ( .DIN1(n5873), .DIN2(n5874), .Q(n4255) );
  xnr2s3 U3101 ( .DIN1(n3289), .DIN2(n5875), .Q(n4254) );
  nnd2s3 U3102 ( .DIN1(n3070), .DIN2(n6671), .Q(n4252) );
  xor2s3 U3103 ( .DIN1(n4256), .DIN2(n4257), .Q(n3070) );
  xor2s3 U3104 ( .DIN1(n5876), .DIN2(n5877), .Q(n4257) );
  xnr2s3 U3105 ( .DIN1(n3290), .DIN2(n5878), .Q(n4256) );
  nnd2s3 U3106 ( .DIN1(n6598), .DIN2(n2211), .Q(n4251) );
  nnd2s3 U3107 ( .DIN1(n6567), .DIN2(n2206), .Q(n4250) );
  nnd4s2 U3108 ( .DIN1(n4258), .DIN2(n4259), .DIN3(n4260), .DIN4(n4261), .Q(
        WX1993) );
  nnd2s3 U3109 ( .DIN1(n3986), .DIN2(n6640), .Q(n4261) );
  xor2s3 U3110 ( .DIN1(n4262), .DIN2(n4263), .Q(n3986) );
  xor2s3 U3111 ( .DIN1(n5880), .DIN2(n5881), .Q(n4263) );
  xnr2s3 U3112 ( .DIN1(n3291), .DIN2(n5882), .Q(n4262) );
  nnd2s3 U3113 ( .DIN1(n3076), .DIN2(n6671), .Q(n4260) );
  xor2s3 U3114 ( .DIN1(n4264), .DIN2(n4265), .Q(n3076) );
  xor2s3 U3115 ( .DIN1(n5883), .DIN2(n5884), .Q(n4265) );
  xnr2s3 U3116 ( .DIN1(n3292), .DIN2(n5885), .Q(n4264) );
  nnd2s3 U3117 ( .DIN1(n6598), .DIN2(n2212), .Q(n4259) );
  nnd2s3 U3118 ( .DIN1(n6567), .DIN2(n2205), .Q(n4258) );
  nnd4s2 U3119 ( .DIN1(n4266), .DIN2(n4267), .DIN3(n4268), .DIN4(n4269), .Q(
        WX1991) );
  nnd2s3 U3120 ( .DIN1(n3993), .DIN2(n6640), .Q(n4269) );
  xor2s3 U3121 ( .DIN1(n4270), .DIN2(n4271), .Q(n3993) );
  xor2s3 U3122 ( .DIN1(n5887), .DIN2(n5888), .Q(n4271) );
  xnr2s3 U3123 ( .DIN1(n3293), .DIN2(n5889), .Q(n4270) );
  nnd2s3 U3124 ( .DIN1(n3082), .DIN2(n6671), .Q(n4268) );
  xor2s3 U3125 ( .DIN1(n4272), .DIN2(n4273), .Q(n3082) );
  xor2s3 U3126 ( .DIN1(n5890), .DIN2(n5891), .Q(n4273) );
  xnr2s3 U3127 ( .DIN1(n3294), .DIN2(n5892), .Q(n4272) );
  nnd2s3 U3128 ( .DIN1(n6598), .DIN2(n2213), .Q(n4267) );
  nnd2s3 U3129 ( .DIN1(n6567), .DIN2(n2204), .Q(n4266) );
  nnd4s2 U3130 ( .DIN1(n4274), .DIN2(n4275), .DIN3(n4276), .DIN4(n4277), .Q(
        WX1989) );
  nnd2s3 U3131 ( .DIN1(n4000), .DIN2(n6640), .Q(n4277) );
  xor2s3 U3132 ( .DIN1(n4278), .DIN2(n4279), .Q(n4000) );
  xor2s3 U3133 ( .DIN1(n5894), .DIN2(n5895), .Q(n4279) );
  xnr2s3 U3134 ( .DIN1(n3295), .DIN2(n5896), .Q(n4278) );
  nnd2s3 U3135 ( .DIN1(n3088), .DIN2(n6671), .Q(n4276) );
  xor2s3 U3136 ( .DIN1(n4280), .DIN2(n4281), .Q(n3088) );
  xor2s3 U3137 ( .DIN1(n5897), .DIN2(n5898), .Q(n4281) );
  xnr2s3 U3138 ( .DIN1(n3296), .DIN2(n5899), .Q(n4280) );
  nnd2s3 U3139 ( .DIN1(n6598), .DIN2(n2214), .Q(n4275) );
  nnd2s3 U3140 ( .DIN1(n6567), .DIN2(n2203), .Q(n4274) );
  nnd4s2 U3141 ( .DIN1(n4282), .DIN2(n4283), .DIN3(n4284), .DIN4(n4285), .Q(
        WX1987) );
  nnd2s3 U3142 ( .DIN1(n4007), .DIN2(n6640), .Q(n4285) );
  xor2s3 U3143 ( .DIN1(n4286), .DIN2(n4287), .Q(n4007) );
  xor2s3 U3144 ( .DIN1(n5901), .DIN2(n5902), .Q(n4287) );
  xnr2s3 U3145 ( .DIN1(n3297), .DIN2(n5903), .Q(n4286) );
  nnd2s3 U3146 ( .DIN1(n3094), .DIN2(n6671), .Q(n4284) );
  xor2s3 U3147 ( .DIN1(n4288), .DIN2(n4289), .Q(n3094) );
  xor2s3 U3148 ( .DIN1(n5904), .DIN2(n5905), .Q(n4289) );
  xnr2s3 U3149 ( .DIN1(n3298), .DIN2(n5906), .Q(n4288) );
  nnd2s3 U3150 ( .DIN1(n6598), .DIN2(n2215), .Q(n4283) );
  nnd2s3 U3151 ( .DIN1(n6567), .DIN2(n2202), .Q(n4282) );
  nnd4s2 U3152 ( .DIN1(n4290), .DIN2(n4291), .DIN3(n4292), .DIN4(n4293), .Q(
        WX1985) );
  nnd2s3 U3153 ( .DIN1(n4014), .DIN2(n6640), .Q(n4293) );
  xor2s3 U3154 ( .DIN1(n4294), .DIN2(n4295), .Q(n4014) );
  xor2s3 U3155 ( .DIN1(n5908), .DIN2(n5909), .Q(n4295) );
  xnr2s3 U3156 ( .DIN1(n3299), .DIN2(n5910), .Q(n4294) );
  nnd2s3 U3157 ( .DIN1(n3100), .DIN2(n6671), .Q(n4292) );
  xor2s3 U3158 ( .DIN1(n4296), .DIN2(n4297), .Q(n3100) );
  xor2s3 U3159 ( .DIN1(n5911), .DIN2(n5912), .Q(n4297) );
  xnr2s3 U3160 ( .DIN1(n3300), .DIN2(n5913), .Q(n4296) );
  nnd2s3 U3161 ( .DIN1(n6598), .DIN2(n2216), .Q(n4291) );
  nnd2s3 U3162 ( .DIN1(n6567), .DIN2(n2201), .Q(n4290) );
  nnd4s2 U3163 ( .DIN1(n4298), .DIN2(n4299), .DIN3(n4300), .DIN4(n4301), .Q(
        WX1983) );
  nnd2s3 U3164 ( .DIN1(n4021), .DIN2(n6640), .Q(n4301) );
  xor2s3 U3165 ( .DIN1(n4302), .DIN2(n4303), .Q(n4021) );
  xor2s3 U3166 ( .DIN1(n5915), .DIN2(n5916), .Q(n4303) );
  xnr2s3 U3167 ( .DIN1(n3301), .DIN2(n5917), .Q(n4302) );
  nnd2s3 U3168 ( .DIN1(n3106), .DIN2(n6671), .Q(n4300) );
  xor2s3 U3169 ( .DIN1(n4304), .DIN2(n4305), .Q(n3106) );
  xor2s3 U3170 ( .DIN1(n5918), .DIN2(n5919), .Q(n4305) );
  xnr2s3 U3171 ( .DIN1(n3302), .DIN2(n5920), .Q(n4304) );
  nnd2s3 U3172 ( .DIN1(n6598), .DIN2(n2217), .Q(n4299) );
  nnd2s3 U3173 ( .DIN1(n6567), .DIN2(n2200), .Q(n4298) );
  nnd4s2 U3174 ( .DIN1(n4306), .DIN2(n4307), .DIN3(n4308), .DIN4(n4309), .Q(
        WX1981) );
  nnd2s3 U3175 ( .DIN1(n4028), .DIN2(n6640), .Q(n4309) );
  xor2s3 U3176 ( .DIN1(n4310), .DIN2(n4311), .Q(n4028) );
  xor2s3 U3177 ( .DIN1(n5922), .DIN2(n5923), .Q(n4311) );
  xnr2s3 U3178 ( .DIN1(n3303), .DIN2(n5924), .Q(n4310) );
  nnd2s3 U3179 ( .DIN1(n3112), .DIN2(n6671), .Q(n4308) );
  xor2s3 U3180 ( .DIN1(n4312), .DIN2(n4313), .Q(n3112) );
  xor2s3 U3181 ( .DIN1(n5925), .DIN2(n5926), .Q(n4313) );
  xnr2s3 U3182 ( .DIN1(n3304), .DIN2(n5927), .Q(n4312) );
  nnd2s3 U3183 ( .DIN1(n6598), .DIN2(n2218), .Q(n4307) );
  nnd2s3 U3184 ( .DIN1(n6567), .DIN2(n2199), .Q(n4306) );
  nnd4s2 U3185 ( .DIN1(n4314), .DIN2(n4315), .DIN3(n4316), .DIN4(n4317), .Q(
        WX1979) );
  nnd2s3 U3186 ( .DIN1(n4035), .DIN2(n6640), .Q(n4317) );
  xor2s3 U3187 ( .DIN1(n4318), .DIN2(n4319), .Q(n4035) );
  xor2s3 U3188 ( .DIN1(n5929), .DIN2(n5930), .Q(n4319) );
  xnr2s3 U3189 ( .DIN1(n3305), .DIN2(n5931), .Q(n4318) );
  nnd2s3 U3190 ( .DIN1(n3118), .DIN2(n6671), .Q(n4316) );
  xor2s3 U3191 ( .DIN1(n4320), .DIN2(n4321), .Q(n3118) );
  xor2s3 U3192 ( .DIN1(n5932), .DIN2(n5933), .Q(n4321) );
  xnr2s3 U3193 ( .DIN1(n3306), .DIN2(n5934), .Q(n4320) );
  nnd2s3 U3194 ( .DIN1(n6598), .DIN2(n2219), .Q(n4315) );
  nnd2s3 U3195 ( .DIN1(n6567), .DIN2(n2198), .Q(n4314) );
  nnd4s2 U3196 ( .DIN1(n4322), .DIN2(n4323), .DIN3(n4324), .DIN4(n4325), .Q(
        WX1977) );
  nnd2s3 U3197 ( .DIN1(n4042), .DIN2(n6640), .Q(n4325) );
  xor2s3 U3198 ( .DIN1(n4326), .DIN2(n4327), .Q(n4042) );
  xor2s3 U3199 ( .DIN1(n5936), .DIN2(n5937), .Q(n4327) );
  xnr2s3 U3200 ( .DIN1(n3307), .DIN2(n5938), .Q(n4326) );
  nnd2s3 U3201 ( .DIN1(n3124), .DIN2(n6671), .Q(n4324) );
  xor2s3 U3202 ( .DIN1(n4328), .DIN2(n4329), .Q(n3124) );
  xor2s3 U3203 ( .DIN1(n5939), .DIN2(n5940), .Q(n4329) );
  xnr2s3 U3204 ( .DIN1(n3308), .DIN2(n5941), .Q(n4328) );
  nnd2s3 U3205 ( .DIN1(n6598), .DIN2(n2220), .Q(n4323) );
  nnd2s3 U3206 ( .DIN1(n6567), .DIN2(n2197), .Q(n4322) );
  nnd4s2 U3207 ( .DIN1(n4330), .DIN2(n4331), .DIN3(n4332), .DIN4(n4333), .Q(
        WX1975) );
  nnd2s3 U3208 ( .DIN1(n4049), .DIN2(n6639), .Q(n4333) );
  xor2s3 U3209 ( .DIN1(n4334), .DIN2(n4335), .Q(n4049) );
  xor2s3 U3210 ( .DIN1(n5943), .DIN2(n5944), .Q(n4335) );
  xnr2s3 U3211 ( .DIN1(n3309), .DIN2(n5945), .Q(n4334) );
  nnd2s3 U3212 ( .DIN1(n3130), .DIN2(n6670), .Q(n4332) );
  xor2s3 U3213 ( .DIN1(n4336), .DIN2(n4337), .Q(n3130) );
  xor2s3 U3214 ( .DIN1(n5946), .DIN2(n5947), .Q(n4337) );
  xnr2s3 U3215 ( .DIN1(n3310), .DIN2(n5948), .Q(n4336) );
  nnd2s3 U3216 ( .DIN1(n6597), .DIN2(n2221), .Q(n4331) );
  nnd2s3 U3217 ( .DIN1(n6566), .DIN2(n2196), .Q(n4330) );
  nnd4s2 U3218 ( .DIN1(n4338), .DIN2(n4339), .DIN3(n4340), .DIN4(n4341), .Q(
        WX1973) );
  nnd2s3 U3219 ( .DIN1(n4056), .DIN2(n6639), .Q(n4341) );
  xor2s3 U3220 ( .DIN1(n4342), .DIN2(n4343), .Q(n4056) );
  xor2s3 U3221 ( .DIN1(n5950), .DIN2(n5951), .Q(n4343) );
  xnr2s3 U3222 ( .DIN1(n3311), .DIN2(n5952), .Q(n4342) );
  nnd2s3 U3223 ( .DIN1(n3136), .DIN2(n6670), .Q(n4340) );
  xor2s3 U3224 ( .DIN1(n4344), .DIN2(n4345), .Q(n3136) );
  xor2s3 U3225 ( .DIN1(n5953), .DIN2(n5954), .Q(n4345) );
  xnr2s3 U3226 ( .DIN1(n3312), .DIN2(n5955), .Q(n4344) );
  nnd2s3 U3227 ( .DIN1(n6597), .DIN2(n2222), .Q(n4339) );
  nnd2s3 U3228 ( .DIN1(n6566), .DIN2(n2195), .Q(n4338) );
  nnd4s2 U3229 ( .DIN1(n4346), .DIN2(n4347), .DIN3(n4348), .DIN4(n4349), .Q(
        WX1971) );
  nnd2s3 U3230 ( .DIN1(n4063), .DIN2(n6639), .Q(n4349) );
  xor2s3 U3231 ( .DIN1(n4350), .DIN2(n4351), .Q(n4063) );
  xor2s3 U3232 ( .DIN1(n5957), .DIN2(n5958), .Q(n4351) );
  xnr2s3 U3233 ( .DIN1(n3313), .DIN2(n5959), .Q(n4350) );
  nnd2s3 U3234 ( .DIN1(n3142), .DIN2(n6670), .Q(n4348) );
  xor2s3 U3235 ( .DIN1(n4352), .DIN2(n4353), .Q(n3142) );
  xor2s3 U3236 ( .DIN1(n5960), .DIN2(n5961), .Q(n4353) );
  xnr2s3 U3237 ( .DIN1(n3314), .DIN2(n5962), .Q(n4352) );
  nnd2s3 U3238 ( .DIN1(n6597), .DIN2(n2223), .Q(n4347) );
  nnd2s3 U3239 ( .DIN1(n6566), .DIN2(n2194), .Q(n4346) );
  nnd4s2 U3240 ( .DIN1(n4354), .DIN2(n4355), .DIN3(n4356), .DIN4(n4357), .Q(
        WX1969) );
  nnd2s3 U3241 ( .DIN1(n4070), .DIN2(n6639), .Q(n4357) );
  xor2s3 U3242 ( .DIN1(n4358), .DIN2(n4359), .Q(n4070) );
  xor2s3 U3243 ( .DIN1(n5964), .DIN2(n5965), .Q(n4359) );
  xnr2s3 U3244 ( .DIN1(n3315), .DIN2(n5966), .Q(n4358) );
  nnd2s3 U3245 ( .DIN1(n3148), .DIN2(n6670), .Q(n4356) );
  xor2s3 U3246 ( .DIN1(n4360), .DIN2(n4361), .Q(n3148) );
  xor2s3 U3247 ( .DIN1(n5967), .DIN2(n5968), .Q(n4361) );
  xnr2s3 U3248 ( .DIN1(n3316), .DIN2(n5969), .Q(n4360) );
  nnd2s3 U3249 ( .DIN1(n6597), .DIN2(n2224), .Q(n4355) );
  nnd2s3 U3250 ( .DIN1(n6566), .DIN2(n2193), .Q(n4354) );
  nnd4s2 U3251 ( .DIN1(n4362), .DIN2(n4363), .DIN3(n4364), .DIN4(n4365), .Q(
        WX1967) );
  nnd2s3 U3252 ( .DIN1(n4078), .DIN2(n6639), .Q(n4365) );
  xor2s3 U3253 ( .DIN1(n4366), .DIN2(n4367), .Q(n4078) );
  xor2s3 U3254 ( .DIN1(n5973), .DIN2(n4368), .Q(n4367) );
  xor2s3 U3255 ( .DIN1(n5971), .DIN2(n5972), .Q(n4368) );
  xor2s3 U3256 ( .DIN1(n5974), .DIN2(n6693), .Q(n4366) );
  nnd2s3 U3257 ( .DIN1(n3154), .DIN2(n6670), .Q(n4364) );
  xor2s3 U3258 ( .DIN1(n4369), .DIN2(n4370), .Q(n3154) );
  xor2s3 U3259 ( .DIN1(n5977), .DIN2(n4371), .Q(n4370) );
  xor2s3 U3260 ( .DIN1(n5975), .DIN2(n5976), .Q(n4371) );
  xor2s3 U3261 ( .DIN1(n5978), .DIN2(n6693), .Q(n4369) );
  nnd2s3 U3262 ( .DIN1(n6597), .DIN2(n2225), .Q(n4363) );
  nnd2s3 U3263 ( .DIN1(n6566), .DIN2(n2192), .Q(n4362) );
  nnd4s2 U3264 ( .DIN1(n4372), .DIN2(n4373), .DIN3(n4374), .DIN4(n4375), .Q(
        WX1965) );
  nnd2s3 U3265 ( .DIN1(n4086), .DIN2(n6639), .Q(n4375) );
  xor2s3 U3266 ( .DIN1(n4376), .DIN2(n4377), .Q(n4086) );
  xor2s3 U3267 ( .DIN1(n5982), .DIN2(n4378), .Q(n4377) );
  xor2s3 U3268 ( .DIN1(n5980), .DIN2(n5981), .Q(n4378) );
  xor2s3 U3269 ( .DIN1(n5983), .DIN2(n6693), .Q(n4376) );
  nnd2s3 U3270 ( .DIN1(n3160), .DIN2(n6670), .Q(n4374) );
  xor2s3 U3271 ( .DIN1(n4379), .DIN2(n4380), .Q(n3160) );
  xor2s3 U3272 ( .DIN1(n5986), .DIN2(n4381), .Q(n4380) );
  xor2s3 U3273 ( .DIN1(n5984), .DIN2(n5985), .Q(n4381) );
  xor2s3 U3274 ( .DIN1(n5987), .DIN2(n6693), .Q(n4379) );
  nnd2s3 U3275 ( .DIN1(n6597), .DIN2(n2226), .Q(n4373) );
  nnd2s3 U3276 ( .DIN1(n6566), .DIN2(n2191), .Q(n4372) );
  nnd4s2 U3277 ( .DIN1(n4382), .DIN2(n4383), .DIN3(n4384), .DIN4(n4385), .Q(
        WX1963) );
  nnd2s3 U3278 ( .DIN1(n4094), .DIN2(n6639), .Q(n4385) );
  xor2s3 U3279 ( .DIN1(n4386), .DIN2(n4387), .Q(n4094) );
  xor2s3 U3280 ( .DIN1(n5991), .DIN2(n4388), .Q(n4387) );
  xor2s3 U3281 ( .DIN1(n5989), .DIN2(n5990), .Q(n4388) );
  xor2s3 U3282 ( .DIN1(n5992), .DIN2(n6693), .Q(n4386) );
  nnd2s3 U3283 ( .DIN1(n3166), .DIN2(n6670), .Q(n4384) );
  xor2s3 U3284 ( .DIN1(n4389), .DIN2(n4390), .Q(n3166) );
  xor2s3 U3285 ( .DIN1(n5995), .DIN2(n4391), .Q(n4390) );
  xor2s3 U3286 ( .DIN1(n5993), .DIN2(n5994), .Q(n4391) );
  xor2s3 U3287 ( .DIN1(n5996), .DIN2(n6693), .Q(n4389) );
  nnd2s3 U3288 ( .DIN1(n6597), .DIN2(n2227), .Q(n4383) );
  nnd2s3 U3289 ( .DIN1(n6566), .DIN2(n2190), .Q(n4382) );
  nnd4s2 U3290 ( .DIN1(n4392), .DIN2(n4393), .DIN3(n4394), .DIN4(n4395), .Q(
        WX1961) );
  nnd2s3 U3291 ( .DIN1(n4102), .DIN2(n6639), .Q(n4395) );
  xor2s3 U3292 ( .DIN1(n4396), .DIN2(n4397), .Q(n4102) );
  xor2s3 U3293 ( .DIN1(n6000), .DIN2(n4398), .Q(n4397) );
  xor2s3 U3294 ( .DIN1(n5998), .DIN2(n5999), .Q(n4398) );
  xor2s3 U3295 ( .DIN1(n6001), .DIN2(n6693), .Q(n4396) );
  nnd2s3 U3296 ( .DIN1(n3172), .DIN2(n6670), .Q(n4394) );
  xor2s3 U3297 ( .DIN1(n4399), .DIN2(n4400), .Q(n3172) );
  xor2s3 U3298 ( .DIN1(n6004), .DIN2(n4401), .Q(n4400) );
  xor2s3 U3299 ( .DIN1(n6002), .DIN2(n6003), .Q(n4401) );
  xor2s3 U3300 ( .DIN1(n6005), .DIN2(n6693), .Q(n4399) );
  nnd2s3 U3301 ( .DIN1(n6597), .DIN2(n2228), .Q(n4393) );
  nnd2s3 U3302 ( .DIN1(n6566), .DIN2(n2189), .Q(n4392) );
  nnd4s2 U3303 ( .DIN1(n4402), .DIN2(n4403), .DIN3(n4404), .DIN4(n4405), .Q(
        WX1959) );
  nnd2s3 U3304 ( .DIN1(n4110), .DIN2(n6639), .Q(n4405) );
  xor2s3 U3305 ( .DIN1(n4406), .DIN2(n4407), .Q(n4110) );
  xor2s3 U3306 ( .DIN1(n6009), .DIN2(n4408), .Q(n4407) );
  xor2s3 U3307 ( .DIN1(n6007), .DIN2(n6008), .Q(n4408) );
  xor2s3 U3308 ( .DIN1(n6010), .DIN2(n6693), .Q(n4406) );
  nnd2s3 U3309 ( .DIN1(n3178), .DIN2(n6670), .Q(n4404) );
  xor2s3 U3310 ( .DIN1(n4409), .DIN2(n4410), .Q(n3178) );
  xor2s3 U3311 ( .DIN1(n6013), .DIN2(n4411), .Q(n4410) );
  xor2s3 U3312 ( .DIN1(n6011), .DIN2(n6012), .Q(n4411) );
  xor2s3 U3313 ( .DIN1(n6014), .DIN2(n6693), .Q(n4409) );
  nnd2s3 U3314 ( .DIN1(n6597), .DIN2(n2229), .Q(n4403) );
  nnd2s3 U3315 ( .DIN1(n6566), .DIN2(n2188), .Q(n4402) );
  nnd4s2 U3316 ( .DIN1(n4412), .DIN2(n4413), .DIN3(n4414), .DIN4(n4415), .Q(
        WX1957) );
  nnd2s3 U3317 ( .DIN1(n4118), .DIN2(n6639), .Q(n4415) );
  xor2s3 U3318 ( .DIN1(n4416), .DIN2(n4417), .Q(n4118) );
  xor2s3 U3319 ( .DIN1(n6018), .DIN2(n4418), .Q(n4417) );
  xor2s3 U3320 ( .DIN1(n6016), .DIN2(n6017), .Q(n4418) );
  xor2s3 U3321 ( .DIN1(n6019), .DIN2(n6694), .Q(n4416) );
  nnd2s3 U3322 ( .DIN1(n3184), .DIN2(n6670), .Q(n4414) );
  xor2s3 U3323 ( .DIN1(n4419), .DIN2(n4420), .Q(n3184) );
  xor2s3 U3324 ( .DIN1(n6022), .DIN2(n4421), .Q(n4420) );
  xor2s3 U3325 ( .DIN1(n6020), .DIN2(n6021), .Q(n4421) );
  xor2s3 U3326 ( .DIN1(n6023), .DIN2(n6694), .Q(n4419) );
  nnd2s3 U3327 ( .DIN1(n6597), .DIN2(n2230), .Q(n4413) );
  nnd2s3 U3328 ( .DIN1(n6566), .DIN2(n2187), .Q(n4412) );
  nnd4s2 U3329 ( .DIN1(n4422), .DIN2(n4423), .DIN3(n4424), .DIN4(n4425), .Q(
        WX1955) );
  nnd2s3 U3330 ( .DIN1(n4126), .DIN2(n6639), .Q(n4425) );
  xor2s3 U3331 ( .DIN1(n4426), .DIN2(n4427), .Q(n4126) );
  xor2s3 U3332 ( .DIN1(n6027), .DIN2(n4428), .Q(n4427) );
  xor2s3 U3333 ( .DIN1(n6025), .DIN2(n6026), .Q(n4428) );
  xor2s3 U3334 ( .DIN1(n6028), .DIN2(n6694), .Q(n4426) );
  nnd2s3 U3335 ( .DIN1(n3190), .DIN2(n6670), .Q(n4424) );
  xor2s3 U3336 ( .DIN1(n4429), .DIN2(n4430), .Q(n3190) );
  xor2s3 U3337 ( .DIN1(n6031), .DIN2(n4431), .Q(n4430) );
  xor2s3 U3338 ( .DIN1(n6029), .DIN2(n6030), .Q(n4431) );
  xor2s3 U3339 ( .DIN1(n6032), .DIN2(n6694), .Q(n4429) );
  nnd2s3 U3340 ( .DIN1(n6597), .DIN2(n2231), .Q(n4423) );
  nnd2s3 U3341 ( .DIN1(n6566), .DIN2(n2186), .Q(n4422) );
  nnd4s2 U3342 ( .DIN1(n4432), .DIN2(n4433), .DIN3(n4434), .DIN4(n4435), .Q(
        WX1953) );
  nnd2s3 U3343 ( .DIN1(n4134), .DIN2(n6639), .Q(n4435) );
  xor2s3 U3344 ( .DIN1(n4436), .DIN2(n4437), .Q(n4134) );
  xor2s3 U3345 ( .DIN1(n6036), .DIN2(n4438), .Q(n4437) );
  xor2s3 U3346 ( .DIN1(n6034), .DIN2(n6035), .Q(n4438) );
  xor2s3 U3347 ( .DIN1(n6037), .DIN2(n6694), .Q(n4436) );
  nnd2s3 U3348 ( .DIN1(n3196), .DIN2(n6670), .Q(n4434) );
  xor2s3 U3349 ( .DIN1(n4439), .DIN2(n4440), .Q(n3196) );
  xor2s3 U3350 ( .DIN1(n6040), .DIN2(n4441), .Q(n4440) );
  xor2s3 U3351 ( .DIN1(n6038), .DIN2(n6039), .Q(n4441) );
  xor2s3 U3352 ( .DIN1(n6041), .DIN2(n6694), .Q(n4439) );
  nnd2s3 U3353 ( .DIN1(n6597), .DIN2(n2232), .Q(n4433) );
  nnd2s3 U3354 ( .DIN1(n6566), .DIN2(n2185), .Q(n4432) );
  nnd4s2 U3355 ( .DIN1(n4442), .DIN2(n4443), .DIN3(n4444), .DIN4(n4445), .Q(
        WX1951) );
  nnd2s3 U3356 ( .DIN1(n4142), .DIN2(n6639), .Q(n4445) );
  xor2s3 U3357 ( .DIN1(n4446), .DIN2(n4447), .Q(n4142) );
  xor2s3 U3358 ( .DIN1(n6045), .DIN2(n4448), .Q(n4447) );
  xor2s3 U3359 ( .DIN1(n6043), .DIN2(n6044), .Q(n4448) );
  xor2s3 U3360 ( .DIN1(n6046), .DIN2(n6694), .Q(n4446) );
  nnd2s3 U3361 ( .DIN1(n3202), .DIN2(n6670), .Q(n4444) );
  xor2s3 U3362 ( .DIN1(n4449), .DIN2(n4450), .Q(n3202) );
  xor2s3 U3363 ( .DIN1(n6049), .DIN2(n4451), .Q(n4450) );
  xor2s3 U3364 ( .DIN1(n6047), .DIN2(n6048), .Q(n4451) );
  xor2s3 U3365 ( .DIN1(n6050), .DIN2(n6694), .Q(n4449) );
  nnd2s3 U3366 ( .DIN1(n6597), .DIN2(n2233), .Q(n4443) );
  nnd2s3 U3367 ( .DIN1(n6566), .DIN2(n2184), .Q(n4442) );
  nnd4s2 U3368 ( .DIN1(n4452), .DIN2(n4453), .DIN3(n4454), .DIN4(n4455), .Q(
        WX1949) );
  nnd2s3 U3369 ( .DIN1(n4150), .DIN2(n6638), .Q(n4455) );
  xor2s3 U3370 ( .DIN1(n4456), .DIN2(n4457), .Q(n4150) );
  xor2s3 U3371 ( .DIN1(n6054), .DIN2(n4458), .Q(n4457) );
  xor2s3 U3372 ( .DIN1(n6052), .DIN2(n6053), .Q(n4458) );
  xor2s3 U3373 ( .DIN1(n6055), .DIN2(n6694), .Q(n4456) );
  nnd2s3 U3374 ( .DIN1(n3336), .DIN2(n6669), .Q(n4454) );
  xor2s3 U3375 ( .DIN1(n4459), .DIN2(n4460), .Q(n3336) );
  xor2s3 U3376 ( .DIN1(n6058), .DIN2(n4461), .Q(n4460) );
  xor2s3 U3377 ( .DIN1(n6056), .DIN2(n6057), .Q(n4461) );
  xor2s3 U3378 ( .DIN1(n6059), .DIN2(n6694), .Q(n4459) );
  nnd2s3 U3379 ( .DIN1(n6596), .DIN2(n2234), .Q(n4453) );
  nnd2s3 U3380 ( .DIN1(n6565), .DIN2(n2183), .Q(n4452) );
  nnd4s2 U3381 ( .DIN1(n4462), .DIN2(n4463), .DIN3(n4464), .DIN4(n4465), .Q(
        WX1947) );
  nnd2s3 U3382 ( .DIN1(n4158), .DIN2(n6638), .Q(n4465) );
  xor2s3 U3383 ( .DIN1(n4466), .DIN2(n4467), .Q(n4158) );
  xor2s3 U3384 ( .DIN1(n6063), .DIN2(n4468), .Q(n4467) );
  xor2s3 U3385 ( .DIN1(n6061), .DIN2(n6062), .Q(n4468) );
  xor2s3 U3386 ( .DIN1(n6064), .DIN2(n6694), .Q(n4466) );
  nnd2s3 U3387 ( .DIN1(n3342), .DIN2(n6669), .Q(n4464) );
  xor2s3 U3388 ( .DIN1(n4469), .DIN2(n4470), .Q(n3342) );
  xor2s3 U3389 ( .DIN1(n6067), .DIN2(n4471), .Q(n4470) );
  xor2s3 U3390 ( .DIN1(n6065), .DIN2(n6066), .Q(n4471) );
  xor2s3 U3391 ( .DIN1(n6068), .DIN2(n6694), .Q(n4469) );
  nnd2s3 U3392 ( .DIN1(n6596), .DIN2(n2235), .Q(n4463) );
  nnd2s3 U3393 ( .DIN1(n6565), .DIN2(n2182), .Q(n4462) );
  nnd4s2 U3394 ( .DIN1(n4472), .DIN2(n4473), .DIN3(n4474), .DIN4(n4475), .Q(
        WX1945) );
  nnd2s3 U3395 ( .DIN1(n4166), .DIN2(n6638), .Q(n4475) );
  xor2s3 U3396 ( .DIN1(n4476), .DIN2(n4477), .Q(n4166) );
  xor2s3 U3397 ( .DIN1(n6072), .DIN2(n4478), .Q(n4477) );
  xor2s3 U3398 ( .DIN1(n6070), .DIN2(n6071), .Q(n4478) );
  xor2s3 U3399 ( .DIN1(n6073), .DIN2(n6694), .Q(n4476) );
  nnd2s3 U3400 ( .DIN1(n3348), .DIN2(n6669), .Q(n4474) );
  xor2s3 U3401 ( .DIN1(n4479), .DIN2(n4480), .Q(n3348) );
  xor2s3 U3402 ( .DIN1(n6076), .DIN2(n4481), .Q(n4480) );
  xor2s3 U3403 ( .DIN1(n6074), .DIN2(n6075), .Q(n4481) );
  xor2s3 U3404 ( .DIN1(n6077), .DIN2(n6695), .Q(n4479) );
  nnd2s3 U3405 ( .DIN1(n6596), .DIN2(n2236), .Q(n4473) );
  nnd2s3 U3406 ( .DIN1(n6565), .DIN2(n2181), .Q(n4472) );
  nnd4s2 U3407 ( .DIN1(n4482), .DIN2(n4483), .DIN3(n4484), .DIN4(n4485), .Q(
        WX1943) );
  nnd2s3 U3408 ( .DIN1(n4174), .DIN2(n6638), .Q(n4485) );
  xor2s3 U3409 ( .DIN1(n4486), .DIN2(n4487), .Q(n4174) );
  xor2s3 U3410 ( .DIN1(n6081), .DIN2(n4488), .Q(n4487) );
  xor2s3 U3411 ( .DIN1(n6079), .DIN2(n6080), .Q(n4488) );
  xor2s3 U3412 ( .DIN1(n6082), .DIN2(n6695), .Q(n4486) );
  nnd2s3 U3413 ( .DIN1(n3354), .DIN2(n6669), .Q(n4484) );
  xor2s3 U3414 ( .DIN1(n4489), .DIN2(n4490), .Q(n3354) );
  xor2s3 U3415 ( .DIN1(n6085), .DIN2(n4491), .Q(n4490) );
  xor2s3 U3416 ( .DIN1(n6083), .DIN2(n6084), .Q(n4491) );
  xor2s3 U3417 ( .DIN1(n6086), .DIN2(n6695), .Q(n4489) );
  nnd2s3 U3418 ( .DIN1(n6596), .DIN2(n2237), .Q(n4483) );
  nnd2s3 U3419 ( .DIN1(n6565), .DIN2(n2180), .Q(n4482) );
  nnd4s2 U3420 ( .DIN1(n4492), .DIN2(n4493), .DIN3(n4494), .DIN4(n4495), .Q(
        WX1941) );
  nnd2s3 U3421 ( .DIN1(n4182), .DIN2(n6638), .Q(n4495) );
  xor2s3 U3422 ( .DIN1(n4496), .DIN2(n4497), .Q(n4182) );
  xor2s3 U3423 ( .DIN1(n6090), .DIN2(n4498), .Q(n4497) );
  xor2s3 U3424 ( .DIN1(n6088), .DIN2(n6089), .Q(n4498) );
  xor2s3 U3425 ( .DIN1(n6091), .DIN2(n6695), .Q(n4496) );
  nnd2s3 U3426 ( .DIN1(n3370), .DIN2(n6669), .Q(n4494) );
  xor2s3 U3427 ( .DIN1(n4499), .DIN2(n4500), .Q(n3370) );
  xor2s3 U3428 ( .DIN1(n6094), .DIN2(n4501), .Q(n4500) );
  xor2s3 U3429 ( .DIN1(n6092), .DIN2(n6093), .Q(n4501) );
  xor2s3 U3430 ( .DIN1(n6095), .DIN2(n6695), .Q(n4499) );
  nnd2s3 U3431 ( .DIN1(n6596), .DIN2(n2238), .Q(n4493) );
  nnd2s3 U3432 ( .DIN1(n6565), .DIN2(n2179), .Q(n4492) );
  nnd4s2 U3433 ( .DIN1(n4502), .DIN2(n4503), .DIN3(n4504), .DIN4(n4505), .Q(
        WX1939) );
  nnd2s3 U3434 ( .DIN1(n4190), .DIN2(n6638), .Q(n4505) );
  xor2s3 U3435 ( .DIN1(n4506), .DIN2(n4507), .Q(n4190) );
  xor2s3 U3436 ( .DIN1(n6099), .DIN2(n4508), .Q(n4507) );
  xor2s3 U3437 ( .DIN1(n6097), .DIN2(n6098), .Q(n4508) );
  xor2s3 U3438 ( .DIN1(n6100), .DIN2(n6695), .Q(n4506) );
  nnd2s3 U3439 ( .DIN1(n3387), .DIN2(n6669), .Q(n4504) );
  xor2s3 U3440 ( .DIN1(n4509), .DIN2(n4510), .Q(n3387) );
  xor2s3 U3441 ( .DIN1(n6103), .DIN2(n4511), .Q(n4510) );
  xor2s3 U3442 ( .DIN1(n6101), .DIN2(n6102), .Q(n4511) );
  xor2s3 U3443 ( .DIN1(n6104), .DIN2(n6695), .Q(n4509) );
  nnd2s3 U3444 ( .DIN1(n6596), .DIN2(n2239), .Q(n4503) );
  nnd2s3 U3445 ( .DIN1(n6565), .DIN2(n2178), .Q(n4502) );
  nnd4s2 U3446 ( .DIN1(n4512), .DIN2(n4513), .DIN3(n4514), .DIN4(n4515), .Q(
        WX1937) );
  nnd2s3 U3447 ( .DIN1(n4198), .DIN2(n6638), .Q(n4515) );
  xor2s3 U3448 ( .DIN1(n4516), .DIN2(n4517), .Q(n4198) );
  xor2s3 U3449 ( .DIN1(n6108), .DIN2(n4518), .Q(n4517) );
  xor2s3 U3450 ( .DIN1(n6106), .DIN2(n6107), .Q(n4518) );
  xor2s3 U3451 ( .DIN1(n6109), .DIN2(n6695), .Q(n4516) );
  nnd2s3 U3452 ( .DIN1(n3405), .DIN2(n6669), .Q(n4514) );
  xor2s3 U3453 ( .DIN1(n4519), .DIN2(n4520), .Q(n3405) );
  xor2s3 U3454 ( .DIN1(n6112), .DIN2(n4521), .Q(n4520) );
  xor2s3 U3455 ( .DIN1(n6110), .DIN2(n6111), .Q(n4521) );
  xor2s3 U3456 ( .DIN1(n6113), .DIN2(n6695), .Q(n4519) );
  nnd2s3 U3457 ( .DIN1(n6596), .DIN2(n2240), .Q(n4513) );
  nnd2s3 U3458 ( .DIN1(n6565), .DIN2(n2177), .Q(n4512) );
  nor2s3 U3459 ( .DIN1(n6803), .DIN2(n2240), .Q(WX1839) );
  nor2s3 U3460 ( .DIN1(n6116), .DIN2(n6757), .Q(WX1837) );
  nor2s3 U3461 ( .DIN1(n6117), .DIN2(n6757), .Q(WX1835) );
  nor2s3 U3462 ( .DIN1(n6118), .DIN2(n6757), .Q(WX1833) );
  nor2s3 U3463 ( .DIN1(n6119), .DIN2(n6757), .Q(WX1831) );
  nor2s3 U3464 ( .DIN1(n6120), .DIN2(n6757), .Q(WX1829) );
  nor2s3 U3465 ( .DIN1(n6121), .DIN2(n6757), .Q(WX1827) );
  nor2s3 U3466 ( .DIN1(n6122), .DIN2(n6757), .Q(WX1825) );
  nor2s3 U3467 ( .DIN1(n6123), .DIN2(n6756), .Q(WX1823) );
  nor2s3 U3468 ( .DIN1(n6124), .DIN2(n6756), .Q(WX1821) );
  nor2s3 U3469 ( .DIN1(n6125), .DIN2(n6756), .Q(WX1819) );
  nor2s3 U3470 ( .DIN1(n6126), .DIN2(n6756), .Q(WX1817) );
  nor2s3 U3471 ( .DIN1(n6127), .DIN2(n6756), .Q(WX1815) );
  nor2s3 U3472 ( .DIN1(n6128), .DIN2(n6756), .Q(WX1813) );
  nor2s3 U3473 ( .DIN1(n6129), .DIN2(n6756), .Q(WX1811) );
  nor2s3 U3474 ( .DIN1(n6130), .DIN2(n6756), .Q(WX1809) );
  nor2s3 U3475 ( .DIN1(n6131), .DIN2(n6761), .Q(WX1807) );
  nor2s3 U3476 ( .DIN1(n6132), .DIN2(n6775), .Q(WX1805) );
  nor2s3 U3477 ( .DIN1(n6133), .DIN2(n6775), .Q(WX1803) );
  nor2s3 U3478 ( .DIN1(n6134), .DIN2(n6775), .Q(WX1801) );
  nor2s3 U3479 ( .DIN1(n6135), .DIN2(n6775), .Q(WX1799) );
  nor2s3 U3480 ( .DIN1(n6136), .DIN2(n6775), .Q(WX1797) );
  nor2s3 U3481 ( .DIN1(n6137), .DIN2(n6775), .Q(WX1795) );
  nor2s3 U3482 ( .DIN1(n6138), .DIN2(n6775), .Q(WX1793) );
  nor2s3 U3483 ( .DIN1(n6139), .DIN2(n6775), .Q(WX1791) );
  nor2s3 U3484 ( .DIN1(n6140), .DIN2(n6775), .Q(WX1789) );
  nor2s3 U3485 ( .DIN1(n6141), .DIN2(n6775), .Q(WX1787) );
  nor2s3 U3486 ( .DIN1(n6142), .DIN2(n6775), .Q(WX1785) );
  nor2s3 U3487 ( .DIN1(n6143), .DIN2(n6775), .Q(WX1783) );
  nor2s3 U3488 ( .DIN1(n6144), .DIN2(n6774), .Q(WX1781) );
  nor2s3 U3489 ( .DIN1(n6145), .DIN2(n6774), .Q(WX1779) );
  nor2s3 U3490 ( .DIN1(n6146), .DIN2(n6774), .Q(WX1777) );
  nor2s3 U3491 ( .DIN1(n6805), .DIN2(n4522), .Q(WX1326) );
  xor2s3 U3492 ( .DIN1(n6147), .DIN2(n6534), .Q(n4522) );
  nor2s3 U3493 ( .DIN1(n6805), .DIN2(n4523), .Q(WX1324) );
  xor2s3 U3494 ( .DIN1(n6148), .DIN2(n6474), .Q(n4523) );
  nor2s3 U3495 ( .DIN1(n6805), .DIN2(n4524), .Q(WX1322) );
  xor2s3 U3496 ( .DIN1(n6149), .DIN2(n6482), .Q(n4524) );
  nor2s3 U3497 ( .DIN1(n6805), .DIN2(n4525), .Q(WX1320) );
  xor2s3 U3498 ( .DIN1(n6150), .DIN2(n6483), .Q(n4525) );
  nor2s3 U3499 ( .DIN1(n6805), .DIN2(n4526), .Q(WX1318) );
  xor2s3 U3500 ( .DIN1(n6151), .DIN2(n6486), .Q(n4526) );
  nor2s3 U3501 ( .DIN1(n6805), .DIN2(n4527), .Q(WX1316) );
  xor2s3 U3502 ( .DIN1(n6152), .DIN2(n6492), .Q(n4527) );
  nor2s3 U3503 ( .DIN1(n6805), .DIN2(n4528), .Q(WX1314) );
  xor2s3 U3504 ( .DIN1(n6153), .DIN2(n6500), .Q(n4528) );
  nor2s3 U3505 ( .DIN1(n6805), .DIN2(n4529), .Q(WX1312) );
  xor2s3 U3506 ( .DIN1(n6154), .DIN2(n6501), .Q(n4529) );
  nor2s3 U3507 ( .DIN1(n6805), .DIN2(n4530), .Q(WX1310) );
  xor2s3 U3508 ( .DIN1(n6155), .DIN2(n6511), .Q(n4530) );
  nor2s3 U3509 ( .DIN1(n6805), .DIN2(n4531), .Q(WX1308) );
  xor2s3 U3510 ( .DIN1(n6156), .DIN2(n6516), .Q(n4531) );
  nor2s3 U3511 ( .DIN1(n6805), .DIN2(n4532), .Q(WX1306) );
  xor2s3 U3512 ( .DIN1(n6157), .DIN2(n6517), .Q(n4532) );
  nor2s3 U3513 ( .DIN1(n6806), .DIN2(n4533), .Q(WX1304) );
  xor2s3 U3514 ( .DIN1(n6158), .DIN2(n6522), .Q(n4533) );
  nor2s3 U3515 ( .DIN1(n6806), .DIN2(n4534), .Q(WX1302) );
  xor2s3 U3516 ( .DIN1(n6159), .DIN2(n6477), .Q(n4534) );
  nor2s3 U3517 ( .DIN1(n6806), .DIN2(n4535), .Q(WX1300) );
  xor2s3 U3518 ( .DIN1(n6160), .DIN2(n6491), .Q(n4535) );
  nor2s3 U3519 ( .DIN1(n6806), .DIN2(n4536), .Q(WX1298) );
  xor2s3 U3520 ( .DIN1(n6161), .DIN2(n6495), .Q(n4536) );
  nor2s3 U3521 ( .DIN1(n4537), .DIN2(n6774), .Q(WX1296) );
  xnr2s3 U3522 ( .DIN1(n6510), .DIN2(n4538), .Q(n4537) );
  xor2s3 U3523 ( .DIN1(n6162), .DIN2(n6178), .Q(n4538) );
  nor2s3 U3524 ( .DIN1(n6806), .DIN2(n4539), .Q(WX1294) );
  xor2s3 U3525 ( .DIN1(n6163), .DIN2(n6438), .Q(n4539) );
  nor2s3 U3526 ( .DIN1(n6806), .DIN2(n4540), .Q(WX1292) );
  xor2s3 U3527 ( .DIN1(n6164), .DIN2(n6525), .Q(n4540) );
  nor2s3 U3528 ( .DIN1(n6806), .DIN2(n4541), .Q(WX1290) );
  xor2s3 U3529 ( .DIN1(n6165), .DIN2(n6447), .Q(n4541) );
  nor2s3 U3530 ( .DIN1(n6806), .DIN2(n4542), .Q(WX1288) );
  xor2s3 U3531 ( .DIN1(n6166), .DIN2(n6456), .Q(n4542) );
  nor2s3 U3532 ( .DIN1(n4543), .DIN2(n6774), .Q(WX1286) );
  xnr2s3 U3533 ( .DIN1(n6444), .DIN2(n4544), .Q(n4543) );
  xor2s3 U3534 ( .DIN1(n6167), .DIN2(n6178), .Q(n4544) );
  nor2s3 U3535 ( .DIN1(n6806), .DIN2(n4545), .Q(WX1284) );
  xor2s3 U3536 ( .DIN1(n6168), .DIN2(n6450), .Q(n4545) );
  nor2s3 U3537 ( .DIN1(n6806), .DIN2(n4546), .Q(WX1282) );
  xor2s3 U3538 ( .DIN1(n6169), .DIN2(n6506), .Q(n4546) );
  nor2s3 U3539 ( .DIN1(n6806), .DIN2(n4547), .Q(WX1280) );
  xor2s3 U3540 ( .DIN1(n6170), .DIN2(n6453), .Q(n4547) );
  nor2s3 U3541 ( .DIN1(n6806), .DIN2(n4548), .Q(WX1278) );
  xor2s3 U3542 ( .DIN1(n6171), .DIN2(n6465), .Q(n4548) );
  nor2s3 U3543 ( .DIN1(n6806), .DIN2(n4549), .Q(WX1276) );
  xor2s3 U3544 ( .DIN1(n6172), .DIN2(n6441), .Q(n4549) );
  nor2s3 U3545 ( .DIN1(n6807), .DIN2(n4550), .Q(WX1274) );
  xor2s3 U3546 ( .DIN1(n6173), .DIN2(n6459), .Q(n4550) );
  nor2s3 U3547 ( .DIN1(n4551), .DIN2(n6774), .Q(WX1272) );
  xnr2s3 U3548 ( .DIN1(n6471), .DIN2(n4552), .Q(n4551) );
  xor2s3 U3549 ( .DIN1(n6174), .DIN2(n6178), .Q(n4552) );
  nor2s3 U3550 ( .DIN1(n6807), .DIN2(n4553), .Q(WX1270) );
  xor2s3 U3551 ( .DIN1(n6175), .DIN2(n6468), .Q(n4553) );
  nor2s3 U3552 ( .DIN1(n6807), .DIN2(n4554), .Q(WX1268) );
  xor2s3 U3553 ( .DIN1(n6176), .DIN2(n6437), .Q(n4554) );
  nor2s3 U3554 ( .DIN1(n6807), .DIN2(n4555), .Q(WX1266) );
  xor2s3 U3555 ( .DIN1(n6177), .DIN2(n6530), .Q(n4555) );
  nor2s3 U3556 ( .DIN1(n6807), .DIN2(n4556), .Q(WX1264) );
  xor2s3 U3557 ( .DIN1(n6178), .DIN2(n6462), .Q(n4556) );
  nor2s3 U3558 ( .DIN1(n6807), .DIN2(n4557), .Q(WX11670) );
  xor2s3 U3559 ( .DIN1(n6336), .DIN2(n6341), .Q(n4557) );
  nor2s3 U3560 ( .DIN1(n6807), .DIN2(n4558), .Q(WX11668) );
  xor2s3 U3561 ( .DIN1(n6331), .DIN2(n6335), .Q(n4558) );
  nor2s3 U3562 ( .DIN1(n6807), .DIN2(n4559), .Q(WX11666) );
  xor2s3 U3563 ( .DIN1(n6326), .DIN2(n6330), .Q(n4559) );
  nor2s3 U3564 ( .DIN1(n6807), .DIN2(n4560), .Q(WX11664) );
  xor2s3 U3565 ( .DIN1(n6321), .DIN2(n6325), .Q(n4560) );
  nor2s3 U3566 ( .DIN1(n6807), .DIN2(n4561), .Q(WX11662) );
  xor2s3 U3567 ( .DIN1(n6316), .DIN2(n6320), .Q(n4561) );
  nor2s3 U3568 ( .DIN1(n6807), .DIN2(n4562), .Q(WX11660) );
  xor2s3 U3569 ( .DIN1(n6311), .DIN2(n6315), .Q(n4562) );
  nor2s3 U3570 ( .DIN1(n6807), .DIN2(n4563), .Q(WX11658) );
  xor2s3 U3571 ( .DIN1(n6306), .DIN2(n6310), .Q(n4563) );
  nor2s3 U3572 ( .DIN1(n6807), .DIN2(n4564), .Q(WX11656) );
  xor2s3 U3573 ( .DIN1(n6301), .DIN2(n6305), .Q(n4564) );
  nor2s3 U3574 ( .DIN1(n6808), .DIN2(n4565), .Q(WX11654) );
  xor2s3 U3575 ( .DIN1(n6296), .DIN2(n6300), .Q(n4565) );
  nor2s3 U3576 ( .DIN1(n6808), .DIN2(n4566), .Q(WX11652) );
  xor2s3 U3577 ( .DIN1(n6291), .DIN2(n6295), .Q(n4566) );
  nor2s3 U3578 ( .DIN1(n6808), .DIN2(n4567), .Q(WX11650) );
  xor2s3 U3579 ( .DIN1(n6285), .DIN2(n6290), .Q(n4567) );
  nor2s3 U3580 ( .DIN1(n6808), .DIN2(n4568), .Q(WX11648) );
  xor2s3 U3581 ( .DIN1(n6280), .DIN2(n6284), .Q(n4568) );
  nor2s3 U3582 ( .DIN1(n6808), .DIN2(n4569), .Q(WX11646) );
  xor2s3 U3583 ( .DIN1(n6275), .DIN2(n6279), .Q(n4569) );
  nor2s3 U3584 ( .DIN1(n6808), .DIN2(n4570), .Q(WX11644) );
  xor2s3 U3585 ( .DIN1(n6270), .DIN2(n6274), .Q(n4570) );
  nor2s3 U3586 ( .DIN1(n6808), .DIN2(n4571), .Q(WX11642) );
  xor2s3 U3587 ( .DIN1(n6265), .DIN2(n6269), .Q(n4571) );
  nor2s3 U3588 ( .DIN1(n4572), .DIN2(n6774), .Q(WX11640) );
  xor2s3 U3589 ( .DIN1(n1729), .DIN2(n4573), .Q(n4572) );
  xor2s3 U3590 ( .DIN1(n6260), .DIN2(n6264), .Q(n4573) );
  nor2s3 U3591 ( .DIN1(n6808), .DIN2(n4574), .Q(WX11638) );
  xor2s3 U3592 ( .DIN1(n6256), .DIN2(n3332), .Q(n4574) );
  nor2s3 U3593 ( .DIN1(n6808), .DIN2(n4575), .Q(WX11636) );
  xor2s3 U3594 ( .DIN1(n6252), .DIN2(n3331), .Q(n4575) );
  nor2s3 U3595 ( .DIN1(n6808), .DIN2(n4576), .Q(WX11634) );
  xor2s3 U3596 ( .DIN1(n6248), .DIN2(n3330), .Q(n4576) );
  nor2s3 U3597 ( .DIN1(n6808), .DIN2(n4577), .Q(WX11632) );
  xor2s3 U3598 ( .DIN1(n6244), .DIN2(n3329), .Q(n4577) );
  nor2s3 U3599 ( .DIN1(n4578), .DIN2(n6774), .Q(WX11630) );
  xnr2s3 U3600 ( .DIN1(n3328), .DIN2(n4579), .Q(n4578) );
  xor2s3 U3601 ( .DIN1(n6240), .DIN2(n6337), .Q(n4579) );
  nor2s3 U3602 ( .DIN1(n6808), .DIN2(n4580), .Q(WX11628) );
  xor2s3 U3603 ( .DIN1(n6236), .DIN2(n3327), .Q(n4580) );
  nor2s3 U3604 ( .DIN1(n6788), .DIN2(n4581), .Q(WX11626) );
  xor2s3 U3605 ( .DIN1(n6232), .DIN2(n3326), .Q(n4581) );
  nor2s3 U3606 ( .DIN1(n6788), .DIN2(n4582), .Q(WX11624) );
  xor2s3 U3607 ( .DIN1(n6228), .DIN2(n3325), .Q(n4582) );
  nor2s3 U3608 ( .DIN1(n6789), .DIN2(n4583), .Q(WX11622) );
  xor2s3 U3609 ( .DIN1(n6224), .DIN2(n3324), .Q(n4583) );
  nor2s3 U3610 ( .DIN1(n6788), .DIN2(n4584), .Q(WX11620) );
  xor2s3 U3611 ( .DIN1(n6220), .DIN2(n3323), .Q(n4584) );
  nor2s3 U3612 ( .DIN1(n6789), .DIN2(n4585), .Q(WX11618) );
  xor2s3 U3613 ( .DIN1(n6216), .DIN2(n3322), .Q(n4585) );
  nor2s3 U3614 ( .DIN1(n4586), .DIN2(n6776), .Q(WX11616) );
  xnr2s3 U3615 ( .DIN1(n3321), .DIN2(n4587), .Q(n4586) );
  xor2s3 U3616 ( .DIN1(n6212), .DIN2(n6337), .Q(n4587) );
  nor2s3 U3617 ( .DIN1(n6789), .DIN2(n4588), .Q(WX11614) );
  xor2s3 U3618 ( .DIN1(n6208), .DIN2(n3320), .Q(n4588) );
  nor2s3 U3619 ( .DIN1(n6788), .DIN2(n4589), .Q(WX11612) );
  xor2s3 U3620 ( .DIN1(n6204), .DIN2(n3319), .Q(n4589) );
  nor2s3 U3621 ( .DIN1(n6789), .DIN2(n4590), .Q(WX11610) );
  xor2s3 U3622 ( .DIN1(n6200), .DIN2(n3318), .Q(n4590) );
  nor2s3 U3623 ( .DIN1(n6788), .DIN2(n4591), .Q(WX11608) );
  xor2s3 U3624 ( .DIN1(n6337), .DIN2(n3317), .Q(n4591) );
  nor2s3 U3625 ( .DIN1(n6199), .DIN2(n6774), .Q(WX11242) );
  nor2s3 U3626 ( .DIN1(n6203), .DIN2(n6774), .Q(WX11240) );
  nor2s3 U3627 ( .DIN1(n6207), .DIN2(n6774), .Q(WX11238) );
  nor2s3 U3628 ( .DIN1(n6211), .DIN2(n6774), .Q(WX11236) );
  nor2s3 U3629 ( .DIN1(n6215), .DIN2(n6773), .Q(WX11234) );
  nor2s3 U3630 ( .DIN1(n6219), .DIN2(n6773), .Q(WX11232) );
  nor2s3 U3631 ( .DIN1(n6223), .DIN2(n6773), .Q(WX11230) );
  nor2s3 U3632 ( .DIN1(n6227), .DIN2(n6773), .Q(WX11228) );
  nor2s3 U3633 ( .DIN1(n6231), .DIN2(n6773), .Q(WX11226) );
  nor2s3 U3634 ( .DIN1(n6235), .DIN2(n6773), .Q(WX11224) );
  nor2s3 U3635 ( .DIN1(n6239), .DIN2(n6773), .Q(WX11222) );
  nor2s3 U3636 ( .DIN1(n6243), .DIN2(n6773), .Q(WX11220) );
  nor2s3 U3637 ( .DIN1(n6247), .DIN2(n6773), .Q(WX11218) );
  nor2s3 U3638 ( .DIN1(n6251), .DIN2(n6773), .Q(WX11216) );
  nor2s3 U3639 ( .DIN1(n6255), .DIN2(n6773), .Q(WX11214) );
  nor2s3 U3640 ( .DIN1(n6259), .DIN2(n6773), .Q(WX11212) );
  nor2s3 U3641 ( .DIN1(n6263), .DIN2(n6772), .Q(WX11210) );
  nor2s3 U3642 ( .DIN1(n6268), .DIN2(n6772), .Q(WX11208) );
  nor2s3 U3643 ( .DIN1(n6273), .DIN2(n6772), .Q(WX11206) );
  nor2s3 U3644 ( .DIN1(n6278), .DIN2(n6772), .Q(WX11204) );
  nor2s3 U3645 ( .DIN1(n6283), .DIN2(n6772), .Q(WX11202) );
  nor2s3 U3646 ( .DIN1(n6289), .DIN2(n6772), .Q(WX11200) );
  nor2s3 U3647 ( .DIN1(n6294), .DIN2(n6772), .Q(WX11198) );
  nor2s3 U3648 ( .DIN1(n6299), .DIN2(n6772), .Q(WX11196) );
  nor2s3 U3649 ( .DIN1(n6304), .DIN2(n6772), .Q(WX11194) );
  nor2s3 U3650 ( .DIN1(n6309), .DIN2(n6772), .Q(WX11192) );
  nor2s3 U3651 ( .DIN1(n6314), .DIN2(n6772), .Q(WX11190) );
  nor2s3 U3652 ( .DIN1(n6319), .DIN2(n6772), .Q(WX11188) );
  nor2s3 U3653 ( .DIN1(n6324), .DIN2(n6771), .Q(WX11186) );
  nor2s3 U3654 ( .DIN1(n6329), .DIN2(n6771), .Q(WX11184) );
  nor2s3 U3655 ( .DIN1(n6334), .DIN2(n6771), .Q(WX11182) );
  nor2s3 U3656 ( .DIN1(n6340), .DIN2(n6771), .Q(WX11180) );
  and2s3 U3657 ( .DIN1(RESET), .DIN2(n6198), .Q(WX11178) );
  and2s3 U3658 ( .DIN1(RESET), .DIN2(n6202), .Q(WX11176) );
  and2s3 U3659 ( .DIN1(RESET), .DIN2(n6206), .Q(WX11174) );
  and2s3 U3660 ( .DIN1(RESET), .DIN2(n6210), .Q(WX11172) );
  and2s3 U3661 ( .DIN1(RESET), .DIN2(n6214), .Q(WX11170) );
  and2s3 U3662 ( .DIN1(RESET), .DIN2(n6218), .Q(WX11168) );
  and2s3 U3663 ( .DIN1(RESET), .DIN2(n6222), .Q(WX11166) );
  and2s3 U3664 ( .DIN1(RESET), .DIN2(n6226), .Q(WX11164) );
  and2s3 U3665 ( .DIN1(RESET), .DIN2(n6230), .Q(WX11162) );
  and2s3 U3666 ( .DIN1(RESET), .DIN2(n6234), .Q(WX11160) );
  and2s3 U3667 ( .DIN1(RESET), .DIN2(n6238), .Q(WX11158) );
  and2s3 U3668 ( .DIN1(RESET), .DIN2(n6242), .Q(WX11156) );
  and2s3 U3669 ( .DIN1(RESET), .DIN2(n6246), .Q(WX11154) );
  and2s3 U3670 ( .DIN1(RESET), .DIN2(n6250), .Q(WX11152) );
  and2s3 U3671 ( .DIN1(RESET), .DIN2(n6254), .Q(WX11150) );
  and2s3 U3672 ( .DIN1(RESET), .DIN2(n6258), .Q(WX11148) );
  and2s3 U3673 ( .DIN1(RESET), .DIN2(n6262), .Q(WX11146) );
  and2s3 U3674 ( .DIN1(RESET), .DIN2(n6267), .Q(WX11144) );
  and2s3 U3675 ( .DIN1(RESET), .DIN2(n6272), .Q(WX11142) );
  and2s3 U3676 ( .DIN1(RESET), .DIN2(n6277), .Q(WX11140) );
  and2s3 U3677 ( .DIN1(RESET), .DIN2(n6282), .Q(WX11138) );
  and2s3 U3678 ( .DIN1(RESET), .DIN2(n6288), .Q(WX11136) );
  and2s3 U3679 ( .DIN1(RESET), .DIN2(n6293), .Q(WX11134) );
  and2s3 U3680 ( .DIN1(RESET), .DIN2(n6298), .Q(WX11132) );
  and2s3 U3681 ( .DIN1(RESET), .DIN2(n6303), .Q(WX11130) );
  and2s3 U3682 ( .DIN1(RESET), .DIN2(n6308), .Q(WX11128) );
  and2s3 U3683 ( .DIN1(RESET), .DIN2(n6313), .Q(WX11126) );
  and2s3 U3684 ( .DIN1(RESET), .DIN2(n6318), .Q(WX11124) );
  and2s3 U3685 ( .DIN1(RESET), .DIN2(n6323), .Q(WX11122) );
  and2s3 U3686 ( .DIN1(RESET), .DIN2(n6328), .Q(WX11120) );
  and2s3 U3687 ( .DIN1(RESET), .DIN2(n6333), .Q(WX11118) );
  and2s3 U3688 ( .DIN1(RESET), .DIN2(n6339), .Q(WX11116) );
  nor2s3 U3689 ( .DIN1(n6197), .DIN2(n6771), .Q(WX11114) );
  nor2s3 U3690 ( .DIN1(n6201), .DIN2(n6771), .Q(WX11112) );
  nor2s3 U3691 ( .DIN1(n6205), .DIN2(n6771), .Q(WX11110) );
  nor2s3 U3692 ( .DIN1(n6209), .DIN2(n6771), .Q(WX11108) );
  nor2s3 U3693 ( .DIN1(n6213), .DIN2(n6771), .Q(WX11106) );
  nor2s3 U3694 ( .DIN1(n6217), .DIN2(n6771), .Q(WX11104) );
  nor2s3 U3695 ( .DIN1(n6221), .DIN2(n6771), .Q(WX11102) );
  nor2s3 U3696 ( .DIN1(n6225), .DIN2(n6770), .Q(WX11100) );
  nor2s3 U3697 ( .DIN1(n6229), .DIN2(n6770), .Q(WX11098) );
  nor2s3 U3698 ( .DIN1(n6233), .DIN2(n6770), .Q(WX11096) );
  nor2s3 U3699 ( .DIN1(n6237), .DIN2(n6770), .Q(WX11094) );
  nor2s3 U3700 ( .DIN1(n6241), .DIN2(n6770), .Q(WX11092) );
  nor2s3 U3701 ( .DIN1(n6245), .DIN2(n6770), .Q(WX11090) );
  nor2s3 U3702 ( .DIN1(n6249), .DIN2(n6770), .Q(WX11088) );
  nor2s3 U3703 ( .DIN1(n6253), .DIN2(n6770), .Q(WX11086) );
  nor2s3 U3704 ( .DIN1(n6257), .DIN2(n6770), .Q(WX11084) );
  nor2s3 U3705 ( .DIN1(n6261), .DIN2(n6770), .Q(WX11082) );
  nor2s3 U3706 ( .DIN1(n6266), .DIN2(n6770), .Q(WX11080) );
  nor2s3 U3707 ( .DIN1(n6271), .DIN2(n6770), .Q(WX11078) );
  nor2s3 U3708 ( .DIN1(n6276), .DIN2(n6769), .Q(WX11076) );
  nor2s3 U3709 ( .DIN1(n6281), .DIN2(n6769), .Q(WX11074) );
  nor2s3 U3710 ( .DIN1(n6287), .DIN2(n6769), .Q(WX11072) );
  nor2s3 U3711 ( .DIN1(n6292), .DIN2(n6769), .Q(WX11070) );
  nor2s3 U3712 ( .DIN1(n6297), .DIN2(n6769), .Q(WX11068) );
  nor2s3 U3713 ( .DIN1(n6302), .DIN2(n6769), .Q(WX11066) );
  nor2s3 U3714 ( .DIN1(n6307), .DIN2(n6769), .Q(WX11064) );
  nor2s3 U3715 ( .DIN1(n6312), .DIN2(n6769), .Q(WX11062) );
  nor2s3 U3716 ( .DIN1(n6317), .DIN2(n6769), .Q(WX11060) );
  nor2s3 U3717 ( .DIN1(n6322), .DIN2(n6769), .Q(WX11058) );
  nor2s3 U3718 ( .DIN1(n6327), .DIN2(n6769), .Q(WX11056) );
  nor2s3 U3719 ( .DIN1(n6332), .DIN2(n6769), .Q(WX11054) );
  nor2s3 U3720 ( .DIN1(n6338), .DIN2(n6768), .Q(WX11052) );
  nnd4s2 U3721 ( .DIN1(n4592), .DIN2(n4593), .DIN3(n4594), .DIN4(n4595), .Q(
        WX11050) );
  nnd2s3 U3722 ( .DIN1(n2315), .DIN2(n6669), .Q(n4595) );
  xor2s3 U3723 ( .DIN1(n4596), .DIN2(n4597), .Q(n2315) );
  xor2s3 U3724 ( .DIN1(n6197), .DIN2(n6198), .Q(n4597) );
  xnr2s3 U3725 ( .DIN1(n3317), .DIN2(n6199), .Q(n4596) );
  nnd2s3 U3726 ( .DIN1(n6596), .DIN2(n1761), .Q(n4594) );
  nnd2s3 U3727 ( .DIN1(DATA_0_0), .DIN2(n6638), .Q(n4593) );
  nnd2s3 U3728 ( .DIN1(n6565), .DIN2(n1760), .Q(n4592) );
  nnd4s2 U3729 ( .DIN1(n4598), .DIN2(n4599), .DIN3(n4600), .DIN4(n4601), .Q(
        WX11048) );
  nnd2s3 U3730 ( .DIN1(n2323), .DIN2(n6669), .Q(n4601) );
  xor2s3 U3731 ( .DIN1(n4602), .DIN2(n4603), .Q(n2323) );
  xor2s3 U3732 ( .DIN1(n6201), .DIN2(n6202), .Q(n4603) );
  xnr2s3 U3733 ( .DIN1(n3318), .DIN2(n6203), .Q(n4602) );
  nnd2s3 U3734 ( .DIN1(n6596), .DIN2(n1762), .Q(n4600) );
  nnd2s3 U3735 ( .DIN1(DATA_0_1), .DIN2(n6638), .Q(n4599) );
  nnd2s3 U3736 ( .DIN1(n6565), .DIN2(n1759), .Q(n4598) );
  nnd4s2 U3737 ( .DIN1(n4604), .DIN2(n4605), .DIN3(n4606), .DIN4(n4607), .Q(
        WX11046) );
  nnd2s3 U3738 ( .DIN1(n2329), .DIN2(n6669), .Q(n4607) );
  xor2s3 U3739 ( .DIN1(n4608), .DIN2(n4609), .Q(n2329) );
  xor2s3 U3740 ( .DIN1(n6205), .DIN2(n6206), .Q(n4609) );
  xnr2s3 U3741 ( .DIN1(n3319), .DIN2(n6207), .Q(n4608) );
  nnd2s3 U3742 ( .DIN1(n6596), .DIN2(n1763), .Q(n4606) );
  nnd2s3 U3743 ( .DIN1(DATA_0_2), .DIN2(n6638), .Q(n4605) );
  nnd2s3 U3744 ( .DIN1(n6565), .DIN2(n1758), .Q(n4604) );
  nnd4s2 U3745 ( .DIN1(n4610), .DIN2(n4611), .DIN3(n4612), .DIN4(n4613), .Q(
        WX11044) );
  nnd2s3 U3746 ( .DIN1(n2335), .DIN2(n6669), .Q(n4613) );
  xor2s3 U3747 ( .DIN1(n4614), .DIN2(n4615), .Q(n2335) );
  xor2s3 U3748 ( .DIN1(n6209), .DIN2(n6210), .Q(n4615) );
  xnr2s3 U3749 ( .DIN1(n3320), .DIN2(n6211), .Q(n4614) );
  nnd2s3 U3750 ( .DIN1(n6596), .DIN2(n1764), .Q(n4612) );
  nnd2s3 U3751 ( .DIN1(DATA_0_3), .DIN2(n6638), .Q(n4611) );
  nnd2s3 U3752 ( .DIN1(n6565), .DIN2(n1757), .Q(n4610) );
  nnd4s2 U3753 ( .DIN1(n4616), .DIN2(n4617), .DIN3(n4618), .DIN4(n4619), .Q(
        WX11042) );
  nnd2s3 U3754 ( .DIN1(n2341), .DIN2(n6669), .Q(n4619) );
  xor2s3 U3755 ( .DIN1(n4620), .DIN2(n4621), .Q(n2341) );
  xor2s3 U3756 ( .DIN1(n6213), .DIN2(n6214), .Q(n4621) );
  xnr2s3 U3757 ( .DIN1(n3321), .DIN2(n6215), .Q(n4620) );
  nnd2s3 U3758 ( .DIN1(n6596), .DIN2(n1765), .Q(n4618) );
  nnd2s3 U3759 ( .DIN1(DATA_0_4), .DIN2(n6638), .Q(n4617) );
  nnd2s3 U3760 ( .DIN1(n6565), .DIN2(n1756), .Q(n4616) );
  nnd4s2 U3761 ( .DIN1(n4622), .DIN2(n4623), .DIN3(n4624), .DIN4(n4625), .Q(
        WX11040) );
  nnd2s3 U3762 ( .DIN1(n2347), .DIN2(n6669), .Q(n4625) );
  xor2s3 U3763 ( .DIN1(n4626), .DIN2(n4627), .Q(n2347) );
  xor2s3 U3764 ( .DIN1(n6217), .DIN2(n6218), .Q(n4627) );
  xnr2s3 U3765 ( .DIN1(n3322), .DIN2(n6219), .Q(n4626) );
  nnd2s3 U3766 ( .DIN1(n6596), .DIN2(n1766), .Q(n4624) );
  nnd2s3 U3767 ( .DIN1(DATA_0_5), .DIN2(n6638), .Q(n4623) );
  nnd2s3 U3768 ( .DIN1(n6565), .DIN2(n1755), .Q(n4622) );
  nnd4s2 U3769 ( .DIN1(n4628), .DIN2(n4629), .DIN3(n4630), .DIN4(n4631), .Q(
        WX11038) );
  nnd2s3 U3770 ( .DIN1(n2353), .DIN2(n6668), .Q(n4631) );
  xor2s3 U3771 ( .DIN1(n4632), .DIN2(n4633), .Q(n2353) );
  xor2s3 U3772 ( .DIN1(n6221), .DIN2(n6222), .Q(n4633) );
  xnr2s3 U3773 ( .DIN1(n3323), .DIN2(n6223), .Q(n4632) );
  nnd2s3 U3774 ( .DIN1(n6595), .DIN2(n1767), .Q(n4630) );
  nnd2s3 U3775 ( .DIN1(DATA_0_6), .DIN2(n6637), .Q(n4629) );
  nnd2s3 U3776 ( .DIN1(n6564), .DIN2(n1754), .Q(n4628) );
  nnd4s2 U3777 ( .DIN1(n4634), .DIN2(n4635), .DIN3(n4636), .DIN4(n4637), .Q(
        WX11036) );
  nnd2s3 U3778 ( .DIN1(n2359), .DIN2(n6668), .Q(n4637) );
  xor2s3 U3779 ( .DIN1(n4638), .DIN2(n4639), .Q(n2359) );
  xor2s3 U3780 ( .DIN1(n6225), .DIN2(n6226), .Q(n4639) );
  xnr2s3 U3781 ( .DIN1(n3324), .DIN2(n6227), .Q(n4638) );
  nnd2s3 U3782 ( .DIN1(n6595), .DIN2(n1768), .Q(n4636) );
  nnd2s3 U3783 ( .DIN1(DATA_0_7), .DIN2(n6637), .Q(n4635) );
  nnd2s3 U3784 ( .DIN1(n6564), .DIN2(n1753), .Q(n4634) );
  nnd4s2 U3785 ( .DIN1(n4640), .DIN2(n4641), .DIN3(n4642), .DIN4(n4643), .Q(
        WX11034) );
  nnd2s3 U3786 ( .DIN1(n2365), .DIN2(n6668), .Q(n4643) );
  xor2s3 U3787 ( .DIN1(n4644), .DIN2(n4645), .Q(n2365) );
  xor2s3 U3788 ( .DIN1(n6229), .DIN2(n6230), .Q(n4645) );
  xnr2s3 U3789 ( .DIN1(n3325), .DIN2(n6231), .Q(n4644) );
  nnd2s3 U3790 ( .DIN1(n6595), .DIN2(n1769), .Q(n4642) );
  nnd2s3 U3791 ( .DIN1(DATA_0_8), .DIN2(n6637), .Q(n4641) );
  nnd2s3 U3792 ( .DIN1(n6564), .DIN2(n1752), .Q(n4640) );
  nnd4s2 U3793 ( .DIN1(n4646), .DIN2(n4647), .DIN3(n4648), .DIN4(n4649), .Q(
        WX11032) );
  nnd2s3 U3794 ( .DIN1(n2371), .DIN2(n6668), .Q(n4649) );
  xor2s3 U3795 ( .DIN1(n4650), .DIN2(n4651), .Q(n2371) );
  xor2s3 U3796 ( .DIN1(n6233), .DIN2(n6234), .Q(n4651) );
  xnr2s3 U3797 ( .DIN1(n3326), .DIN2(n6235), .Q(n4650) );
  nnd2s3 U3798 ( .DIN1(n6595), .DIN2(n1770), .Q(n4648) );
  nnd2s3 U3799 ( .DIN1(DATA_0_9), .DIN2(n6637), .Q(n4647) );
  nnd2s3 U3800 ( .DIN1(n6564), .DIN2(n1751), .Q(n4646) );
  nnd4s2 U3801 ( .DIN1(n4652), .DIN2(n4653), .DIN3(n4654), .DIN4(n4655), .Q(
        WX11030) );
  nnd2s3 U3802 ( .DIN1(n2377), .DIN2(n6668), .Q(n4655) );
  xor2s3 U3803 ( .DIN1(n4656), .DIN2(n4657), .Q(n2377) );
  xor2s3 U3804 ( .DIN1(n6237), .DIN2(n6238), .Q(n4657) );
  xnr2s3 U3805 ( .DIN1(n3327), .DIN2(n6239), .Q(n4656) );
  nnd2s3 U3806 ( .DIN1(n6595), .DIN2(n1771), .Q(n4654) );
  nnd2s3 U3807 ( .DIN1(DATA_0_10), .DIN2(n6637), .Q(n4653) );
  nnd2s3 U3808 ( .DIN1(n6564), .DIN2(n1750), .Q(n4652) );
  nnd4s2 U3809 ( .DIN1(n4658), .DIN2(n4659), .DIN3(n4660), .DIN4(n4661), .Q(
        WX11028) );
  nnd2s3 U3810 ( .DIN1(n2383), .DIN2(n6668), .Q(n4661) );
  xor2s3 U3811 ( .DIN1(n4662), .DIN2(n4663), .Q(n2383) );
  xor2s3 U3812 ( .DIN1(n6241), .DIN2(n6242), .Q(n4663) );
  xnr2s3 U3813 ( .DIN1(n3328), .DIN2(n6243), .Q(n4662) );
  nnd2s3 U3814 ( .DIN1(n6595), .DIN2(n1772), .Q(n4660) );
  nnd2s3 U3815 ( .DIN1(DATA_0_11), .DIN2(n6637), .Q(n4659) );
  nnd2s3 U3816 ( .DIN1(n6564), .DIN2(n1749), .Q(n4658) );
  nnd4s2 U3817 ( .DIN1(n4664), .DIN2(n4665), .DIN3(n4666), .DIN4(n4667), .Q(
        WX11026) );
  nnd2s3 U3818 ( .DIN1(n2389), .DIN2(n6668), .Q(n4667) );
  xor2s3 U3819 ( .DIN1(n4668), .DIN2(n4669), .Q(n2389) );
  xor2s3 U3820 ( .DIN1(n6245), .DIN2(n6246), .Q(n4669) );
  xnr2s3 U3821 ( .DIN1(n3329), .DIN2(n6247), .Q(n4668) );
  nnd2s3 U3822 ( .DIN1(n6595), .DIN2(n1773), .Q(n4666) );
  nnd2s3 U3823 ( .DIN1(DATA_0_12), .DIN2(n6637), .Q(n4665) );
  nnd2s3 U3824 ( .DIN1(n6564), .DIN2(n1748), .Q(n4664) );
  nnd4s2 U3825 ( .DIN1(n4670), .DIN2(n4671), .DIN3(n4672), .DIN4(n4673), .Q(
        WX11024) );
  nnd2s3 U3826 ( .DIN1(n2395), .DIN2(n6668), .Q(n4673) );
  xor2s3 U3827 ( .DIN1(n4674), .DIN2(n4675), .Q(n2395) );
  xor2s3 U3828 ( .DIN1(n6249), .DIN2(n6250), .Q(n4675) );
  xnr2s3 U3829 ( .DIN1(n3330), .DIN2(n6251), .Q(n4674) );
  nnd2s3 U3830 ( .DIN1(n6595), .DIN2(n1774), .Q(n4672) );
  nnd2s3 U3831 ( .DIN1(DATA_0_13), .DIN2(n6637), .Q(n4671) );
  nnd2s3 U3832 ( .DIN1(n6564), .DIN2(n1747), .Q(n4670) );
  nnd4s2 U3833 ( .DIN1(n4676), .DIN2(n4677), .DIN3(n4678), .DIN4(n4679), .Q(
        WX11022) );
  nnd2s3 U3834 ( .DIN1(n2401), .DIN2(n6668), .Q(n4679) );
  xor2s3 U3835 ( .DIN1(n4680), .DIN2(n4681), .Q(n2401) );
  xor2s3 U3836 ( .DIN1(n6253), .DIN2(n6254), .Q(n4681) );
  xnr2s3 U3837 ( .DIN1(n3331), .DIN2(n6255), .Q(n4680) );
  nnd2s3 U3838 ( .DIN1(n6595), .DIN2(n1775), .Q(n4678) );
  nnd2s3 U3839 ( .DIN1(DATA_0_14), .DIN2(n6637), .Q(n4677) );
  nnd2s3 U3840 ( .DIN1(n6564), .DIN2(n1746), .Q(n4676) );
  nnd4s2 U3841 ( .DIN1(n4682), .DIN2(n4683), .DIN3(n4684), .DIN4(n4685), .Q(
        WX11020) );
  nnd2s3 U3842 ( .DIN1(n2407), .DIN2(n6668), .Q(n4685) );
  xor2s3 U3843 ( .DIN1(n4686), .DIN2(n4687), .Q(n2407) );
  xor2s3 U3844 ( .DIN1(n6257), .DIN2(n6258), .Q(n4687) );
  xnr2s3 U3845 ( .DIN1(n3332), .DIN2(n6259), .Q(n4686) );
  nnd2s3 U3846 ( .DIN1(n6595), .DIN2(n1776), .Q(n4684) );
  nnd2s3 U3847 ( .DIN1(DATA_0_15), .DIN2(n6637), .Q(n4683) );
  nnd2s3 U3848 ( .DIN1(n6564), .DIN2(n1745), .Q(n4682) );
  nnd4s2 U3849 ( .DIN1(n4688), .DIN2(n4689), .DIN3(n4690), .DIN4(n4691), .Q(
        WX11018) );
  nnd2s3 U3850 ( .DIN1(n2413), .DIN2(n6668), .Q(n4691) );
  xor2s3 U3851 ( .DIN1(n4692), .DIN2(n4693), .Q(n2413) );
  xor2s3 U3852 ( .DIN1(n6263), .DIN2(n4694), .Q(n4693) );
  xor2s3 U3853 ( .DIN1(n6261), .DIN2(n6262), .Q(n4694) );
  xor2s3 U3854 ( .DIN1(n6264), .DIN2(n6695), .Q(n4692) );
  nnd2s3 U3855 ( .DIN1(n6595), .DIN2(n1777), .Q(n4690) );
  nnd2s3 U3856 ( .DIN1(DATA_0_16), .DIN2(n6637), .Q(n4689) );
  nnd2s3 U3857 ( .DIN1(n6564), .DIN2(n1744), .Q(n4688) );
  nnd4s2 U3858 ( .DIN1(n4695), .DIN2(n4696), .DIN3(n4697), .DIN4(n4698), .Q(
        WX11016) );
  nnd2s3 U3859 ( .DIN1(n2419), .DIN2(n6668), .Q(n4698) );
  xor2s3 U3860 ( .DIN1(n4699), .DIN2(n4700), .Q(n2419) );
  xor2s3 U3861 ( .DIN1(n6268), .DIN2(n4701), .Q(n4700) );
  xor2s3 U3862 ( .DIN1(n6266), .DIN2(n6267), .Q(n4701) );
  xor2s3 U3863 ( .DIN1(n6269), .DIN2(n6695), .Q(n4699) );
  nnd2s3 U3864 ( .DIN1(n6595), .DIN2(n1778), .Q(n4697) );
  nnd2s3 U3865 ( .DIN1(DATA_0_17), .DIN2(n6637), .Q(n4696) );
  nnd2s3 U3866 ( .DIN1(n6564), .DIN2(n1743), .Q(n4695) );
  nnd4s2 U3867 ( .DIN1(n4702), .DIN2(n4703), .DIN3(n4704), .DIN4(n4705), .Q(
        WX11014) );
  nnd2s3 U3868 ( .DIN1(n2425), .DIN2(n6668), .Q(n4705) );
  xor2s3 U3869 ( .DIN1(n4706), .DIN2(n4707), .Q(n2425) );
  xor2s3 U3870 ( .DIN1(n6273), .DIN2(n4708), .Q(n4707) );
  xor2s3 U3871 ( .DIN1(n6271), .DIN2(n6272), .Q(n4708) );
  xor2s3 U3872 ( .DIN1(n6274), .DIN2(n6695), .Q(n4706) );
  nnd2s3 U3873 ( .DIN1(n6595), .DIN2(n1779), .Q(n4704) );
  nnd2s3 U3874 ( .DIN1(DATA_0_18), .DIN2(n6637), .Q(n4703) );
  nnd2s3 U3875 ( .DIN1(n6564), .DIN2(n1742), .Q(n4702) );
  nnd4s2 U3876 ( .DIN1(n4709), .DIN2(n4710), .DIN3(n4711), .DIN4(n4712), .Q(
        WX11012) );
  nnd2s3 U3877 ( .DIN1(n2431), .DIN2(n6667), .Q(n4712) );
  xor2s3 U3878 ( .DIN1(n4713), .DIN2(n4714), .Q(n2431) );
  xor2s3 U3879 ( .DIN1(n6278), .DIN2(n4715), .Q(n4714) );
  xor2s3 U3880 ( .DIN1(n6276), .DIN2(n6277), .Q(n4715) );
  xor2s3 U3881 ( .DIN1(n6279), .DIN2(n6695), .Q(n4713) );
  nnd2s3 U3882 ( .DIN1(n6594), .DIN2(n1780), .Q(n4711) );
  nnd2s3 U3883 ( .DIN1(DATA_0_19), .DIN2(n6636), .Q(n4710) );
  nnd2s3 U3884 ( .DIN1(n6563), .DIN2(n1741), .Q(n4709) );
  nnd4s2 U3885 ( .DIN1(n4716), .DIN2(n4717), .DIN3(n4718), .DIN4(n4719), .Q(
        WX11010) );
  nnd2s3 U3886 ( .DIN1(n2437), .DIN2(n6667), .Q(n4719) );
  xor2s3 U3887 ( .DIN1(n4720), .DIN2(n4721), .Q(n2437) );
  xor2s3 U3888 ( .DIN1(n6283), .DIN2(n4722), .Q(n4721) );
  xor2s3 U3889 ( .DIN1(n6281), .DIN2(n6282), .Q(n4722) );
  xor2s3 U3890 ( .DIN1(n6284), .DIN2(n6696), .Q(n4720) );
  nnd2s3 U3891 ( .DIN1(n6594), .DIN2(n1781), .Q(n4718) );
  nnd2s3 U3892 ( .DIN1(DATA_0_20), .DIN2(n6636), .Q(n4717) );
  nnd2s3 U3893 ( .DIN1(n6563), .DIN2(n1740), .Q(n4716) );
  nnd4s2 U3894 ( .DIN1(n4723), .DIN2(n4724), .DIN3(n4725), .DIN4(n4726), .Q(
        WX11008) );
  nnd2s3 U3895 ( .DIN1(n2443), .DIN2(n6667), .Q(n4726) );
  xor2s3 U3896 ( .DIN1(n4727), .DIN2(n4728), .Q(n2443) );
  xor2s3 U3897 ( .DIN1(n6289), .DIN2(n4729), .Q(n4728) );
  xor2s3 U3898 ( .DIN1(n6287), .DIN2(n6288), .Q(n4729) );
  xor2s3 U3899 ( .DIN1(n6290), .DIN2(n6696), .Q(n4727) );
  nnd2s3 U3900 ( .DIN1(n6594), .DIN2(n1782), .Q(n4725) );
  nnd2s3 U3901 ( .DIN1(DATA_0_21), .DIN2(n6636), .Q(n4724) );
  nnd2s3 U3902 ( .DIN1(n6563), .DIN2(n1739), .Q(n4723) );
  nnd4s2 U3903 ( .DIN1(n4730), .DIN2(n4731), .DIN3(n4732), .DIN4(n4733), .Q(
        WX11006) );
  nnd2s3 U3904 ( .DIN1(n2449), .DIN2(n6667), .Q(n4733) );
  xor2s3 U3905 ( .DIN1(n4734), .DIN2(n4735), .Q(n2449) );
  xor2s3 U3906 ( .DIN1(n6294), .DIN2(n4736), .Q(n4735) );
  xor2s3 U3907 ( .DIN1(n6292), .DIN2(n6293), .Q(n4736) );
  xor2s3 U3908 ( .DIN1(n6295), .DIN2(n6696), .Q(n4734) );
  nnd2s3 U3909 ( .DIN1(n6594), .DIN2(n1783), .Q(n4732) );
  nnd2s3 U3910 ( .DIN1(DATA_0_22), .DIN2(n6636), .Q(n4731) );
  nnd2s3 U3911 ( .DIN1(n6563), .DIN2(n1738), .Q(n4730) );
  nnd4s2 U3912 ( .DIN1(n4737), .DIN2(n4738), .DIN3(n4739), .DIN4(n4740), .Q(
        WX11004) );
  nnd2s3 U3913 ( .DIN1(n2455), .DIN2(n6667), .Q(n4740) );
  xor2s3 U3914 ( .DIN1(n4741), .DIN2(n4742), .Q(n2455) );
  xor2s3 U3915 ( .DIN1(n6299), .DIN2(n4743), .Q(n4742) );
  xor2s3 U3916 ( .DIN1(n6297), .DIN2(n6298), .Q(n4743) );
  xor2s3 U3917 ( .DIN1(n6300), .DIN2(n6696), .Q(n4741) );
  nnd2s3 U3918 ( .DIN1(n6594), .DIN2(n1784), .Q(n4739) );
  nnd2s3 U3919 ( .DIN1(DATA_0_23), .DIN2(n6636), .Q(n4738) );
  nnd2s3 U3920 ( .DIN1(n6563), .DIN2(n1737), .Q(n4737) );
  nnd4s2 U3921 ( .DIN1(n4744), .DIN2(n4745), .DIN3(n4746), .DIN4(n4747), .Q(
        WX11002) );
  nnd2s3 U3922 ( .DIN1(n2461), .DIN2(n6667), .Q(n4747) );
  xor2s3 U3923 ( .DIN1(n4748), .DIN2(n4749), .Q(n2461) );
  xor2s3 U3924 ( .DIN1(n6304), .DIN2(n4750), .Q(n4749) );
  xor2s3 U3925 ( .DIN1(n6302), .DIN2(n6303), .Q(n4750) );
  xor2s3 U3926 ( .DIN1(n6305), .DIN2(n6696), .Q(n4748) );
  nnd2s3 U3927 ( .DIN1(n6594), .DIN2(n1785), .Q(n4746) );
  nnd2s3 U3928 ( .DIN1(DATA_0_24), .DIN2(n6636), .Q(n4745) );
  nnd2s3 U3929 ( .DIN1(n6563), .DIN2(n1736), .Q(n4744) );
  nnd4s2 U3930 ( .DIN1(n4751), .DIN2(n4752), .DIN3(n4753), .DIN4(n4754), .Q(
        WX11000) );
  nnd2s3 U3931 ( .DIN1(n2467), .DIN2(n6667), .Q(n4754) );
  xor2s3 U3932 ( .DIN1(n4755), .DIN2(n4756), .Q(n2467) );
  xor2s3 U3933 ( .DIN1(n6309), .DIN2(n4757), .Q(n4756) );
  xor2s3 U3934 ( .DIN1(n6307), .DIN2(n6308), .Q(n4757) );
  xor2s3 U3935 ( .DIN1(n6310), .DIN2(n6696), .Q(n4755) );
  nnd2s3 U3936 ( .DIN1(n6594), .DIN2(n1786), .Q(n4753) );
  nnd2s3 U3937 ( .DIN1(DATA_0_25), .DIN2(n6636), .Q(n4752) );
  nnd2s3 U3938 ( .DIN1(n6563), .DIN2(n1735), .Q(n4751) );
  nnd4s2 U3939 ( .DIN1(n4758), .DIN2(n4759), .DIN3(n4760), .DIN4(n4761), .Q(
        WX10998) );
  nnd2s3 U3940 ( .DIN1(n2473), .DIN2(n6667), .Q(n4761) );
  xor2s3 U3941 ( .DIN1(n4762), .DIN2(n4763), .Q(n2473) );
  xor2s3 U3942 ( .DIN1(n6314), .DIN2(n4764), .Q(n4763) );
  xor2s3 U3943 ( .DIN1(n6312), .DIN2(n6313), .Q(n4764) );
  xor2s3 U3944 ( .DIN1(n6315), .DIN2(n6696), .Q(n4762) );
  nnd2s3 U3945 ( .DIN1(n6594), .DIN2(n1787), .Q(n4760) );
  nnd2s3 U3946 ( .DIN1(DATA_0_26), .DIN2(n6636), .Q(n4759) );
  nnd2s3 U3947 ( .DIN1(n6563), .DIN2(n1734), .Q(n4758) );
  nnd4s2 U3948 ( .DIN1(n4765), .DIN2(n4766), .DIN3(n4767), .DIN4(n4768), .Q(
        WX10996) );
  nnd2s3 U3949 ( .DIN1(n2479), .DIN2(n6667), .Q(n4768) );
  xor2s3 U3950 ( .DIN1(n4769), .DIN2(n4770), .Q(n2479) );
  xor2s3 U3951 ( .DIN1(n6319), .DIN2(n4771), .Q(n4770) );
  xor2s3 U3952 ( .DIN1(n6317), .DIN2(n6318), .Q(n4771) );
  xor2s3 U3953 ( .DIN1(n6320), .DIN2(n6696), .Q(n4769) );
  nnd2s3 U3954 ( .DIN1(n6594), .DIN2(n1788), .Q(n4767) );
  nnd2s3 U3955 ( .DIN1(DATA_0_27), .DIN2(n6636), .Q(n4766) );
  nnd2s3 U3956 ( .DIN1(n6563), .DIN2(n1733), .Q(n4765) );
  nnd4s2 U3957 ( .DIN1(n4772), .DIN2(n4773), .DIN3(n4774), .DIN4(n4775), .Q(
        WX10994) );
  nnd2s3 U3958 ( .DIN1(n2485), .DIN2(n6667), .Q(n4775) );
  xor2s3 U3959 ( .DIN1(n4776), .DIN2(n4777), .Q(n2485) );
  xor2s3 U3960 ( .DIN1(n6324), .DIN2(n4778), .Q(n4777) );
  xor2s3 U3961 ( .DIN1(n6322), .DIN2(n6323), .Q(n4778) );
  xor2s3 U3962 ( .DIN1(n6325), .DIN2(n6696), .Q(n4776) );
  nnd2s3 U3963 ( .DIN1(n6594), .DIN2(n1789), .Q(n4774) );
  nnd2s3 U3964 ( .DIN1(DATA_0_28), .DIN2(n6636), .Q(n4773) );
  nnd2s3 U3965 ( .DIN1(n6563), .DIN2(n1732), .Q(n4772) );
  nnd4s2 U3966 ( .DIN1(n4779), .DIN2(n4780), .DIN3(n4781), .DIN4(n4782), .Q(
        WX10992) );
  nnd2s3 U3967 ( .DIN1(n2491), .DIN2(n6667), .Q(n4782) );
  xor2s3 U3968 ( .DIN1(n4783), .DIN2(n4784), .Q(n2491) );
  xor2s3 U3969 ( .DIN1(n6329), .DIN2(n4785), .Q(n4784) );
  xor2s3 U3970 ( .DIN1(n6327), .DIN2(n6328), .Q(n4785) );
  xor2s3 U3971 ( .DIN1(n6330), .DIN2(n6696), .Q(n4783) );
  nnd2s3 U3972 ( .DIN1(n6594), .DIN2(n1790), .Q(n4781) );
  nnd2s3 U3973 ( .DIN1(DATA_0_29), .DIN2(n6636), .Q(n4780) );
  nnd2s3 U3974 ( .DIN1(n6563), .DIN2(n1731), .Q(n4779) );
  nnd4s2 U3975 ( .DIN1(n4786), .DIN2(n4787), .DIN3(n4788), .DIN4(n4789), .Q(
        WX10990) );
  nnd2s3 U3976 ( .DIN1(n2497), .DIN2(n6672), .Q(n4789) );
  xor2s3 U3977 ( .DIN1(n4790), .DIN2(n4791), .Q(n2497) );
  xor2s3 U3978 ( .DIN1(n6334), .DIN2(n4792), .Q(n4791) );
  xor2s3 U3979 ( .DIN1(n6332), .DIN2(n6333), .Q(n4792) );
  xor2s3 U3980 ( .DIN1(n6335), .DIN2(n6696), .Q(n4790) );
  nnd2s3 U3981 ( .DIN1(n6594), .DIN2(n1791), .Q(n4788) );
  nnd2s3 U3982 ( .DIN1(DATA_0_30), .DIN2(n6641), .Q(n4787) );
  nnd2s3 U3983 ( .DIN1(n6563), .DIN2(n1730), .Q(n4786) );
  nnd4s2 U3984 ( .DIN1(n4793), .DIN2(n4794), .DIN3(n4795), .DIN4(n4796), .Q(
        WX10988) );
  nnd2s3 U3985 ( .DIN1(n6594), .DIN2(n1792), .Q(n4796) );
  and3s3 U3986 ( .DIN1(TM1), .DIN2(RESET), .DIN3(n6703), .Q(n2316) );
  nnd2s3 U3987 ( .DIN1(DATA_0_31), .DIN2(n6625), .Q(n4795) );
  and3s3 U3988 ( .DIN1(n6711), .DIN2(n6698), .DIN3(RESET), .Q(n2314) );
  nnd2s3 U3989 ( .DIN1(n6563), .DIN2(n1729), .Q(n4794) );
  and3s3 U3990 ( .DIN1(RESET), .DIN2(n6698), .DIN3(n6703), .Q(n2317) );
  nnd2s3 U3991 ( .DIN1(n2503), .DIN2(n6661), .Q(n4793) );
  and3s3 U3992 ( .DIN1(RESET), .DIN2(n6711), .DIN3(TM1), .Q(n2312) );
  xor2s3 U3993 ( .DIN1(n4797), .DIN2(n4798), .Q(n2503) );
  xor2s3 U3994 ( .DIN1(n6340), .DIN2(n4799), .Q(n4798) );
  xor2s3 U3995 ( .DIN1(n6338), .DIN2(n6339), .Q(n4799) );
  xor2s3 U3996 ( .DIN1(n6341), .DIN2(n6696), .Q(n4797) );
  nor2s3 U3997 ( .DIN1(n6789), .DIN2(n1792), .Q(WX10890) );
  nor2s3 U3998 ( .DIN1(n6344), .DIN2(n6768), .Q(WX10888) );
  nor2s3 U3999 ( .DIN1(n6345), .DIN2(n6768), .Q(WX10886) );
  nor2s3 U4000 ( .DIN1(n6346), .DIN2(n6768), .Q(WX10884) );
  nor2s3 U4001 ( .DIN1(n6347), .DIN2(n6768), .Q(WX10882) );
  nor2s3 U4002 ( .DIN1(n6348), .DIN2(n6768), .Q(WX10880) );
  nor2s3 U4003 ( .DIN1(n6349), .DIN2(n6768), .Q(WX10878) );
  nor2s3 U4004 ( .DIN1(n6350), .DIN2(n6768), .Q(WX10876) );
  nor2s3 U4005 ( .DIN1(n6351), .DIN2(n6768), .Q(WX10874) );
  nor2s3 U4006 ( .DIN1(n6352), .DIN2(n6768), .Q(WX10872) );
  nor2s3 U4007 ( .DIN1(n6353), .DIN2(n6768), .Q(WX10870) );
  nor2s3 U4008 ( .DIN1(n6355), .DIN2(n6768), .Q(WX10868) );
  nor2s3 U4009 ( .DIN1(n6356), .DIN2(n6767), .Q(WX10866) );
  nor2s3 U4010 ( .DIN1(n6357), .DIN2(n6767), .Q(WX10864) );
  nor2s3 U4011 ( .DIN1(n6358), .DIN2(n6767), .Q(WX10862) );
  nor2s3 U4012 ( .DIN1(n6359), .DIN2(n6767), .Q(WX10860) );
  nor2s3 U4013 ( .DIN1(n6360), .DIN2(n6767), .Q(WX10858) );
  nor2s3 U4014 ( .DIN1(n6361), .DIN2(n6767), .Q(WX10856) );
  nor2s3 U4015 ( .DIN1(n6362), .DIN2(n6767), .Q(WX10854) );
  nor2s3 U4016 ( .DIN1(n6363), .DIN2(n6767), .Q(WX10852) );
  nor2s3 U4017 ( .DIN1(n6364), .DIN2(n6767), .Q(WX10850) );
  nor2s3 U4018 ( .DIN1(n6365), .DIN2(n6767), .Q(WX10848) );
  nor2s3 U4019 ( .DIN1(n6366), .DIN2(n6767), .Q(WX10846) );
  nor2s3 U4020 ( .DIN1(n6367), .DIN2(n6767), .Q(WX10844) );
  nor2s3 U4021 ( .DIN1(n6368), .DIN2(n6766), .Q(WX10842) );
  nor2s3 U4022 ( .DIN1(n6369), .DIN2(n6766), .Q(WX10840) );
  nor2s3 U4023 ( .DIN1(n6370), .DIN2(n6766), .Q(WX10838) );
  nor2s3 U4024 ( .DIN1(n6371), .DIN2(n6766), .Q(WX10836) );
  nor2s3 U4025 ( .DIN1(n6372), .DIN2(n6766), .Q(WX10834) );
  nor2s3 U4026 ( .DIN1(n6373), .DIN2(n6766), .Q(WX10832) );
  nor2s3 U4027 ( .DIN1(n6374), .DIN2(n6766), .Q(WX10830) );
  nor2s3 U4028 ( .DIN1(n6375), .DIN2(n6766), .Q(WX10828) );
  nor2s3 U4029 ( .DIN1(n6795), .DIN2(n4800), .Q(WX10377) );
  xor2s3 U4030 ( .DIN1(n6383), .DIN2(n6384), .Q(n4800) );
  nor2s3 U4031 ( .DIN1(n6795), .DIN2(n4801), .Q(WX10375) );
  xor2s3 U4032 ( .DIN1(n6385), .DIN2(n6386), .Q(n4801) );
  nor2s3 U4033 ( .DIN1(n6795), .DIN2(n4802), .Q(WX10373) );
  xor2s3 U4034 ( .DIN1(n6387), .DIN2(n6388), .Q(n4802) );
  nor2s3 U4035 ( .DIN1(n6795), .DIN2(n4803), .Q(WX10371) );
  xor2s3 U4036 ( .DIN1(n6389), .DIN2(n6390), .Q(n4803) );
  nor2s3 U4037 ( .DIN1(n6794), .DIN2(n4804), .Q(WX10369) );
  xor2s3 U4038 ( .DIN1(n6391), .DIN2(n6392), .Q(n4804) );
  nor2s3 U4039 ( .DIN1(n6794), .DIN2(n4805), .Q(WX10367) );
  xor2s3 U4040 ( .DIN1(n6393), .DIN2(n6394), .Q(n4805) );
  nor2s3 U4041 ( .DIN1(n6794), .DIN2(n4806), .Q(WX10365) );
  xor2s3 U4042 ( .DIN1(n6395), .DIN2(n6396), .Q(n4806) );
  nor2s3 U4043 ( .DIN1(n6794), .DIN2(n4807), .Q(WX10363) );
  xor2s3 U4044 ( .DIN1(n6397), .DIN2(n6398), .Q(n4807) );
  nor2s3 U4045 ( .DIN1(n6794), .DIN2(n4808), .Q(WX10361) );
  xor2s3 U4046 ( .DIN1(n6399), .DIN2(n6400), .Q(n4808) );
  nor2s3 U4047 ( .DIN1(n6794), .DIN2(n4809), .Q(WX10359) );
  xor2s3 U4048 ( .DIN1(n6401), .DIN2(n6402), .Q(n4809) );
  nor2s3 U4049 ( .DIN1(n6794), .DIN2(n4810), .Q(WX10357) );
  xor2s3 U4050 ( .DIN1(n6403), .DIN2(n6404), .Q(n4810) );
  nor2s3 U4051 ( .DIN1(n6794), .DIN2(n4811), .Q(WX10355) );
  xor2s3 U4052 ( .DIN1(n6405), .DIN2(n6406), .Q(n4811) );
  nor2s3 U4053 ( .DIN1(n6794), .DIN2(n4812), .Q(WX10353) );
  xor2s3 U4054 ( .DIN1(n6407), .DIN2(n6408), .Q(n4812) );
  nor2s3 U4055 ( .DIN1(n6793), .DIN2(n4813), .Q(WX10351) );
  xor2s3 U4056 ( .DIN1(n6409), .DIN2(n6410), .Q(n4813) );
  nor2s3 U4057 ( .DIN1(n6793), .DIN2(n4814), .Q(WX10349) );
  xor2s3 U4058 ( .DIN1(n6411), .DIN2(n6412), .Q(n4814) );
  nor2s3 U4059 ( .DIN1(n4815), .DIN2(n6766), .Q(WX10347) );
  xor2s3 U4060 ( .DIN1(n1793), .DIN2(n4816), .Q(n4815) );
  xor2s3 U4061 ( .DIN1(n6413), .DIN2(n6414), .Q(n4816) );
  nor2s3 U4062 ( .DIN1(n6793), .DIN2(n4817), .Q(WX10345) );
  xor2s3 U4063 ( .DIN1(n6415), .DIN2(n3220), .Q(n4817) );
  nor2s3 U4064 ( .DIN1(n6793), .DIN2(n4818), .Q(WX10343) );
  xor2s3 U4065 ( .DIN1(n6416), .DIN2(n3219), .Q(n4818) );
  nor2s3 U4066 ( .DIN1(n6792), .DIN2(n4819), .Q(WX10341) );
  xor2s3 U4067 ( .DIN1(n6417), .DIN2(n3218), .Q(n4819) );
  nor2s3 U4068 ( .DIN1(n6792), .DIN2(n4820), .Q(WX10339) );
  xor2s3 U4069 ( .DIN1(n6418), .DIN2(n3217), .Q(n4820) );
  nor2s3 U4070 ( .DIN1(n4821), .DIN2(n6766), .Q(WX10337) );
  xnr2s3 U4071 ( .DIN1(n3216), .DIN2(n4822), .Q(n4821) );
  xor2s3 U4072 ( .DIN1(n6419), .DIN2(n6430), .Q(n4822) );
  nor2s3 U4073 ( .DIN1(n6791), .DIN2(n4823), .Q(WX10335) );
  xor2s3 U4074 ( .DIN1(n6420), .DIN2(n3215), .Q(n4823) );
  nor2s3 U4075 ( .DIN1(n6791), .DIN2(n4824), .Q(WX10333) );
  xor2s3 U4076 ( .DIN1(n6421), .DIN2(n3214), .Q(n4824) );
  nor2s3 U4077 ( .DIN1(n6791), .DIN2(n4825), .Q(WX10331) );
  xor2s3 U4078 ( .DIN1(n6422), .DIN2(n3213), .Q(n4825) );
  nor2s3 U4079 ( .DIN1(n6791), .DIN2(n4826), .Q(WX10329) );
  xor2s3 U4080 ( .DIN1(n6423), .DIN2(n3212), .Q(n4826) );
  nor2s3 U4081 ( .DIN1(n6791), .DIN2(n4827), .Q(WX10327) );
  xor2s3 U4082 ( .DIN1(n6424), .DIN2(n3211), .Q(n4827) );
  nor2s3 U4083 ( .DIN1(n6791), .DIN2(n4828), .Q(WX10325) );
  xor2s3 U4084 ( .DIN1(n6425), .DIN2(n3210), .Q(n4828) );
  nor2s3 U4085 ( .DIN1(n4829), .DIN2(n6771), .Q(WX10323) );
  xnr2s3 U4086 ( .DIN1(n3209), .DIN2(n4830), .Q(n4829) );
  xor2s3 U4087 ( .DIN1(n6426), .DIN2(n6430), .Q(n4830) );
  nor2s3 U4088 ( .DIN1(n6791), .DIN2(n4831), .Q(WX10321) );
  xor2s3 U4089 ( .DIN1(n6427), .DIN2(n3208), .Q(n4831) );
  nor2s3 U4090 ( .DIN1(n6790), .DIN2(n4832), .Q(WX10319) );
  xor2s3 U4091 ( .DIN1(n6428), .DIN2(n3207), .Q(n4832) );
  nor2s3 U4092 ( .DIN1(n6788), .DIN2(n4833), .Q(WX10317) );
  xor2s3 U4093 ( .DIN1(n6429), .DIN2(n3206), .Q(n4833) );
  nor2s3 U4094 ( .DIN1(n6788), .DIN2(n4834), .Q(WX10315) );
  xor2s3 U4095 ( .DIN1(n6430), .DIN2(n3205), .Q(n4834) );
  xnr2s3 U4096 ( .DIN1(n4835), .DIN2(n3113), .Q(DATA_9_9) );
  xnr2s3 U4097 ( .DIN1(n4836), .DIN2(n4837), .Q(n3113) );
  xor2s3 U4098 ( .DIN1(n6506), .DIN2(n4838), .Q(n4837) );
  xor2s3 U4099 ( .DIN1(n6504), .DIN2(n6505), .Q(n4838) );
  xor2s3 U4100 ( .DIN1(n6507), .DIN2(n6710), .Q(n4836) );
  nnd2s3 U4101 ( .DIN1(n6703), .DIN2(n2282), .Q(n4835) );
  xnr2s3 U4102 ( .DIN1(n4839), .DIN2(n3107), .Q(DATA_9_8) );
  xnr2s3 U4103 ( .DIN1(n4840), .DIN2(n4841), .Q(n3107) );
  xor2s3 U4104 ( .DIN1(n6455), .DIN2(n4842), .Q(n4841) );
  xor2s3 U4105 ( .DIN1(n6453), .DIN2(n6454), .Q(n4842) );
  xor2s3 U4106 ( .DIN1(n6556), .DIN2(n6710), .Q(n4840) );
  nnd2s3 U4107 ( .DIN1(n6703), .DIN2(n2281), .Q(n4839) );
  xnr2s3 U4108 ( .DIN1(n4843), .DIN2(n3101), .Q(DATA_9_7) );
  xnr2s3 U4109 ( .DIN1(n4844), .DIN2(n4845), .Q(n3101) );
  xor2s3 U4110 ( .DIN1(n6467), .DIN2(n4846), .Q(n4845) );
  xor2s3 U4111 ( .DIN1(n6465), .DIN2(n6466), .Q(n4846) );
  xor2s3 U4112 ( .DIN1(n6552), .DIN2(n6710), .Q(n4844) );
  nnd2s3 U4113 ( .DIN1(n6703), .DIN2(n2280), .Q(n4843) );
  xnr2s3 U4114 ( .DIN1(n4847), .DIN2(n3095), .Q(DATA_9_6) );
  xnr2s3 U4115 ( .DIN1(n4848), .DIN2(n4849), .Q(n3095) );
  xor2s3 U4116 ( .DIN1(n6443), .DIN2(n4850), .Q(n4849) );
  xor2s3 U4117 ( .DIN1(n6441), .DIN2(n6442), .Q(n4850) );
  xor2s3 U4118 ( .DIN1(n6560), .DIN2(n6710), .Q(n4848) );
  nnd2s3 U4119 ( .DIN1(n6703), .DIN2(n2279), .Q(n4847) );
  xnr2s3 U4120 ( .DIN1(n4851), .DIN2(n3089), .Q(DATA_9_5) );
  xnr2s3 U4121 ( .DIN1(n4852), .DIN2(n4853), .Q(n3089) );
  xor2s3 U4122 ( .DIN1(n6461), .DIN2(n4854), .Q(n4853) );
  xor2s3 U4123 ( .DIN1(n6459), .DIN2(n6460), .Q(n4854) );
  xor2s3 U4124 ( .DIN1(n6554), .DIN2(n6709), .Q(n4852) );
  nnd2s3 U4125 ( .DIN1(n6703), .DIN2(n2278), .Q(n4851) );
  xnr2s3 U4126 ( .DIN1(n4855), .DIN2(n3083), .Q(DATA_9_4) );
  xnr2s3 U4127 ( .DIN1(n4856), .DIN2(n4857), .Q(n3083) );
  xor2s3 U4128 ( .DIN1(n6473), .DIN2(n4858), .Q(n4857) );
  xor2s3 U4129 ( .DIN1(n6471), .DIN2(n6472), .Q(n4858) );
  xor2s3 U4130 ( .DIN1(n6550), .DIN2(n6709), .Q(n4856) );
  nnd2s3 U4131 ( .DIN1(n6703), .DIN2(n2277), .Q(n4855) );
  xnr2s3 U4132 ( .DIN1(n4859), .DIN2(n3406), .Q(DATA_9_31) );
  xnr2s3 U4133 ( .DIN1(n4860), .DIN2(n4861), .Q(n3406) );
  xor2s3 U4134 ( .DIN1(n6533), .DIN2(n4862), .Q(n4861) );
  xor2s3 U4135 ( .DIN1(n6531), .DIN2(n6532), .Q(n4862) );
  xor2s3 U4136 ( .DIN1(n6534), .DIN2(n6696), .Q(n4860) );
  nnd2s3 U4137 ( .DIN1(n6703), .DIN2(n2304), .Q(n4859) );
  xnr2s3 U4138 ( .DIN1(n4863), .DIN2(n3388), .Q(DATA_9_30) );
  xnr2s3 U4139 ( .DIN1(n4864), .DIN2(n4865), .Q(n3388) );
  xor2s3 U4140 ( .DIN1(n6476), .DIN2(n4866), .Q(n4865) );
  xor2s3 U4141 ( .DIN1(n6474), .DIN2(n6475), .Q(n4866) );
  xor2s3 U4142 ( .DIN1(n6549), .DIN2(n6697), .Q(n4864) );
  nnd2s3 U4143 ( .DIN1(n6703), .DIN2(n2303), .Q(n4863) );
  xnr2s3 U4144 ( .DIN1(n4867), .DIN2(n3077), .Q(DATA_9_3) );
  xnr2s3 U4145 ( .DIN1(n4868), .DIN2(n4869), .Q(n3077) );
  xor2s3 U4146 ( .DIN1(n6470), .DIN2(n4870), .Q(n4869) );
  xor2s3 U4147 ( .DIN1(n6468), .DIN2(n6469), .Q(n4870) );
  xor2s3 U4148 ( .DIN1(n6551), .DIN2(n6709), .Q(n4868) );
  nnd2s3 U4149 ( .DIN1(n6703), .DIN2(n2276), .Q(n4867) );
  xnr2s3 U4150 ( .DIN1(n4871), .DIN2(n3371), .Q(DATA_9_29) );
  xnr2s3 U4151 ( .DIN1(n4872), .DIN2(n4873), .Q(n3371) );
  xor2s3 U4152 ( .DIN1(n6482), .DIN2(n4874), .Q(n4873) );
  xor2s3 U4153 ( .DIN1(n6480), .DIN2(n6481), .Q(n4874) );
  xor2s3 U4154 ( .DIN1(n6547), .DIN2(n6697), .Q(n4872) );
  nnd2s3 U4155 ( .DIN1(n6703), .DIN2(n2302), .Q(n4871) );
  xnr2s3 U4156 ( .DIN1(n4875), .DIN2(n3355), .Q(DATA_9_28) );
  xnr2s3 U4157 ( .DIN1(n4876), .DIN2(n4877), .Q(n3355) );
  xor2s3 U4158 ( .DIN1(n6485), .DIN2(n4878), .Q(n4877) );
  xor2s3 U4159 ( .DIN1(n6483), .DIN2(n6484), .Q(n4878) );
  xor2s3 U4160 ( .DIN1(n6546), .DIN2(n6697), .Q(n4876) );
  nnd2s3 U4161 ( .DIN1(n6703), .DIN2(n2301), .Q(n4875) );
  xnr2s3 U4162 ( .DIN1(n4879), .DIN2(n3349), .Q(DATA_9_27) );
  xnr2s3 U4163 ( .DIN1(n4880), .DIN2(n4881), .Q(n3349) );
  xor2s3 U4164 ( .DIN1(n6488), .DIN2(n4882), .Q(n4881) );
  xor2s3 U4165 ( .DIN1(n6486), .DIN2(n6487), .Q(n4882) );
  xor2s3 U4166 ( .DIN1(n6545), .DIN2(n6697), .Q(n4880) );
  nnd2s3 U4167 ( .DIN1(n6703), .DIN2(n2300), .Q(n4879) );
  xnr2s3 U4168 ( .DIN1(n4883), .DIN2(n3343), .Q(DATA_9_26) );
  xnr2s3 U4169 ( .DIN1(n4884), .DIN2(n4885), .Q(n3343) );
  xor2s3 U4170 ( .DIN1(n6494), .DIN2(n4886), .Q(n4885) );
  xor2s3 U4171 ( .DIN1(n6492), .DIN2(n6493), .Q(n4886) );
  xor2s3 U4172 ( .DIN1(n6543), .DIN2(n6697), .Q(n4884) );
  nnd2s3 U4173 ( .DIN1(n6703), .DIN2(n2299), .Q(n4883) );
  xnr2s3 U4174 ( .DIN1(n4887), .DIN2(n3337), .Q(DATA_9_25) );
  xnr2s3 U4175 ( .DIN1(n4888), .DIN2(n4889), .Q(n3337) );
  xor2s3 U4176 ( .DIN1(n6500), .DIN2(n4890), .Q(n4889) );
  xor2s3 U4177 ( .DIN1(n6498), .DIN2(n6499), .Q(n4890) );
  xor2s3 U4178 ( .DIN1(n6541), .DIN2(n6697), .Q(n4888) );
  nnd2s3 U4179 ( .DIN1(n6704), .DIN2(n2298), .Q(n4887) );
  xnr2s3 U4180 ( .DIN1(n4891), .DIN2(n3203), .Q(DATA_9_24) );
  xnr2s3 U4181 ( .DIN1(n4892), .DIN2(n4893), .Q(n3203) );
  xor2s3 U4182 ( .DIN1(n6503), .DIN2(n4894), .Q(n4893) );
  xor2s3 U4183 ( .DIN1(n6501), .DIN2(n6502), .Q(n4894) );
  xor2s3 U4184 ( .DIN1(n6540), .DIN2(n6697), .Q(n4892) );
  nnd2s3 U4185 ( .DIN1(n6704), .DIN2(n2297), .Q(n4891) );
  xnr2s3 U4186 ( .DIN1(n4895), .DIN2(n3197), .Q(DATA_9_23) );
  xnr2s3 U4187 ( .DIN1(n4896), .DIN2(n4897), .Q(n3197) );
  xor2s3 U4188 ( .DIN1(n6513), .DIN2(n4898), .Q(n4897) );
  xor2s3 U4189 ( .DIN1(n6511), .DIN2(n6512), .Q(n4898) );
  xor2s3 U4190 ( .DIN1(n6538), .DIN2(n6697), .Q(n4896) );
  nnd2s3 U4191 ( .DIN1(n6704), .DIN2(n2296), .Q(n4895) );
  xnr2s3 U4192 ( .DIN1(n4899), .DIN2(n3191), .Q(DATA_9_22) );
  xnr2s3 U4193 ( .DIN1(n4900), .DIN2(n4901), .Q(n3191) );
  xor2s3 U4194 ( .DIN1(n6516), .DIN2(n4902), .Q(n4901) );
  xor2s3 U4195 ( .DIN1(n6514), .DIN2(n6515), .Q(n4902) );
  xor2s3 U4196 ( .DIN1(n6537), .DIN2(n6697), .Q(n4900) );
  nnd2s3 U4197 ( .DIN1(n6704), .DIN2(n2295), .Q(n4899) );
  xnr2s3 U4198 ( .DIN1(n4903), .DIN2(n3185), .Q(DATA_9_21) );
  xnr2s3 U4199 ( .DIN1(n4904), .DIN2(n4905), .Q(n3185) );
  xor2s3 U4200 ( .DIN1(n6519), .DIN2(n4906), .Q(n4905) );
  xor2s3 U4201 ( .DIN1(n6517), .DIN2(n6518), .Q(n4906) );
  xor2s3 U4202 ( .DIN1(n6536), .DIN2(n6697), .Q(n4904) );
  nnd2s3 U4203 ( .DIN1(n6704), .DIN2(n2294), .Q(n4903) );
  xnr2s3 U4204 ( .DIN1(n4907), .DIN2(n3179), .Q(DATA_9_20) );
  xnr2s3 U4205 ( .DIN1(n4908), .DIN2(n4909), .Q(n3179) );
  xor2s3 U4206 ( .DIN1(n6522), .DIN2(n4910), .Q(n4909) );
  xor2s3 U4207 ( .DIN1(n6520), .DIN2(n6521), .Q(n4910) );
  xor2s3 U4208 ( .DIN1(n6535), .DIN2(n6697), .Q(n4908) );
  nnd2s3 U4209 ( .DIN1(n6704), .DIN2(n2293), .Q(n4907) );
  xnr2s3 U4210 ( .DIN1(n4911), .DIN2(n3071), .Q(DATA_9_2) );
  xnr2s3 U4211 ( .DIN1(n4912), .DIN2(n4913), .Q(n3071) );
  xor2s3 U4212 ( .DIN1(n6437), .DIN2(n4914), .Q(n4913) );
  xor2s3 U4213 ( .DIN1(n6435), .DIN2(n6436), .Q(n4914) );
  xor2s3 U4214 ( .DIN1(n6562), .DIN2(n6709), .Q(n4912) );
  nnd2s3 U4215 ( .DIN1(n6704), .DIN2(n2275), .Q(n4911) );
  xnr2s3 U4216 ( .DIN1(n4915), .DIN2(n3173), .Q(DATA_9_19) );
  xnr2s3 U4217 ( .DIN1(n4916), .DIN2(n4917), .Q(n3173) );
  xor2s3 U4218 ( .DIN1(n6479), .DIN2(n4918), .Q(n4917) );
  xor2s3 U4219 ( .DIN1(n6477), .DIN2(n6478), .Q(n4918) );
  xor2s3 U4220 ( .DIN1(n6548), .DIN2(n6697), .Q(n4916) );
  nnd2s3 U4221 ( .DIN1(n6704), .DIN2(n2292), .Q(n4915) );
  xnr2s3 U4222 ( .DIN1(n4919), .DIN2(n3167), .Q(DATA_9_18) );
  xnr2s3 U4223 ( .DIN1(n4920), .DIN2(n4921), .Q(n3167) );
  xor2s3 U4224 ( .DIN1(n6491), .DIN2(n4922), .Q(n4921) );
  xor2s3 U4225 ( .DIN1(n6489), .DIN2(n6490), .Q(n4922) );
  xor2s3 U4226 ( .DIN1(n6544), .DIN2(n6698), .Q(n4920) );
  nnd2s3 U4227 ( .DIN1(n6704), .DIN2(n2291), .Q(n4919) );
  xnr2s3 U4228 ( .DIN1(n4923), .DIN2(n3161), .Q(DATA_9_17) );
  xnr2s3 U4229 ( .DIN1(n4924), .DIN2(n4925), .Q(n3161) );
  xor2s3 U4230 ( .DIN1(n6497), .DIN2(n4926), .Q(n4925) );
  xor2s3 U4231 ( .DIN1(n6495), .DIN2(n6496), .Q(n4926) );
  xor2s3 U4232 ( .DIN1(n6542), .DIN2(n6697), .Q(n4924) );
  nnd2s3 U4233 ( .DIN1(n6704), .DIN2(n2290), .Q(n4923) );
  xnr2s3 U4234 ( .DIN1(n4927), .DIN2(n3155), .Q(DATA_9_16) );
  xnr2s3 U4235 ( .DIN1(n4928), .DIN2(n4929), .Q(n3155) );
  xor2s3 U4236 ( .DIN1(n6510), .DIN2(n4930), .Q(n4929) );
  xor2s3 U4237 ( .DIN1(n6508), .DIN2(n6509), .Q(n4930) );
  xor2s3 U4238 ( .DIN1(n6539), .DIN2(n6687), .Q(n4928) );
  nnd2s3 U4239 ( .DIN1(n6704), .DIN2(n2289), .Q(n4927) );
  xnr2s3 U4240 ( .DIN1(n4931), .DIN2(n3149), .Q(DATA_9_15) );
  xnr2s3 U4241 ( .DIN1(n4932), .DIN2(n4933), .Q(n3149) );
  xor2s3 U4242 ( .DIN1(n6440), .DIN2(n4934), .Q(n4933) );
  xor2s3 U4243 ( .DIN1(n6438), .DIN2(n6439), .Q(n4934) );
  xor2s3 U4244 ( .DIN1(n6561), .DIN2(n6708), .Q(n4932) );
  nnd2s3 U4245 ( .DIN1(n6704), .DIN2(n2288), .Q(n4931) );
  xnr2s3 U4246 ( .DIN1(n4935), .DIN2(n3143), .Q(DATA_9_14) );
  xnr2s3 U4247 ( .DIN1(n4936), .DIN2(n4937), .Q(n3143) );
  xor2s3 U4248 ( .DIN1(n6525), .DIN2(n4938), .Q(n4937) );
  xor2s3 U4249 ( .DIN1(n6523), .DIN2(n6524), .Q(n4938) );
  xor2s3 U4250 ( .DIN1(n6526), .DIN2(n6708), .Q(n4936) );
  nnd2s3 U4251 ( .DIN1(n6704), .DIN2(n2287), .Q(n4935) );
  xnr2s3 U4252 ( .DIN1(n4939), .DIN2(n3137), .Q(DATA_9_13) );
  xnr2s3 U4253 ( .DIN1(n4940), .DIN2(n4941), .Q(n3137) );
  xor2s3 U4254 ( .DIN1(n6449), .DIN2(n4942), .Q(n4941) );
  xor2s3 U4255 ( .DIN1(n6447), .DIN2(n6448), .Q(n4942) );
  xor2s3 U4256 ( .DIN1(n6558), .DIN2(n6708), .Q(n4940) );
  nnd2s3 U4257 ( .DIN1(n6704), .DIN2(n2286), .Q(n4939) );
  xnr2s3 U4258 ( .DIN1(n4943), .DIN2(n3131), .Q(DATA_9_12) );
  xnr2s3 U4259 ( .DIN1(n4944), .DIN2(n4945), .Q(n3131) );
  xor2s3 U4260 ( .DIN1(n6458), .DIN2(n4946), .Q(n4945) );
  xor2s3 U4261 ( .DIN1(n6456), .DIN2(n6457), .Q(n4946) );
  xor2s3 U4262 ( .DIN1(n6555), .DIN2(n6708), .Q(n4944) );
  nnd2s3 U4263 ( .DIN1(n6704), .DIN2(n2285), .Q(n4943) );
  xnr2s3 U4264 ( .DIN1(n4947), .DIN2(n3125), .Q(DATA_9_11) );
  xnr2s3 U4265 ( .DIN1(n4948), .DIN2(n4949), .Q(n3125) );
  xor2s3 U4266 ( .DIN1(n6446), .DIN2(n4950), .Q(n4949) );
  xor2s3 U4267 ( .DIN1(n6444), .DIN2(n6445), .Q(n4950) );
  xor2s3 U4268 ( .DIN1(n6559), .DIN2(n6707), .Q(n4948) );
  nnd2s3 U4269 ( .DIN1(n6704), .DIN2(n2284), .Q(n4947) );
  xnr2s3 U4270 ( .DIN1(n4951), .DIN2(n3119), .Q(DATA_9_10) );
  xnr2s3 U4271 ( .DIN1(n4952), .DIN2(n4953), .Q(n3119) );
  xor2s3 U4272 ( .DIN1(n6452), .DIN2(n4954), .Q(n4953) );
  xor2s3 U4273 ( .DIN1(n6450), .DIN2(n6451), .Q(n4954) );
  xor2s3 U4274 ( .DIN1(n6557), .DIN2(n6707), .Q(n4952) );
  nnd2s3 U4275 ( .DIN1(n6705), .DIN2(n2283), .Q(n4951) );
  xnr2s3 U4276 ( .DIN1(n4955), .DIN2(n3065), .Q(DATA_9_1) );
  xnr2s3 U4277 ( .DIN1(n4956), .DIN2(n4957), .Q(n3065) );
  xor2s3 U4278 ( .DIN1(n6529), .DIN2(n4958), .Q(n4957) );
  xor2s3 U4279 ( .DIN1(n6527), .DIN2(n6528), .Q(n4958) );
  xor2s3 U4280 ( .DIN1(n6530), .DIN2(n6707), .Q(n4956) );
  nnd2s3 U4281 ( .DIN1(n6705), .DIN2(n2274), .Q(n4955) );
  xnr2s3 U4282 ( .DIN1(n4959), .DIN2(n3059), .Q(DATA_9_0) );
  xnr2s3 U4283 ( .DIN1(n4960), .DIN2(n4961), .Q(n3059) );
  xor2s3 U4284 ( .DIN1(n6464), .DIN2(n4962), .Q(n4961) );
  xor2s3 U4285 ( .DIN1(n6462), .DIN2(n6463), .Q(n4962) );
  xor2s3 U4286 ( .DIN1(n6553), .DIN2(n6707), .Q(n4960) );
  nnd2s3 U4287 ( .DIN1(n6705), .DIN2(n2273), .Q(n4959) );
  i1s3 U4288 ( .DIN(n6337), .Q(n1729) );
  i1s3 U4289 ( .DIN(n6336), .Q(n1730) );
  i1s3 U4290 ( .DIN(n6331), .Q(n1731) );
  i1s3 U4291 ( .DIN(n6326), .Q(n1732) );
  i1s3 U4292 ( .DIN(n6321), .Q(n1733) );
  i1s3 U4293 ( .DIN(n6316), .Q(n1734) );
  i1s3 U4294 ( .DIN(n6311), .Q(n1735) );
  i1s3 U4295 ( .DIN(n6306), .Q(n1736) );
  i1s3 U4296 ( .DIN(n6301), .Q(n1737) );
  i1s3 U4297 ( .DIN(n6296), .Q(n1738) );
  i1s3 U4298 ( .DIN(n6291), .Q(n1739) );
  i1s3 U4299 ( .DIN(n6285), .Q(n1740) );
  i1s3 U4300 ( .DIN(n6280), .Q(n1741) );
  i1s3 U4301 ( .DIN(n6275), .Q(n1742) );
  i1s3 U4302 ( .DIN(n6270), .Q(n1743) );
  i1s3 U4303 ( .DIN(n6265), .Q(n1744) );
  i1s3 U4304 ( .DIN(n6260), .Q(n1745) );
  i1s3 U4305 ( .DIN(n6256), .Q(n1746) );
  i1s3 U4306 ( .DIN(n6252), .Q(n1747) );
  i1s3 U4307 ( .DIN(n6248), .Q(n1748) );
  i1s3 U4308 ( .DIN(n6244), .Q(n1749) );
  i1s3 U4309 ( .DIN(n6240), .Q(n1750) );
  i1s3 U4310 ( .DIN(n6236), .Q(n1751) );
  i1s3 U4311 ( .DIN(n6232), .Q(n1752) );
  i1s3 U4312 ( .DIN(n6228), .Q(n1753) );
  i1s3 U4313 ( .DIN(n6224), .Q(n1754) );
  i1s3 U4314 ( .DIN(n6220), .Q(n1755) );
  i1s3 U4315 ( .DIN(n6216), .Q(n1756) );
  i1s3 U4316 ( .DIN(n6212), .Q(n1757) );
  i1s3 U4317 ( .DIN(n6208), .Q(n1758) );
  i1s3 U4318 ( .DIN(n6204), .Q(n1759) );
  i1s3 U4319 ( .DIN(n6200), .Q(n1760) );
  i1s3 U4320 ( .DIN(n6344), .Q(n1761) );
  i1s3 U4321 ( .DIN(n6345), .Q(n1762) );
  i1s3 U4322 ( .DIN(n6346), .Q(n1763) );
  i1s3 U4323 ( .DIN(n6347), .Q(n1764) );
  i1s3 U4324 ( .DIN(n6348), .Q(n1765) );
  i1s3 U4325 ( .DIN(n6349), .Q(n1766) );
  i1s3 U4326 ( .DIN(n6350), .Q(n1767) );
  i1s3 U4327 ( .DIN(n6351), .Q(n1768) );
  i1s3 U4328 ( .DIN(n6352), .Q(n1769) );
  i1s3 U4329 ( .DIN(n6353), .Q(n1770) );
  i1s3 U4330 ( .DIN(n6355), .Q(n1771) );
  i1s3 U4331 ( .DIN(n6356), .Q(n1772) );
  i1s3 U4332 ( .DIN(n6357), .Q(n1773) );
  i1s3 U4333 ( .DIN(n6358), .Q(n1774) );
  i1s3 U4334 ( .DIN(n6359), .Q(n1775) );
  i1s3 U4335 ( .DIN(n6360), .Q(n1776) );
  i1s3 U4336 ( .DIN(n6361), .Q(n1777) );
  i1s3 U4337 ( .DIN(n6362), .Q(n1778) );
  i1s3 U4338 ( .DIN(n6363), .Q(n1779) );
  i1s3 U4339 ( .DIN(n6364), .Q(n1780) );
  i1s3 U4340 ( .DIN(n6365), .Q(n1781) );
  i1s3 U4341 ( .DIN(n6366), .Q(n1782) );
  i1s3 U4342 ( .DIN(n6367), .Q(n1783) );
  i1s3 U4343 ( .DIN(n6368), .Q(n1784) );
  i1s3 U4344 ( .DIN(n6369), .Q(n1785) );
  i1s3 U4345 ( .DIN(n6370), .Q(n1786) );
  i1s3 U4346 ( .DIN(n6371), .Q(n1787) );
  i1s3 U4347 ( .DIN(n6372), .Q(n1788) );
  i1s3 U4348 ( .DIN(n6373), .Q(n1789) );
  i1s3 U4349 ( .DIN(n6374), .Q(n1790) );
  i1s3 U4350 ( .DIN(n6375), .Q(n1791) );
  i1s3 U4351 ( .DIN(n6343), .Q(n1792) );
  i1s3 U4352 ( .DIN(n6430), .Q(n1793) );
  i1s3 U4353 ( .DIN(n6383), .Q(n1794) );
  i1s3 U4354 ( .DIN(n6385), .Q(n1795) );
  i1s3 U4355 ( .DIN(n6387), .Q(n1796) );
  i1s3 U4356 ( .DIN(n6389), .Q(n1797) );
  i1s3 U4357 ( .DIN(n6391), .Q(n1798) );
  i1s3 U4358 ( .DIN(n6393), .Q(n1799) );
  i1s3 U4359 ( .DIN(n6395), .Q(n1800) );
  i1s3 U4360 ( .DIN(n6397), .Q(n1801) );
  i1s3 U4361 ( .DIN(n6399), .Q(n1802) );
  i1s3 U4362 ( .DIN(n6401), .Q(n1803) );
  i1s3 U4363 ( .DIN(n6403), .Q(n1804) );
  i1s3 U4364 ( .DIN(n6405), .Q(n1805) );
  i1s3 U4365 ( .DIN(n6407), .Q(n1806) );
  i1s3 U4366 ( .DIN(n6409), .Q(n1807) );
  i1s3 U4367 ( .DIN(n6411), .Q(n1808) );
  i1s3 U4368 ( .DIN(n6413), .Q(n1809) );
  i1s3 U4369 ( .DIN(n6415), .Q(n1810) );
  i1s3 U4370 ( .DIN(n6416), .Q(n1811) );
  i1s3 U4371 ( .DIN(n6417), .Q(n1812) );
  i1s3 U4372 ( .DIN(n6418), .Q(n1813) );
  i1s3 U4373 ( .DIN(n6419), .Q(n1814) );
  i1s3 U4374 ( .DIN(n6420), .Q(n1815) );
  i1s3 U4375 ( .DIN(n6421), .Q(n1816) );
  i1s3 U4376 ( .DIN(n6422), .Q(n1817) );
  i1s3 U4377 ( .DIN(n6423), .Q(n1818) );
  i1s3 U4378 ( .DIN(n6424), .Q(n1819) );
  i1s3 U4379 ( .DIN(n6425), .Q(n1820) );
  i1s3 U4380 ( .DIN(n6426), .Q(n1821) );
  i1s3 U4381 ( .DIN(n6427), .Q(n1822) );
  i1s3 U4382 ( .DIN(n6428), .Q(n1823) );
  i1s3 U4383 ( .DIN(n6429), .Q(n1824) );
  i1s3 U4384 ( .DIN(n4964), .Q(n1825) );
  i1s3 U4385 ( .DIN(n4965), .Q(n1826) );
  i1s3 U4386 ( .DIN(n4966), .Q(n1827) );
  i1s3 U4387 ( .DIN(n4967), .Q(n1828) );
  i1s3 U4388 ( .DIN(n4968), .Q(n1829) );
  i1s3 U4389 ( .DIN(n4969), .Q(n1830) );
  i1s3 U4390 ( .DIN(n4970), .Q(n1831) );
  i1s3 U4391 ( .DIN(n4971), .Q(n1832) );
  i1s3 U4392 ( .DIN(n4972), .Q(n1833) );
  i1s3 U4393 ( .DIN(n4973), .Q(n1834) );
  i1s3 U4394 ( .DIN(n4974), .Q(n1835) );
  i1s3 U4395 ( .DIN(n4975), .Q(n1836) );
  i1s3 U4396 ( .DIN(n4976), .Q(n1837) );
  i1s3 U4397 ( .DIN(n4977), .Q(n1838) );
  i1s3 U4398 ( .DIN(n4978), .Q(n1839) );
  i1s3 U4399 ( .DIN(n4979), .Q(n1840) );
  i1s3 U4400 ( .DIN(n4980), .Q(n1841) );
  i1s3 U4401 ( .DIN(n4981), .Q(n1842) );
  i1s3 U4402 ( .DIN(n4982), .Q(n1843) );
  i1s3 U4403 ( .DIN(n4983), .Q(n1844) );
  i1s3 U4404 ( .DIN(n4984), .Q(n1845) );
  i1s3 U4405 ( .DIN(n4985), .Q(n1846) );
  i1s3 U4406 ( .DIN(n4986), .Q(n1847) );
  i1s3 U4407 ( .DIN(n4987), .Q(n1848) );
  i1s3 U4408 ( .DIN(n4988), .Q(n1849) );
  i1s3 U4409 ( .DIN(n4989), .Q(n1850) );
  i1s3 U4410 ( .DIN(n4990), .Q(n1851) );
  i1s3 U4411 ( .DIN(n4991), .Q(n1852) );
  i1s3 U4412 ( .DIN(n4992), .Q(n1853) );
  i1s3 U4413 ( .DIN(n4993), .Q(n1854) );
  i1s3 U4414 ( .DIN(n4994), .Q(n1855) );
  i1s3 U4415 ( .DIN(n4963), .Q(n1856) );
  i1s3 U4416 ( .DIN(n5122), .Q(n1857) );
  i1s3 U4417 ( .DIN(n5118), .Q(n1858) );
  i1s3 U4418 ( .DIN(n5114), .Q(n1859) );
  i1s3 U4419 ( .DIN(n5110), .Q(n1860) );
  i1s3 U4420 ( .DIN(n5106), .Q(n1861) );
  i1s3 U4421 ( .DIN(n5102), .Q(n1862) );
  i1s3 U4422 ( .DIN(n5098), .Q(n1863) );
  i1s3 U4423 ( .DIN(n5094), .Q(n1864) );
  i1s3 U4424 ( .DIN(n5090), .Q(n1865) );
  i1s3 U4425 ( .DIN(n5086), .Q(n1866) );
  i1s3 U4426 ( .DIN(n5082), .Q(n1867) );
  i1s3 U4427 ( .DIN(n5078), .Q(n1868) );
  i1s3 U4428 ( .DIN(n5074), .Q(n1869) );
  i1s3 U4429 ( .DIN(n5070), .Q(n1870) );
  i1s3 U4430 ( .DIN(n5066), .Q(n1871) );
  i1s3 U4431 ( .DIN(n5062), .Q(n1872) );
  i1s3 U4432 ( .DIN(n5058), .Q(n1873) );
  i1s3 U4433 ( .DIN(n5054), .Q(n1874) );
  i1s3 U4434 ( .DIN(n5050), .Q(n1875) );
  i1s3 U4435 ( .DIN(n5046), .Q(n1876) );
  i1s3 U4436 ( .DIN(n5042), .Q(n1877) );
  i1s3 U4437 ( .DIN(n5038), .Q(n1878) );
  i1s3 U4438 ( .DIN(n5034), .Q(n1879) );
  i1s3 U4439 ( .DIN(n5030), .Q(n1880) );
  i1s3 U4440 ( .DIN(n5026), .Q(n1881) );
  i1s3 U4441 ( .DIN(n5022), .Q(n1882) );
  i1s3 U4442 ( .DIN(n5018), .Q(n1883) );
  i1s3 U4443 ( .DIN(n5014), .Q(n1884) );
  i1s3 U4444 ( .DIN(n5010), .Q(n1885) );
  i1s3 U4445 ( .DIN(n5006), .Q(n1886) );
  i1s3 U4446 ( .DIN(n5002), .Q(n1887) );
  i1s3 U4447 ( .DIN(n4998), .Q(n1888) );
  i1s3 U4448 ( .DIN(n5124), .Q(n1889) );
  i1s3 U4449 ( .DIN(n5125), .Q(n1890) );
  i1s3 U4450 ( .DIN(n5126), .Q(n1891) );
  i1s3 U4451 ( .DIN(n5127), .Q(n1892) );
  i1s3 U4452 ( .DIN(n5128), .Q(n1893) );
  i1s3 U4453 ( .DIN(n5129), .Q(n1894) );
  i1s3 U4454 ( .DIN(n5130), .Q(n1895) );
  i1s3 U4455 ( .DIN(n5131), .Q(n1896) );
  i1s3 U4456 ( .DIN(n5132), .Q(n1897) );
  i1s3 U4457 ( .DIN(n5133), .Q(n1898) );
  i1s3 U4458 ( .DIN(n5134), .Q(n1899) );
  i1s3 U4459 ( .DIN(n5135), .Q(n1900) );
  i1s3 U4460 ( .DIN(n5136), .Q(n1901) );
  i1s3 U4461 ( .DIN(n5137), .Q(n1902) );
  i1s3 U4462 ( .DIN(n5138), .Q(n1903) );
  i1s3 U4463 ( .DIN(n5139), .Q(n1904) );
  i1s3 U4464 ( .DIN(n5140), .Q(n1905) );
  i1s3 U4465 ( .DIN(n5141), .Q(n1906) );
  i1s3 U4466 ( .DIN(n5142), .Q(n1907) );
  i1s3 U4467 ( .DIN(n5143), .Q(n1908) );
  i1s3 U4468 ( .DIN(n5144), .Q(n1909) );
  i1s3 U4469 ( .DIN(n5145), .Q(n1910) );
  i1s3 U4470 ( .DIN(n5146), .Q(n1911) );
  i1s3 U4471 ( .DIN(n5147), .Q(n1912) );
  i1s3 U4472 ( .DIN(n5148), .Q(n1913) );
  i1s3 U4473 ( .DIN(n5149), .Q(n1914) );
  i1s3 U4474 ( .DIN(n5150), .Q(n1915) );
  i1s3 U4475 ( .DIN(n5151), .Q(n1916) );
  i1s3 U4476 ( .DIN(n5152), .Q(n1917) );
  i1s3 U4477 ( .DIN(n5153), .Q(n1918) );
  i1s3 U4478 ( .DIN(n5154), .Q(n1919) );
  i1s3 U4479 ( .DIN(n5123), .Q(n1920) );
  i1s3 U4480 ( .DIN(n5298), .Q(n1921) );
  i1s3 U4481 ( .DIN(n5293), .Q(n1922) );
  i1s3 U4482 ( .DIN(n5288), .Q(n1923) );
  i1s3 U4483 ( .DIN(n5283), .Q(n1924) );
  i1s3 U4484 ( .DIN(n5278), .Q(n1925) );
  i1s3 U4485 ( .DIN(n5273), .Q(n1926) );
  i1s3 U4486 ( .DIN(n5268), .Q(n1927) );
  i1s3 U4487 ( .DIN(n5263), .Q(n1928) );
  i1s3 U4488 ( .DIN(n5258), .Q(n1929) );
  i1s3 U4489 ( .DIN(n5253), .Q(n1930) );
  i1s3 U4490 ( .DIN(n5248), .Q(n1931) );
  i1s3 U4491 ( .DIN(n5243), .Q(n1932) );
  i1s3 U4492 ( .DIN(n5238), .Q(n1933) );
  i1s3 U4493 ( .DIN(n5233), .Q(n1934) );
  i1s3 U4494 ( .DIN(n5228), .Q(n1935) );
  i1s3 U4495 ( .DIN(n5223), .Q(n1936) );
  i1s3 U4496 ( .DIN(n5218), .Q(n1937) );
  i1s3 U4497 ( .DIN(n5214), .Q(n1938) );
  i1s3 U4498 ( .DIN(n5210), .Q(n1939) );
  i1s3 U4499 ( .DIN(n5206), .Q(n1940) );
  i1s3 U4500 ( .DIN(n5202), .Q(n1941) );
  i1s3 U4501 ( .DIN(n5198), .Q(n1942) );
  i1s3 U4502 ( .DIN(n5194), .Q(n1943) );
  i1s3 U4503 ( .DIN(n5190), .Q(n1944) );
  i1s3 U4504 ( .DIN(n5186), .Q(n1945) );
  i1s3 U4505 ( .DIN(n5182), .Q(n1946) );
  i1s3 U4506 ( .DIN(n5178), .Q(n1947) );
  i1s3 U4507 ( .DIN(n5174), .Q(n1948) );
  i1s3 U4508 ( .DIN(n5170), .Q(n1949) );
  i1s3 U4509 ( .DIN(n5166), .Q(n1950) );
  i1s3 U4510 ( .DIN(n5162), .Q(n1951) );
  i1s3 U4511 ( .DIN(n5158), .Q(n1952) );
  i1s3 U4512 ( .DIN(n5300), .Q(n1953) );
  i1s3 U4513 ( .DIN(n5301), .Q(n1954) );
  i1s3 U4514 ( .DIN(n5302), .Q(n1955) );
  i1s3 U4515 ( .DIN(n5303), .Q(n1956) );
  i1s3 U4516 ( .DIN(n5304), .Q(n1957) );
  i1s3 U4517 ( .DIN(n5305), .Q(n1958) );
  i1s3 U4518 ( .DIN(n5306), .Q(n1959) );
  i1s3 U4519 ( .DIN(n5307), .Q(n1960) );
  i1s3 U4520 ( .DIN(n5308), .Q(n1961) );
  i1s3 U4521 ( .DIN(n5309), .Q(n1962) );
  i1s3 U4522 ( .DIN(n5310), .Q(n1963) );
  i1s3 U4523 ( .DIN(n5311), .Q(n1964) );
  i1s3 U4524 ( .DIN(n5312), .Q(n1965) );
  i1s3 U4525 ( .DIN(n5313), .Q(n1966) );
  i1s3 U4526 ( .DIN(n5314), .Q(n1967) );
  i1s3 U4527 ( .DIN(n5315), .Q(n1968) );
  i1s3 U4528 ( .DIN(n5316), .Q(n1969) );
  i1s3 U4529 ( .DIN(n5317), .Q(n1970) );
  i1s3 U4530 ( .DIN(n5318), .Q(n1971) );
  i1s3 U4531 ( .DIN(n5319), .Q(n1972) );
  i1s3 U4532 ( .DIN(n5320), .Q(n1973) );
  i1s3 U4533 ( .DIN(n5321), .Q(n1974) );
  i1s3 U4534 ( .DIN(n5322), .Q(n1975) );
  i1s3 U4535 ( .DIN(n5323), .Q(n1976) );
  i1s3 U4536 ( .DIN(n5324), .Q(n1977) );
  i1s3 U4537 ( .DIN(n5325), .Q(n1978) );
  i1s3 U4538 ( .DIN(n5326), .Q(n1979) );
  i1s3 U4539 ( .DIN(n5327), .Q(n1980) );
  i1s3 U4540 ( .DIN(n5328), .Q(n1981) );
  i1s3 U4541 ( .DIN(n5329), .Q(n1982) );
  i1s3 U4542 ( .DIN(n5330), .Q(n1983) );
  i1s3 U4543 ( .DIN(n5299), .Q(n1984) );
  i1s3 U4544 ( .DIN(n5474), .Q(n1985) );
  i1s3 U4545 ( .DIN(n5469), .Q(n1986) );
  i1s3 U4546 ( .DIN(n5464), .Q(n1987) );
  i1s3 U4547 ( .DIN(n5459), .Q(n1988) );
  i1s3 U4548 ( .DIN(n5454), .Q(n1989) );
  i1s3 U4549 ( .DIN(n5449), .Q(n1990) );
  i1s3 U4550 ( .DIN(n5444), .Q(n1991) );
  i1s3 U4551 ( .DIN(n5439), .Q(n1992) );
  i1s3 U4552 ( .DIN(n5434), .Q(n1993) );
  i1s3 U4553 ( .DIN(n5429), .Q(n1994) );
  i1s3 U4554 ( .DIN(n5424), .Q(n1995) );
  i1s3 U4555 ( .DIN(n5419), .Q(n1996) );
  i1s3 U4556 ( .DIN(n5414), .Q(n1997) );
  i1s3 U4557 ( .DIN(n5409), .Q(n1998) );
  i1s3 U4558 ( .DIN(n5404), .Q(n1999) );
  i1s3 U4559 ( .DIN(n5399), .Q(n2000) );
  i1s3 U4560 ( .DIN(n5394), .Q(n2001) );
  i1s3 U4561 ( .DIN(n5390), .Q(n2002) );
  i1s3 U4562 ( .DIN(n5386), .Q(n2003) );
  i1s3 U4563 ( .DIN(n5382), .Q(n2004) );
  i1s3 U4564 ( .DIN(n5378), .Q(n2005) );
  i1s3 U4565 ( .DIN(n5374), .Q(n2006) );
  i1s3 U4566 ( .DIN(n5370), .Q(n2007) );
  i1s3 U4567 ( .DIN(n5366), .Q(n2008) );
  i1s3 U4568 ( .DIN(n5362), .Q(n2009) );
  i1s3 U4569 ( .DIN(n5358), .Q(n2010) );
  i1s3 U4570 ( .DIN(n5354), .Q(n2011) );
  i1s3 U4571 ( .DIN(n5350), .Q(n2012) );
  i1s3 U4572 ( .DIN(n5346), .Q(n2013) );
  i1s3 U4573 ( .DIN(n5342), .Q(n2014) );
  i1s3 U4574 ( .DIN(n5338), .Q(n2015) );
  i1s3 U4575 ( .DIN(n5334), .Q(n2016) );
  i1s3 U4576 ( .DIN(n5476), .Q(n2017) );
  i1s3 U4577 ( .DIN(n5477), .Q(n2018) );
  i1s3 U4578 ( .DIN(n5478), .Q(n2019) );
  i1s3 U4579 ( .DIN(n5479), .Q(n2020) );
  i1s3 U4580 ( .DIN(n5480), .Q(n2021) );
  i1s3 U4581 ( .DIN(n5481), .Q(n2022) );
  i1s3 U4582 ( .DIN(n5482), .Q(n2023) );
  i1s3 U4583 ( .DIN(n5483), .Q(n2024) );
  i1s3 U4584 ( .DIN(n5484), .Q(n2025) );
  i1s3 U4585 ( .DIN(n5485), .Q(n2026) );
  i1s3 U4586 ( .DIN(n5486), .Q(n2027) );
  i1s3 U4587 ( .DIN(n5487), .Q(n2028) );
  i1s3 U4588 ( .DIN(n5488), .Q(n2029) );
  i1s3 U4589 ( .DIN(n5489), .Q(n2030) );
  i1s3 U4590 ( .DIN(n5490), .Q(n2031) );
  i1s3 U4591 ( .DIN(n5491), .Q(n2032) );
  i1s3 U4592 ( .DIN(n5492), .Q(n2033) );
  i1s3 U4593 ( .DIN(n5493), .Q(n2034) );
  i1s3 U4594 ( .DIN(n5494), .Q(n2035) );
  i1s3 U4595 ( .DIN(n5495), .Q(n2036) );
  i1s3 U4596 ( .DIN(n5496), .Q(n2037) );
  i1s3 U4597 ( .DIN(n5497), .Q(n2038) );
  i1s3 U4598 ( .DIN(n5498), .Q(n2039) );
  i1s3 U4599 ( .DIN(n5499), .Q(n2040) );
  i1s3 U4600 ( .DIN(n5500), .Q(n2041) );
  i1s3 U4601 ( .DIN(n5501), .Q(n2042) );
  i1s3 U4602 ( .DIN(n5502), .Q(n2043) );
  i1s3 U4603 ( .DIN(n5503), .Q(n2044) );
  i1s3 U4604 ( .DIN(n5504), .Q(n2045) );
  i1s3 U4605 ( .DIN(n5505), .Q(n2046) );
  i1s3 U4606 ( .DIN(n5506), .Q(n2047) );
  i1s3 U4607 ( .DIN(n5475), .Q(n2048) );
  i1s3 U4608 ( .DIN(n5650), .Q(n2049) );
  i1s3 U4609 ( .DIN(n5645), .Q(n2050) );
  i1s3 U4610 ( .DIN(n5640), .Q(n2051) );
  i1s3 U4611 ( .DIN(n5635), .Q(n2052) );
  i1s3 U4612 ( .DIN(n5630), .Q(n2053) );
  i1s3 U4613 ( .DIN(n5625), .Q(n2054) );
  i1s3 U4614 ( .DIN(n5620), .Q(n2055) );
  i1s3 U4615 ( .DIN(n5615), .Q(n2056) );
  i1s3 U4616 ( .DIN(n5610), .Q(n2057) );
  i1s3 U4617 ( .DIN(n5605), .Q(n2058) );
  i1s3 U4618 ( .DIN(n5600), .Q(n2059) );
  i1s3 U4619 ( .DIN(n5595), .Q(n2060) );
  i1s3 U4620 ( .DIN(n5590), .Q(n2061) );
  i1s3 U4621 ( .DIN(n5585), .Q(n2062) );
  i1s3 U4622 ( .DIN(n5580), .Q(n2063) );
  i1s3 U4623 ( .DIN(n5575), .Q(n2064) );
  i1s3 U4624 ( .DIN(n5570), .Q(n2065) );
  i1s3 U4625 ( .DIN(n5566), .Q(n2066) );
  i1s3 U4626 ( .DIN(n5562), .Q(n2067) );
  i1s3 U4627 ( .DIN(n5558), .Q(n2068) );
  i1s3 U4628 ( .DIN(n5554), .Q(n2069) );
  i1s3 U4629 ( .DIN(n5550), .Q(n2070) );
  i1s3 U4630 ( .DIN(n5546), .Q(n2071) );
  i1s3 U4631 ( .DIN(n5542), .Q(n2072) );
  i1s3 U4632 ( .DIN(n5538), .Q(n2073) );
  i1s3 U4633 ( .DIN(n5534), .Q(n2074) );
  i1s3 U4634 ( .DIN(n5530), .Q(n2075) );
  i1s3 U4635 ( .DIN(n5526), .Q(n2076) );
  i1s3 U4636 ( .DIN(n5522), .Q(n2077) );
  i1s3 U4637 ( .DIN(n5518), .Q(n2078) );
  i1s3 U4638 ( .DIN(n5514), .Q(n2079) );
  i1s3 U4639 ( .DIN(n5510), .Q(n2080) );
  i1s3 U4640 ( .DIN(n5652), .Q(n2081) );
  i1s3 U4641 ( .DIN(n5653), .Q(n2082) );
  i1s3 U4642 ( .DIN(n5654), .Q(n2083) );
  i1s3 U4643 ( .DIN(n5655), .Q(n2084) );
  i1s3 U4644 ( .DIN(n5656), .Q(n2085) );
  i1s3 U4645 ( .DIN(n5657), .Q(n2086) );
  i1s3 U4646 ( .DIN(n5658), .Q(n2087) );
  i1s3 U4647 ( .DIN(n5659), .Q(n2088) );
  i1s3 U4648 ( .DIN(n5660), .Q(n2089) );
  i1s3 U4649 ( .DIN(n5661), .Q(n2090) );
  i1s3 U4650 ( .DIN(n5662), .Q(n2091) );
  i1s3 U4651 ( .DIN(n5663), .Q(n2092) );
  i1s3 U4652 ( .DIN(n5664), .Q(n2093) );
  i1s3 U4653 ( .DIN(n5665), .Q(n2094) );
  i1s3 U4654 ( .DIN(n5666), .Q(n2095) );
  i1s3 U4655 ( .DIN(n5667), .Q(n2096) );
  i1s3 U4656 ( .DIN(n5668), .Q(n2097) );
  i1s3 U4657 ( .DIN(n5669), .Q(n2098) );
  i1s3 U4658 ( .DIN(n5670), .Q(n2099) );
  i1s3 U4659 ( .DIN(n5671), .Q(n2100) );
  i1s3 U4660 ( .DIN(n5672), .Q(n2101) );
  i1s3 U4661 ( .DIN(n5673), .Q(n2102) );
  i1s3 U4662 ( .DIN(n5674), .Q(n2103) );
  i1s3 U4663 ( .DIN(n5675), .Q(n2104) );
  i1s3 U4664 ( .DIN(n5676), .Q(n2105) );
  i1s3 U4665 ( .DIN(n5677), .Q(n2106) );
  i1s3 U4666 ( .DIN(n5678), .Q(n2107) );
  i1s3 U4667 ( .DIN(n5679), .Q(n2108) );
  i1s3 U4668 ( .DIN(n5680), .Q(n2109) );
  i1s3 U4669 ( .DIN(n5681), .Q(n2110) );
  i1s3 U4670 ( .DIN(n5682), .Q(n2111) );
  i1s3 U4671 ( .DIN(n5651), .Q(n2112) );
  i1s3 U4672 ( .DIN(n5826), .Q(n2113) );
  i1s3 U4673 ( .DIN(n5821), .Q(n2114) );
  i1s3 U4674 ( .DIN(n5816), .Q(n2115) );
  i1s3 U4675 ( .DIN(n5811), .Q(n2116) );
  i1s3 U4676 ( .DIN(n5806), .Q(n2117) );
  i1s3 U4677 ( .DIN(n5801), .Q(n2118) );
  i1s3 U4678 ( .DIN(n5796), .Q(n2119) );
  i1s3 U4679 ( .DIN(n5791), .Q(n2120) );
  i1s3 U4680 ( .DIN(n5786), .Q(n2121) );
  i1s3 U4681 ( .DIN(n5781), .Q(n2122) );
  i1s3 U4682 ( .DIN(n5776), .Q(n2123) );
  i1s3 U4683 ( .DIN(n5771), .Q(n2124) );
  i1s3 U4684 ( .DIN(n5766), .Q(n2125) );
  i1s3 U4685 ( .DIN(n5761), .Q(n2126) );
  i1s3 U4686 ( .DIN(n5756), .Q(n2127) );
  i1s3 U4687 ( .DIN(n5751), .Q(n2128) );
  i1s3 U4688 ( .DIN(n5746), .Q(n2129) );
  i1s3 U4689 ( .DIN(n5742), .Q(n2130) );
  i1s3 U4690 ( .DIN(n5738), .Q(n2131) );
  i1s3 U4691 ( .DIN(n5734), .Q(n2132) );
  i1s3 U4692 ( .DIN(n5730), .Q(n2133) );
  i1s3 U4693 ( .DIN(n5726), .Q(n2134) );
  i1s3 U4694 ( .DIN(n5722), .Q(n2135) );
  i1s3 U4695 ( .DIN(n5718), .Q(n2136) );
  i1s3 U4696 ( .DIN(n5714), .Q(n2137) );
  i1s3 U4697 ( .DIN(n5710), .Q(n2138) );
  i1s3 U4698 ( .DIN(n5706), .Q(n2139) );
  i1s3 U4699 ( .DIN(n5702), .Q(n2140) );
  i1s3 U4700 ( .DIN(n5698), .Q(n2141) );
  i1s3 U4701 ( .DIN(n5694), .Q(n2142) );
  i1s3 U4702 ( .DIN(n5690), .Q(n2143) );
  i1s3 U4703 ( .DIN(n5686), .Q(n2144) );
  i1s3 U4704 ( .DIN(n5828), .Q(n2145) );
  i1s3 U4705 ( .DIN(n5829), .Q(n2146) );
  i1s3 U4706 ( .DIN(n5830), .Q(n2147) );
  i1s3 U4707 ( .DIN(n5831), .Q(n2148) );
  i1s3 U4708 ( .DIN(n5832), .Q(n2149) );
  i1s3 U4709 ( .DIN(n5833), .Q(n2150) );
  i1s3 U4710 ( .DIN(n5834), .Q(n2151) );
  i1s3 U4711 ( .DIN(n5835), .Q(n2152) );
  i1s3 U4712 ( .DIN(n5836), .Q(n2153) );
  i1s3 U4713 ( .DIN(n5837), .Q(n2154) );
  i1s3 U4714 ( .DIN(n5838), .Q(n2155) );
  i1s3 U4715 ( .DIN(n5839), .Q(n2156) );
  i1s3 U4716 ( .DIN(n5840), .Q(n2157) );
  i1s3 U4717 ( .DIN(n5841), .Q(n2158) );
  i1s3 U4718 ( .DIN(n5842), .Q(n2159) );
  i1s3 U4719 ( .DIN(n5843), .Q(n2160) );
  i1s3 U4720 ( .DIN(n5844), .Q(n2161) );
  i1s3 U4721 ( .DIN(n5845), .Q(n2162) );
  i1s3 U4722 ( .DIN(n5846), .Q(n2163) );
  i1s3 U4723 ( .DIN(n5847), .Q(n2164) );
  i1s3 U4724 ( .DIN(n5848), .Q(n2165) );
  i1s3 U4725 ( .DIN(n5849), .Q(n2166) );
  i1s3 U4726 ( .DIN(n5850), .Q(n2167) );
  i1s3 U4727 ( .DIN(n5851), .Q(n2168) );
  i1s3 U4728 ( .DIN(n5852), .Q(n2169) );
  i1s3 U4729 ( .DIN(n5853), .Q(n2170) );
  i1s3 U4730 ( .DIN(n5854), .Q(n2171) );
  i1s3 U4731 ( .DIN(n5855), .Q(n2172) );
  i1s3 U4732 ( .DIN(n5856), .Q(n2173) );
  i1s3 U4733 ( .DIN(n5857), .Q(n2174) );
  i1s3 U4734 ( .DIN(n5858), .Q(n2175) );
  i1s3 U4735 ( .DIN(n5827), .Q(n2176) );
  i1s3 U4736 ( .DIN(n6114), .Q(n2177) );
  i1s3 U4737 ( .DIN(n6105), .Q(n2178) );
  i1s3 U4738 ( .DIN(n6096), .Q(n2179) );
  i1s3 U4739 ( .DIN(n6087), .Q(n2180) );
  i1s3 U4740 ( .DIN(n6078), .Q(n2181) );
  i1s3 U4741 ( .DIN(n6069), .Q(n2182) );
  i1s3 U4742 ( .DIN(n6060), .Q(n2183) );
  i1s3 U4743 ( .DIN(n6051), .Q(n2184) );
  i1s3 U4744 ( .DIN(n6042), .Q(n2185) );
  i1s3 U4745 ( .DIN(n6033), .Q(n2186) );
  i1s3 U4746 ( .DIN(n6024), .Q(n2187) );
  i1s3 U4747 ( .DIN(n6015), .Q(n2188) );
  i1s3 U4748 ( .DIN(n6006), .Q(n2189) );
  i1s3 U4749 ( .DIN(n5997), .Q(n2190) );
  i1s3 U4750 ( .DIN(n5988), .Q(n2191) );
  i1s3 U4751 ( .DIN(n5979), .Q(n2192) );
  i1s3 U4752 ( .DIN(n5970), .Q(n2193) );
  i1s3 U4753 ( .DIN(n5963), .Q(n2194) );
  i1s3 U4754 ( .DIN(n5956), .Q(n2195) );
  i1s3 U4755 ( .DIN(n5949), .Q(n2196) );
  i1s3 U4756 ( .DIN(n5942), .Q(n2197) );
  i1s3 U4757 ( .DIN(n5935), .Q(n2198) );
  i1s3 U4758 ( .DIN(n5928), .Q(n2199) );
  i1s3 U4759 ( .DIN(n5921), .Q(n2200) );
  i1s3 U4760 ( .DIN(n5914), .Q(n2201) );
  i1s3 U4761 ( .DIN(n5907), .Q(n2202) );
  i1s3 U4762 ( .DIN(n5900), .Q(n2203) );
  i1s3 U4763 ( .DIN(n5893), .Q(n2204) );
  i1s3 U4764 ( .DIN(n5886), .Q(n2205) );
  i1s3 U4765 ( .DIN(n5879), .Q(n2206) );
  i1s3 U4766 ( .DIN(n5872), .Q(n2207) );
  i1s3 U4767 ( .DIN(n5865), .Q(n2208) );
  i1s3 U4768 ( .DIN(n6116), .Q(n2209) );
  i1s3 U4769 ( .DIN(n6117), .Q(n2210) );
  i1s3 U4770 ( .DIN(n6118), .Q(n2211) );
  i1s3 U4771 ( .DIN(n6119), .Q(n2212) );
  i1s3 U4772 ( .DIN(n6120), .Q(n2213) );
  i1s3 U4773 ( .DIN(n6121), .Q(n2214) );
  i1s3 U4774 ( .DIN(n6122), .Q(n2215) );
  i1s3 U4775 ( .DIN(n6123), .Q(n2216) );
  i1s3 U4776 ( .DIN(n6124), .Q(n2217) );
  i1s3 U4777 ( .DIN(n6125), .Q(n2218) );
  i1s3 U4778 ( .DIN(n6126), .Q(n2219) );
  i1s3 U4779 ( .DIN(n6127), .Q(n2220) );
  i1s3 U4780 ( .DIN(n6128), .Q(n2221) );
  i1s3 U4781 ( .DIN(n6129), .Q(n2222) );
  i1s3 U4782 ( .DIN(n6130), .Q(n2223) );
  i1s3 U4783 ( .DIN(n6131), .Q(n2224) );
  i1s3 U4784 ( .DIN(n6132), .Q(n2225) );
  i1s3 U4785 ( .DIN(n6133), .Q(n2226) );
  i1s3 U4786 ( .DIN(n6134), .Q(n2227) );
  i1s3 U4787 ( .DIN(n6135), .Q(n2228) );
  i1s3 U4788 ( .DIN(n6136), .Q(n2229) );
  i1s3 U4789 ( .DIN(n6137), .Q(n2230) );
  i1s3 U4790 ( .DIN(n6138), .Q(n2231) );
  i1s3 U4791 ( .DIN(n6139), .Q(n2232) );
  i1s3 U4792 ( .DIN(n6140), .Q(n2233) );
  i1s3 U4793 ( .DIN(n6141), .Q(n2234) );
  i1s3 U4794 ( .DIN(n6142), .Q(n2235) );
  i1s3 U4795 ( .DIN(n6143), .Q(n2236) );
  i1s3 U4796 ( .DIN(n6144), .Q(n2237) );
  i1s3 U4797 ( .DIN(n6145), .Q(n2238) );
  i1s3 U4798 ( .DIN(n6146), .Q(n2239) );
  i1s3 U4799 ( .DIN(n6115), .Q(n2240) );
  i1s3 U4800 ( .DIN(n6178), .Q(n2241) );
  i1s3 U4801 ( .DIN(n6147), .Q(n2242) );
  i1s3 U4802 ( .DIN(n6148), .Q(n2243) );
  i1s3 U4803 ( .DIN(n6149), .Q(n2244) );
  i1s3 U4804 ( .DIN(n6150), .Q(n2245) );
  i1s3 U4805 ( .DIN(n6151), .Q(n2246) );
  i1s3 U4806 ( .DIN(n6152), .Q(n2247) );
  i1s3 U4807 ( .DIN(n6153), .Q(n2248) );
  i1s3 U4808 ( .DIN(n6154), .Q(n2249) );
  i1s3 U4809 ( .DIN(n6155), .Q(n2250) );
  i1s3 U4810 ( .DIN(n6156), .Q(n2251) );
  i1s3 U4811 ( .DIN(n6157), .Q(n2252) );
  i1s3 U4812 ( .DIN(n6158), .Q(n2253) );
  i1s3 U4813 ( .DIN(n6159), .Q(n2254) );
  i1s3 U4814 ( .DIN(n6160), .Q(n2255) );
  i1s3 U4815 ( .DIN(n6161), .Q(n2256) );
  i1s3 U4816 ( .DIN(n6162), .Q(n2257) );
  i1s3 U4817 ( .DIN(n6163), .Q(n2258) );
  i1s3 U4818 ( .DIN(n6164), .Q(n2259) );
  i1s3 U4819 ( .DIN(n6165), .Q(n2260) );
  i1s3 U4820 ( .DIN(n6166), .Q(n2261) );
  i1s3 U4821 ( .DIN(n6167), .Q(n2262) );
  i1s3 U4822 ( .DIN(n6168), .Q(n2263) );
  i1s3 U4823 ( .DIN(n6169), .Q(n2264) );
  i1s3 U4824 ( .DIN(n6170), .Q(n2265) );
  i1s3 U4825 ( .DIN(n6171), .Q(n2266) );
  i1s3 U4826 ( .DIN(n6172), .Q(n2267) );
  i1s3 U4827 ( .DIN(n6173), .Q(n2268) );
  i1s3 U4828 ( .DIN(n6174), .Q(n2269) );
  i1s3 U4829 ( .DIN(n6175), .Q(n2270) );
  i1s3 U4830 ( .DIN(n6176), .Q(n2271) );
  i1s3 U4831 ( .DIN(n6177), .Q(n2272) );
  i1s3 U4832 ( .DIN(n6179), .Q(n2273) );
  i1s3 U4833 ( .DIN(n6180), .Q(n2274) );
  i1s3 U4834 ( .DIN(n6181), .Q(n2275) );
  i1s3 U4835 ( .DIN(n6182), .Q(n2276) );
  i1s3 U4836 ( .DIN(n6183), .Q(n2277) );
  i1s3 U4837 ( .DIN(n6184), .Q(n2278) );
  i1s3 U4838 ( .DIN(n6185), .Q(n2279) );
  i1s3 U4839 ( .DIN(n6186), .Q(n2280) );
  i1s3 U4840 ( .DIN(n6187), .Q(n2281) );
  i1s3 U4841 ( .DIN(n6188), .Q(n2282) );
  i1s3 U4842 ( .DIN(n6189), .Q(n2283) );
  i1s3 U4843 ( .DIN(n6190), .Q(n2284) );
  i1s3 U4844 ( .DIN(n6191), .Q(n2285) );
  i1s3 U4845 ( .DIN(n6192), .Q(n2286) );
  i1s3 U4846 ( .DIN(n6193), .Q(n2287) );
  i1s3 U4847 ( .DIN(n6194), .Q(n2288) );
  i1s3 U4848 ( .DIN(n6195), .Q(n2289) );
  i1s3 U4849 ( .DIN(n6196), .Q(n2290) );
  i1s3 U4850 ( .DIN(n6286), .Q(n2291) );
  i1s3 U4851 ( .DIN(n6342), .Q(n2292) );
  i1s3 U4852 ( .DIN(n6354), .Q(n2293) );
  i1s3 U4853 ( .DIN(n6376), .Q(n2294) );
  i1s3 U4854 ( .DIN(n6377), .Q(n2295) );
  i1s3 U4855 ( .DIN(n6378), .Q(n2296) );
  i1s3 U4856 ( .DIN(n6379), .Q(n2297) );
  i1s3 U4857 ( .DIN(n6380), .Q(n2298) );
  i1s3 U4858 ( .DIN(n6381), .Q(n2299) );
  i1s3 U4859 ( .DIN(n6382), .Q(n2300) );
  i1s3 U4860 ( .DIN(n6431), .Q(n2301) );
  i1s3 U4861 ( .DIN(n6432), .Q(n2302) );
  i1s3 U4862 ( .DIN(n6433), .Q(n2303) );
  i1s3 U4863 ( .DIN(n6434), .Q(n2304) );
  i1s3 U4866 ( .DIN(TM1), .Q(n2307) );
  ib1s9 U4867 ( .DIN(n6593), .Q(n6563) );
  ib1s9 U4868 ( .DIN(n6593), .Q(n6564) );
  ib1s9 U4869 ( .DIN(n6592), .Q(n6565) );
  ib1s9 U4870 ( .DIN(n6592), .Q(n6566) );
  ib1s9 U4871 ( .DIN(n6592), .Q(n6567) );
  ib1s9 U4872 ( .DIN(n6591), .Q(n6568) );
  ib1s9 U4873 ( .DIN(n6591), .Q(n6569) );
  ib1s9 U4874 ( .DIN(n6591), .Q(n6570) );
  ib1s9 U4875 ( .DIN(n6590), .Q(n6571) );
  ib1s9 U4876 ( .DIN(n6590), .Q(n6572) );
  ib1s9 U4877 ( .DIN(n6590), .Q(n6573) );
  ib1s9 U4878 ( .DIN(n6589), .Q(n6574) );
  ib1s9 U4879 ( .DIN(n6589), .Q(n6575) );
  ib1s9 U4880 ( .DIN(n6589), .Q(n6576) );
  ib1s9 U4881 ( .DIN(n6588), .Q(n6577) );
  ib1s9 U4882 ( .DIN(n6588), .Q(n6578) );
  ib1s9 U4883 ( .DIN(n6588), .Q(n6579) );
  ib1s9 U4884 ( .DIN(n6587), .Q(n6580) );
  ib1s9 U4885 ( .DIN(n6587), .Q(n6581) );
  ib1s9 U4886 ( .DIN(n6587), .Q(n6582) );
  ib1s9 U4887 ( .DIN(n6586), .Q(n6583) );
  ib1s9 U4888 ( .DIN(n6586), .Q(n6584) );
  ib1s9 U4889 ( .DIN(n6624), .Q(n6594) );
  ib1s9 U4890 ( .DIN(n6624), .Q(n6595) );
  ib1s9 U4891 ( .DIN(n6623), .Q(n6596) );
  ib1s9 U4892 ( .DIN(n6623), .Q(n6597) );
  ib1s9 U4893 ( .DIN(n6623), .Q(n6598) );
  ib1s9 U4894 ( .DIN(n6622), .Q(n6599) );
  ib1s9 U4895 ( .DIN(n6622), .Q(n6600) );
  ib1s9 U4896 ( .DIN(n6622), .Q(n6601) );
  ib1s9 U4897 ( .DIN(n6621), .Q(n6602) );
  ib1s9 U4898 ( .DIN(n6621), .Q(n6603) );
  ib1s9 U4899 ( .DIN(n6621), .Q(n6604) );
  ib1s9 U4900 ( .DIN(n6620), .Q(n6605) );
  ib1s9 U4901 ( .DIN(n6620), .Q(n6606) );
  ib1s9 U4902 ( .DIN(n6620), .Q(n6607) );
  ib1s9 U4903 ( .DIN(n6619), .Q(n6608) );
  ib1s9 U4904 ( .DIN(n6619), .Q(n6609) );
  ib1s9 U4905 ( .DIN(n6619), .Q(n6610) );
  ib1s9 U4906 ( .DIN(n6618), .Q(n6611) );
  ib1s9 U4907 ( .DIN(n6618), .Q(n6612) );
  ib1s9 U4908 ( .DIN(n6618), .Q(n6613) );
  ib1s9 U4909 ( .DIN(n6617), .Q(n6614) );
  ib1s9 U4910 ( .DIN(n6617), .Q(n6615) );
  ib1s9 U4911 ( .DIN(n6655), .Q(n6625) );
  ib1s9 U4912 ( .DIN(n6655), .Q(n6626) );
  ib1s9 U4913 ( .DIN(n6654), .Q(n6627) );
  ib1s9 U4914 ( .DIN(n6654), .Q(n6628) );
  ib1s9 U4915 ( .DIN(n6654), .Q(n6629) );
  ib1s9 U4916 ( .DIN(n6653), .Q(n6630) );
  ib1s9 U4917 ( .DIN(n6653), .Q(n6631) );
  ib1s9 U4918 ( .DIN(n6653), .Q(n6632) );
  ib1s9 U4919 ( .DIN(n6652), .Q(n6633) );
  ib1s9 U4920 ( .DIN(n6652), .Q(n6634) );
  ib1s9 U4921 ( .DIN(n6652), .Q(n6635) );
  ib1s9 U4922 ( .DIN(n6651), .Q(n6636) );
  ib1s9 U4923 ( .DIN(n6651), .Q(n6637) );
  ib1s9 U4924 ( .DIN(n6651), .Q(n6638) );
  ib1s9 U4925 ( .DIN(n6650), .Q(n6639) );
  ib1s9 U4926 ( .DIN(n6650), .Q(n6640) );
  ib1s9 U4927 ( .DIN(n6650), .Q(n6641) );
  ib1s9 U4928 ( .DIN(n6649), .Q(n6642) );
  ib1s9 U4929 ( .DIN(n6649), .Q(n6643) );
  ib1s9 U4930 ( .DIN(n6649), .Q(n6644) );
  ib1s9 U4931 ( .DIN(n6648), .Q(n6645) );
  ib1s9 U4932 ( .DIN(n6648), .Q(n6646) );
  ib1s9 U4933 ( .DIN(n6686), .Q(n6656) );
  ib1s9 U4934 ( .DIN(n6686), .Q(n6657) );
  ib1s9 U4935 ( .DIN(n6685), .Q(n6658) );
  ib1s9 U4936 ( .DIN(n6685), .Q(n6659) );
  ib1s9 U4937 ( .DIN(n6685), .Q(n6660) );
  ib1s9 U4938 ( .DIN(n6684), .Q(n6661) );
  ib1s9 U4939 ( .DIN(n6684), .Q(n6662) );
  ib1s9 U4940 ( .DIN(n6684), .Q(n6663) );
  ib1s9 U4941 ( .DIN(n6683), .Q(n6664) );
  ib1s9 U4942 ( .DIN(n6683), .Q(n6665) );
  ib1s9 U4943 ( .DIN(n6683), .Q(n6666) );
  ib1s9 U4944 ( .DIN(n6682), .Q(n6667) );
  ib1s9 U4945 ( .DIN(n6682), .Q(n6668) );
  ib1s9 U4946 ( .DIN(n6682), .Q(n6669) );
  ib1s9 U4947 ( .DIN(n6681), .Q(n6670) );
  ib1s9 U4948 ( .DIN(n6681), .Q(n6671) );
  ib1s9 U4949 ( .DIN(n6681), .Q(n6672) );
  ib1s9 U4950 ( .DIN(n6680), .Q(n6673) );
  ib1s9 U4951 ( .DIN(n6680), .Q(n6674) );
  ib1s9 U4952 ( .DIN(n6680), .Q(n6675) );
  ib1s9 U4953 ( .DIN(n6679), .Q(n6676) );
  ib1s9 U4954 ( .DIN(n6679), .Q(n6677) );
  ib1s9 U4955 ( .DIN(n6702), .Q(n6687) );
  ib1s9 U4956 ( .DIN(n6702), .Q(n6688) );
  ib1s9 U4957 ( .DIN(n6702), .Q(n6689) );
  ib1s9 U4958 ( .DIN(n6701), .Q(n6690) );
  ib1s9 U4959 ( .DIN(n6701), .Q(n6691) );
  ib1s9 U4960 ( .DIN(n6701), .Q(n6692) );
  ib1s9 U4961 ( .DIN(n6700), .Q(n6693) );
  ib1s9 U4962 ( .DIN(n6700), .Q(n6694) );
  ib1s9 U4963 ( .DIN(n6700), .Q(n6695) );
  ib1s9 U4964 ( .DIN(n6699), .Q(n6696) );
  ib1s9 U4965 ( .DIN(n6699), .Q(n6697) );
  ib1s9 U4966 ( .DIN(n6706), .Q(n6703) );
  ib1s9 U4967 ( .DIN(n6706), .Q(n6704) );
  ib1s9 U4968 ( .DIN(RESET), .Q(n6712) );
  ib1s9 U4969 ( .DIN(RESET), .Q(n6713) );
  ib1s9 U4970 ( .DIN(RESET), .Q(n6714) );
  ib1s9 U4971 ( .DIN(RESET), .Q(n6715) );
  ib1s9 U4972 ( .DIN(RESET), .Q(n6716) );
  ib1s9 U4973 ( .DIN(RESET), .Q(n6717) );
  ib1s9 U4974 ( .DIN(RESET), .Q(n6718) );
  ib1s9 U4975 ( .DIN(RESET), .Q(n6719) );
  ib1s9 U4976 ( .DIN(RESET), .Q(n6720) );
  ib1s9 U4977 ( .DIN(RESET), .Q(n6721) );
  ib1s9 U4978 ( .DIN(RESET), .Q(n6722) );
  ib1s9 U4979 ( .DIN(RESET), .Q(n6723) );
  ib1s9 U4980 ( .DIN(RESET), .Q(n6724) );
  ib1s9 U4981 ( .DIN(RESET), .Q(n6725) );
  ib1s9 U4982 ( .DIN(RESET), .Q(n6726) );
  ib1s9 U4983 ( .DIN(RESET), .Q(n6727) );
  ib1s9 U4984 ( .DIN(RESET), .Q(n6728) );
  ib1s9 U4985 ( .DIN(RESET), .Q(n6729) );
  ib1s9 U4986 ( .DIN(RESET), .Q(n6730) );
  ib1s9 U4987 ( .DIN(RESET), .Q(n6731) );
  ib1s9 U4988 ( .DIN(RESET), .Q(n6732) );
  ib1s9 U4989 ( .DIN(RESET), .Q(n6733) );
  ib1s9 U4990 ( .DIN(RESET), .Q(n6734) );
  ib1s9 U4991 ( .DIN(RESET), .Q(n6735) );
  ib1s9 U4992 ( .DIN(RESET), .Q(n6736) );
  ib1s9 U4993 ( .DIN(RESET), .Q(n6737) );
  ib1s9 U4994 ( .DIN(RESET), .Q(n6738) );
  ib1s9 U4995 ( .DIN(RESET), .Q(n6739) );
  ib1s9 U4996 ( .DIN(RESET), .Q(n6740) );
  ib1s9 U4997 ( .DIN(RESET), .Q(n6741) );
  ib1s9 U4998 ( .DIN(RESET), .Q(n6742) );
  ib1s9 U4999 ( .DIN(RESET), .Q(n6743) );
  ib1s9 U5000 ( .DIN(RESET), .Q(n6744) );
  ib1s9 U5001 ( .DIN(RESET), .Q(n6745) );
  ib1s9 U5002 ( .DIN(RESET), .Q(n6746) );
  ib1s9 U5003 ( .DIN(RESET), .Q(n6747) );
  ib1s9 U5004 ( .DIN(RESET), .Q(n6748) );
  ib1s9 U5005 ( .DIN(RESET), .Q(n6749) );
  ib1s9 U5006 ( .DIN(RESET), .Q(n6750) );
  ib1s9 U5007 ( .DIN(RESET), .Q(n6751) );
  ib1s9 U5008 ( .DIN(RESET), .Q(n6752) );
  ib1s9 U5009 ( .DIN(RESET), .Q(n6753) );
  ib1s9 U5010 ( .DIN(RESET), .Q(n6754) );
  ib1s9 U5011 ( .DIN(RESET), .Q(n6755) );
  ib1s9 U5012 ( .DIN(RESET), .Q(n6756) );
  ib1s9 U5013 ( .DIN(RESET), .Q(n6757) );
  ib1s9 U5014 ( .DIN(RESET), .Q(n6758) );
  ib1s9 U5015 ( .DIN(RESET), .Q(n6759) );
  ib1s9 U5016 ( .DIN(RESET), .Q(n6760) );
  ib1s9 U5017 ( .DIN(RESET), .Q(n6761) );
  ib1s9 U5018 ( .DIN(RESET), .Q(n6762) );
  ib1s9 U5019 ( .DIN(RESET), .Q(n6763) );
  ib1s9 U5020 ( .DIN(RESET), .Q(n6764) );
  ib1s9 U5021 ( .DIN(RESET), .Q(n6765) );
  ib1s9 U5022 ( .DIN(RESET), .Q(n6766) );
  ib1s9 U5023 ( .DIN(RESET), .Q(n6767) );
  ib1s9 U5024 ( .DIN(RESET), .Q(n6768) );
  ib1s9 U5025 ( .DIN(RESET), .Q(n6769) );
  ib1s9 U5026 ( .DIN(RESET), .Q(n6770) );
  ib1s9 U5027 ( .DIN(RESET), .Q(n6771) );
  ib1s9 U5028 ( .DIN(RESET), .Q(n6772) );
  ib1s9 U5029 ( .DIN(RESET), .Q(n6773) );
  ib1s9 U5030 ( .DIN(RESET), .Q(n6774) );
  ib1s9 U5031 ( .DIN(RESET), .Q(n6775) );
  ib1s9 U5032 ( .DIN(RESET), .Q(n6776) );
  ib1s9 U5033 ( .DIN(RESET), .Q(n6777) );
  ib1s9 U5034 ( .DIN(RESET), .Q(n6778) );
  ib1s9 U5035 ( .DIN(RESET), .Q(n6779) );
  ib1s9 U5036 ( .DIN(RESET), .Q(n6780) );
  ib1s9 U5037 ( .DIN(RESET), .Q(n6781) );
  ib1s9 U5038 ( .DIN(RESET), .Q(n6782) );
  ib1s9 U5039 ( .DIN(RESET), .Q(n6783) );
  ib1s9 U5040 ( .DIN(RESET), .Q(n6784) );
  ib1s9 U5041 ( .DIN(RESET), .Q(n6785) );
  ib1s9 U5042 ( .DIN(RESET), .Q(n6786) );
  ib1s9 U5043 ( .DIN(RESET), .Q(n6787) );
  ib1s9 U5044 ( .DIN(RESET), .Q(n6788) );
  ib1s9 U5045 ( .DIN(RESET), .Q(n6789) );
  ib1s9 U5046 ( .DIN(RESET), .Q(n6790) );
  ib1s9 U5047 ( .DIN(RESET), .Q(n6791) );
  ib1s9 U5048 ( .DIN(RESET), .Q(n6792) );
  ib1s9 U5049 ( .DIN(RESET), .Q(n6793) );
  ib1s9 U5050 ( .DIN(RESET), .Q(n6794) );
  ib1s9 U5051 ( .DIN(RESET), .Q(n6795) );
  ib1s9 U5052 ( .DIN(RESET), .Q(n6796) );
  ib1s9 U5053 ( .DIN(RESET), .Q(n6797) );
  ib1s9 U5054 ( .DIN(RESET), .Q(n6798) );
  ib1s9 U5055 ( .DIN(RESET), .Q(n6799) );
  ib1s9 U5056 ( .DIN(RESET), .Q(n6800) );
  ib1s9 U5057 ( .DIN(RESET), .Q(n6801) );
  ib1s9 U5058 ( .DIN(RESET), .Q(n6802) );
  ib1s9 U5059 ( .DIN(RESET), .Q(n6803) );
  ib1s9 U5060 ( .DIN(RESET), .Q(n6804) );
  ib1s9 U5061 ( .DIN(RESET), .Q(n6805) );
  ib1s9 U5062 ( .DIN(RESET), .Q(n6806) );
  ib1s9 U5063 ( .DIN(RESET), .Q(n6807) );
  ib1s9 U5064 ( .DIN(RESET), .Q(n6808) );
  i1s11 U5065 ( .DIN(n6586), .Q(n6585) );
  i1s11 U5066 ( .DIN(n2317), .Q(n6586) );
  i1s11 U5067 ( .DIN(n2317), .Q(n6587) );
  i1s11 U5068 ( .DIN(n2317), .Q(n6588) );
  i1s11 U5069 ( .DIN(n2317), .Q(n6589) );
  i1s11 U5070 ( .DIN(n2317), .Q(n6590) );
  i1s11 U5071 ( .DIN(n2317), .Q(n6591) );
  i1s11 U5072 ( .DIN(n2317), .Q(n6592) );
  i1s11 U5073 ( .DIN(n2317), .Q(n6593) );
  i1s11 U5074 ( .DIN(n6617), .Q(n6616) );
  i1s11 U5075 ( .DIN(n2316), .Q(n6617) );
  i1s11 U5076 ( .DIN(n2316), .Q(n6618) );
  i1s11 U5077 ( .DIN(n2316), .Q(n6619) );
  i1s11 U5078 ( .DIN(n2316), .Q(n6620) );
  i1s11 U5079 ( .DIN(n2316), .Q(n6621) );
  i1s11 U5080 ( .DIN(n2316), .Q(n6622) );
  i1s11 U5081 ( .DIN(n2316), .Q(n6623) );
  i1s11 U5082 ( .DIN(n2316), .Q(n6624) );
  i1s11 U5083 ( .DIN(n6648), .Q(n6647) );
  i1s11 U5084 ( .DIN(n2314), .Q(n6648) );
  i1s11 U5085 ( .DIN(n2314), .Q(n6649) );
  i1s11 U5086 ( .DIN(n2314), .Q(n6650) );
  i1s11 U5087 ( .DIN(n2314), .Q(n6651) );
  i1s11 U5088 ( .DIN(n2314), .Q(n6652) );
  i1s11 U5089 ( .DIN(n2314), .Q(n6653) );
  i1s11 U5090 ( .DIN(n2314), .Q(n6654) );
  i1s11 U5091 ( .DIN(n2314), .Q(n6655) );
  i1s11 U5092 ( .DIN(n6679), .Q(n6678) );
  i1s11 U5093 ( .DIN(n2312), .Q(n6679) );
  i1s11 U5094 ( .DIN(n2312), .Q(n6680) );
  i1s11 U5095 ( .DIN(n2312), .Q(n6681) );
  i1s11 U5096 ( .DIN(n2312), .Q(n6682) );
  i1s11 U5097 ( .DIN(n2312), .Q(n6683) );
  i1s11 U5098 ( .DIN(n2312), .Q(n6684) );
  i1s11 U5099 ( .DIN(n2312), .Q(n6685) );
  i1s11 U5100 ( .DIN(n2312), .Q(n6686) );
  i1s12 U5101 ( .DIN(n6699), .Q(n6698) );
  i1s12 U5102 ( .DIN(n2307), .Q(n6699) );
  i1s12 U5103 ( .DIN(n2307), .Q(n6700) );
  i1s12 U5104 ( .DIN(n2307), .Q(n6701) );
  i1s12 U5105 ( .DIN(n2307), .Q(n6702) );
  i1s12 U5106 ( .DIN(n6706), .Q(n6705) );
  i1s12 U5107 ( .DIN(TM0), .Q(n6706) );
  i1s12 U5108 ( .DIN(TM0), .Q(n6707) );
  i1s12 U5109 ( .DIN(TM0), .Q(n6708) );
  i1s12 U5110 ( .DIN(TM0), .Q(n6709) );
  i1s12 U5111 ( .DIN(TM0), .Q(n6710) );
  i1s12 U5112 ( .DIN(TM0), .Q(n6711) );
  sdffs1 \DFF_1727/Q_reg  ( .DIN(WX11670), .SDIN(CRC_OUT_1_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_31), .QN(n6337) );
  sdffs1 \DFF_1726/Q_reg  ( .DIN(WX11668), .SDIN(CRC_OUT_1_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_30), .QN(n6336) );
  sdffs1 \DFF_1725/Q_reg  ( .DIN(WX11666), .SDIN(CRC_OUT_1_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_29), .QN(n6331) );
  sdffs1 \DFF_1724/Q_reg  ( .DIN(WX11664), .SDIN(CRC_OUT_1_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_28), .QN(n6326) );
  sdffs1 \DFF_1723/Q_reg  ( .DIN(WX11662), .SDIN(CRC_OUT_1_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_27), .QN(n6321) );
  sdffs1 \DFF_1722/Q_reg  ( .DIN(WX11660), .SDIN(CRC_OUT_1_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_26), .QN(n6316) );
  sdffs1 \DFF_1721/Q_reg  ( .DIN(WX11658), .SDIN(CRC_OUT_1_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_25), .QN(n6311) );
  sdffs1 \DFF_1720/Q_reg  ( .DIN(WX11656), .SDIN(CRC_OUT_1_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_24), .QN(n6306) );
  sdffs1 \DFF_1719/Q_reg  ( .DIN(WX11654), .SDIN(CRC_OUT_1_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_23), .QN(n6301) );
  sdffs1 \DFF_1718/Q_reg  ( .DIN(WX11652), .SDIN(CRC_OUT_1_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_22), .QN(n6296) );
  sdffs1 \DFF_1717/Q_reg  ( .DIN(WX11650), .SDIN(CRC_OUT_1_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_21), .QN(n6291) );
  sdffs1 \DFF_1716/Q_reg  ( .DIN(WX11648), .SDIN(CRC_OUT_1_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_20), .QN(n6285) );
  sdffs1 \DFF_1715/Q_reg  ( .DIN(WX11646), .SDIN(CRC_OUT_1_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_19), .QN(n6280) );
  sdffs1 \DFF_1714/Q_reg  ( .DIN(WX11644), .SDIN(CRC_OUT_1_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_18), .QN(n6275) );
  sdffs1 \DFF_1713/Q_reg  ( .DIN(WX11642), .SDIN(CRC_OUT_1_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_17), .QN(n6270) );
  sdffs1 \DFF_1712/Q_reg  ( .DIN(WX11640), .SDIN(CRC_OUT_1_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_16), .QN(n6265) );
  sdffs1 \DFF_1711/Q_reg  ( .DIN(WX11638), .SDIN(CRC_OUT_1_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_15), .QN(n6260) );
  sdffs1 \DFF_1710/Q_reg  ( .DIN(WX11636), .SDIN(CRC_OUT_1_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_14), .QN(n6256) );
  sdffs1 \DFF_1709/Q_reg  ( .DIN(WX11634), .SDIN(CRC_OUT_1_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_13), .QN(n6252) );
  sdffs1 \DFF_1708/Q_reg  ( .DIN(WX11632), .SDIN(CRC_OUT_1_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_12), .QN(n6248) );
  sdffs1 \DFF_1707/Q_reg  ( .DIN(WX11630), .SDIN(CRC_OUT_1_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_11), .QN(n6244) );
  sdffs1 \DFF_1706/Q_reg  ( .DIN(WX11628), .SDIN(CRC_OUT_1_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_10), .QN(n6240) );
  sdffs1 \DFF_1705/Q_reg  ( .DIN(WX11626), .SDIN(CRC_OUT_1_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_9), .QN(n6236) );
  sdffs1 \DFF_1704/Q_reg  ( .DIN(WX11624), .SDIN(CRC_OUT_1_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_8), .QN(n6232) );
  sdffs1 \DFF_1703/Q_reg  ( .DIN(WX11622), .SDIN(CRC_OUT_1_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_7), .QN(n6228) );
  sdffs1 \DFF_1702/Q_reg  ( .DIN(WX11620), .SDIN(CRC_OUT_1_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_6), .QN(n6224) );
  sdffs1 \DFF_1701/Q_reg  ( .DIN(WX11618), .SDIN(CRC_OUT_1_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_5), .QN(n6220) );
  sdffs1 \DFF_1700/Q_reg  ( .DIN(WX11616), .SDIN(CRC_OUT_1_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_4), .QN(n6216) );
  sdffs1 \DFF_1699/Q_reg  ( .DIN(WX11614), .SDIN(CRC_OUT_1_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_3), .QN(n6212) );
  sdffs1 \DFF_1698/Q_reg  ( .DIN(WX11612), .SDIN(CRC_OUT_1_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_2), .QN(n6208) );
  sdffs1 \DFF_1697/Q_reg  ( .DIN(WX11610), .SDIN(CRC_OUT_1_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_1_1), .QN(n6204) );
  sdffs1 \DFF_1696/Q_reg  ( .DIN(WX11608), .SDIN(n7994), .SSEL(test_se), .CLK(
        CK), .Q(CRC_OUT_1_0), .QN(n6200) );
  sdffs1 \DFF_1695/Q_reg  ( .DIN(WX11242), .SDIN(n7993), .SSEL(test_se), .CLK(
        CK), .Q(n7994), .QN(n3317) );
  sdffs1 \DFF_1694/Q_reg  ( .DIN(WX11240), .SDIN(n7992), .SSEL(test_se), .CLK(
        CK), .Q(n7993), .QN(n3318) );
  sdffs1 \DFF_1693/Q_reg  ( .DIN(WX11238), .SDIN(n7991), .SSEL(test_se), .CLK(
        CK), .Q(n7992), .QN(n3319) );
  sdffs1 \DFF_1692/Q_reg  ( .DIN(WX11236), .SDIN(n7990), .SSEL(test_se), .CLK(
        CK), .Q(n7991), .QN(n3320) );
  sdffs1 \DFF_1691/Q_reg  ( .DIN(WX11234), .SDIN(n7989), .SSEL(test_se), .CLK(
        CK), .Q(n7990), .QN(n3321) );
  sdffs1 \DFF_1690/Q_reg  ( .DIN(WX11232), .SDIN(n7988), .SSEL(test_se), .CLK(
        CK), .Q(n7989), .QN(n3322) );
  sdffs1 \DFF_1689/Q_reg  ( .DIN(WX11230), .SDIN(n7987), .SSEL(test_se), .CLK(
        CK), .Q(n7988), .QN(n3323) );
  sdffs1 \DFF_1688/Q_reg  ( .DIN(WX11228), .SDIN(n7986), .SSEL(test_se), .CLK(
        CK), .Q(n7987), .QN(n3324) );
  sdffs1 \DFF_1687/Q_reg  ( .DIN(WX11226), .SDIN(n7985), .SSEL(test_se), .CLK(
        CK), .Q(n7986), .QN(n3325) );
  sdffs1 \DFF_1686/Q_reg  ( .DIN(WX11224), .SDIN(n7984), .SSEL(test_se), .CLK(
        CK), .Q(n7985), .QN(n3326) );
  sdffs1 \DFF_1685/Q_reg  ( .DIN(WX11222), .SDIN(n7983), .SSEL(test_se), .CLK(
        CK), .Q(n7984), .QN(n3327) );
  sdffs1 \DFF_1684/Q_reg  ( .DIN(WX11220), .SDIN(n7982), .SSEL(test_se), .CLK(
        CK), .Q(n7983), .QN(n3328) );
  sdffs1 \DFF_1683/Q_reg  ( .DIN(WX11218), .SDIN(n7981), .SSEL(test_se), .CLK(
        CK), .Q(n7982), .QN(n3329) );
  sdffs1 \DFF_1682/Q_reg  ( .DIN(WX11216), .SDIN(n7980), .SSEL(test_se), .CLK(
        CK), .Q(n7981), .QN(n3330) );
  sdffs1 \DFF_1681/Q_reg  ( .DIN(WX11214), .SDIN(n7979), .SSEL(test_se), .CLK(
        CK), .Q(n7980), .QN(n3331) );
  sdffs1 \DFF_1680/Q_reg  ( .DIN(WX11212), .SDIN(n7978), .SSEL(test_se), .CLK(
        CK), .Q(n7979), .QN(n3332) );
  sdffs1 \DFF_1679/Q_reg  ( .DIN(WX11210), .SDIN(n7977), .SSEL(test_se), .CLK(
        CK), .Q(n7978), .QN(n6264) );
  sdffs1 \DFF_1678/Q_reg  ( .DIN(WX11208), .SDIN(n7976), .SSEL(test_se), .CLK(
        CK), .Q(n7977), .QN(n6269) );
  sdffs1 \DFF_1677/Q_reg  ( .DIN(WX11206), .SDIN(n7975), .SSEL(test_se), .CLK(
        CK), .Q(n7976), .QN(n6274) );
  sdffs1 \DFF_1676/Q_reg  ( .DIN(WX11204), .SDIN(n7974), .SSEL(test_se), .CLK(
        CK), .Q(n7975), .QN(n6279) );
  sdffs1 \DFF_1675/Q_reg  ( .DIN(WX11202), .SDIN(n7973), .SSEL(test_se), .CLK(
        CK), .Q(n7974), .QN(n6284) );
  sdffs1 \DFF_1674/Q_reg  ( .DIN(WX11200), .SDIN(n7972), .SSEL(test_se), .CLK(
        CK), .Q(n7973), .QN(n6290) );
  sdffs1 \DFF_1673/Q_reg  ( .DIN(WX11198), .SDIN(n7971), .SSEL(test_se), .CLK(
        CK), .Q(n7972), .QN(n6295) );
  sdffs1 \DFF_1672/Q_reg  ( .DIN(WX11196), .SDIN(n7970), .SSEL(test_se), .CLK(
        CK), .Q(n7971), .QN(n6300) );
  sdffs1 \DFF_1671/Q_reg  ( .DIN(WX11194), .SDIN(n7969), .SSEL(test_se), .CLK(
        CK), .Q(n7970), .QN(n6305) );
  sdffs1 \DFF_1670/Q_reg  ( .DIN(WX11192), .SDIN(n7968), .SSEL(test_se), .CLK(
        CK), .Q(n7969), .QN(n6310) );
  sdffs1 \DFF_1669/Q_reg  ( .DIN(WX11190), .SDIN(n7967), .SSEL(test_se), .CLK(
        CK), .Q(n7968), .QN(n6315) );
  sdffs1 \DFF_1668/Q_reg  ( .DIN(WX11188), .SDIN(n7966), .SSEL(test_se), .CLK(
        CK), .Q(n7967), .QN(n6320) );
  sdffs1 \DFF_1667/Q_reg  ( .DIN(WX11186), .SDIN(n7965), .SSEL(test_se), .CLK(
        CK), .Q(n7966), .QN(n6325) );
  sdffs1 \DFF_1666/Q_reg  ( .DIN(WX11184), .SDIN(n7964), .SSEL(test_se), .CLK(
        CK), .Q(n7965), .QN(n6330) );
  sdffs1 \DFF_1665/Q_reg  ( .DIN(WX11182), .SDIN(n7963), .SSEL(test_se), .CLK(
        CK), .Q(n7964), .QN(n6335) );
  sdffs1 \DFF_1664/Q_reg  ( .DIN(WX11180), .SDIN(n7962), .SSEL(test_se), .CLK(
        CK), .Q(n7963), .QN(n6341) );
  sdffs1 \DFF_1663/Q_reg  ( .DIN(WX11178), .SDIN(n7961), .SSEL(test_se), .CLK(
        CK), .Q(n7962), .QN(n6199) );
  sdffs1 \DFF_1662/Q_reg  ( .DIN(WX11176), .SDIN(n7960), .SSEL(test_se), .CLK(
        CK), .Q(n7961), .QN(n6203) );
  sdffs1 \DFF_1661/Q_reg  ( .DIN(WX11174), .SDIN(n7959), .SSEL(test_se), .CLK(
        CK), .Q(n7960), .QN(n6207) );
  sdffs1 \DFF_1660/Q_reg  ( .DIN(WX11172), .SDIN(n7958), .SSEL(test_se), .CLK(
        CK), .Q(n7959), .QN(n6211) );
  sdffs1 \DFF_1659/Q_reg  ( .DIN(WX11170), .SDIN(n7957), .SSEL(test_se), .CLK(
        CK), .Q(n7958), .QN(n6215) );
  sdffs1 \DFF_1658/Q_reg  ( .DIN(WX11168), .SDIN(n7956), .SSEL(test_se), .CLK(
        CK), .Q(n7957), .QN(n6219) );
  sdffs1 \DFF_1657/Q_reg  ( .DIN(WX11166), .SDIN(n7955), .SSEL(test_se), .CLK(
        CK), .Q(n7956), .QN(n6223) );
  sdffs1 \DFF_1656/Q_reg  ( .DIN(WX11164), .SDIN(n7954), .SSEL(test_se), .CLK(
        CK), .Q(n7955), .QN(n6227) );
  sdffs1 \DFF_1655/Q_reg  ( .DIN(WX11162), .SDIN(n7953), .SSEL(test_se), .CLK(
        CK), .Q(n7954), .QN(n6231) );
  sdffs1 \DFF_1654/Q_reg  ( .DIN(WX11160), .SDIN(n7952), .SSEL(test_se), .CLK(
        CK), .Q(n7953), .QN(n6235) );
  sdffs1 \DFF_1653/Q_reg  ( .DIN(WX11158), .SDIN(n7951), .SSEL(test_se), .CLK(
        CK), .Q(n7952), .QN(n6239) );
  sdffs1 \DFF_1652/Q_reg  ( .DIN(WX11156), .SDIN(n7950), .SSEL(test_se), .CLK(
        CK), .Q(n7951), .QN(n6243) );
  sdffs1 \DFF_1651/Q_reg  ( .DIN(WX11154), .SDIN(n7949), .SSEL(test_se), .CLK(
        CK), .Q(n7950), .QN(n6247) );
  sdffs1 \DFF_1650/Q_reg  ( .DIN(WX11152), .SDIN(n7948), .SSEL(test_se), .CLK(
        CK), .Q(n7949), .QN(n6251) );
  sdffs1 \DFF_1649/Q_reg  ( .DIN(WX11150), .SDIN(n7947), .SSEL(test_se), .CLK(
        CK), .Q(n7948), .QN(n6255) );
  sdffs1 \DFF_1648/Q_reg  ( .DIN(WX11148), .SDIN(n7946), .SSEL(test_se), .CLK(
        CK), .Q(n7947), .QN(n6259) );
  sdffs1 \DFF_1647/Q_reg  ( .DIN(WX11146), .SDIN(n7945), .SSEL(test_se), .CLK(
        CK), .Q(n7946), .QN(n6263) );
  sdffs1 \DFF_1646/Q_reg  ( .DIN(WX11144), .SDIN(n7944), .SSEL(test_se), .CLK(
        CK), .Q(n7945), .QN(n6268) );
  sdffs1 \DFF_1645/Q_reg  ( .DIN(WX11142), .SDIN(n7943), .SSEL(test_se), .CLK(
        CK), .Q(n7944), .QN(n6273) );
  sdffs1 \DFF_1644/Q_reg  ( .DIN(WX11140), .SDIN(n7942), .SSEL(test_se), .CLK(
        CK), .Q(n7943), .QN(n6278) );
  sdffs1 \DFF_1643/Q_reg  ( .DIN(WX11138), .SDIN(n7941), .SSEL(test_se), .CLK(
        CK), .Q(n7942), .QN(n6283) );
  sdffs1 \DFF_1642/Q_reg  ( .DIN(WX11136), .SDIN(n7940), .SSEL(test_se), .CLK(
        CK), .Q(n7941), .QN(n6289) );
  sdffs1 \DFF_1641/Q_reg  ( .DIN(WX11134), .SDIN(n7939), .SSEL(test_se), .CLK(
        CK), .Q(n7940), .QN(n6294) );
  sdffs1 \DFF_1640/Q_reg  ( .DIN(WX11132), .SDIN(n7938), .SSEL(test_se), .CLK(
        CK), .Q(n7939), .QN(n6299) );
  sdffs1 \DFF_1639/Q_reg  ( .DIN(WX11130), .SDIN(n7937), .SSEL(test_se), .CLK(
        CK), .Q(n7938), .QN(n6304) );
  sdffs1 \DFF_1638/Q_reg  ( .DIN(WX11128), .SDIN(n7936), .SSEL(test_se), .CLK(
        CK), .Q(n7937), .QN(n6309) );
  sdffs1 \DFF_1637/Q_reg  ( .DIN(WX11126), .SDIN(n7935), .SSEL(test_se), .CLK(
        CK), .Q(n7936), .QN(n6314) );
  sdffs1 \DFF_1636/Q_reg  ( .DIN(WX11124), .SDIN(n7934), .SSEL(test_se), .CLK(
        CK), .Q(n7935), .QN(n6319) );
  sdffs1 \DFF_1635/Q_reg  ( .DIN(WX11122), .SDIN(n7933), .SSEL(test_se), .CLK(
        CK), .Q(n7934), .QN(n6324) );
  sdffs1 \DFF_1634/Q_reg  ( .DIN(WX11120), .SDIN(n7932), .SSEL(test_se), .CLK(
        CK), .Q(n7933), .QN(n6329) );
  sdffs1 \DFF_1633/Q_reg  ( .DIN(WX11118), .SDIN(n7931), .SSEL(test_se), .CLK(
        CK), .Q(n7932), .QN(n6334) );
  sdffs1 \DFF_1632/Q_reg  ( .DIN(WX11116), .SDIN(n6198), .SSEL(test_se), .CLK(
        CK), .Q(n7931), .QN(n6340) );
  sdffs1 \DFF_1631/Q_reg  ( .DIN(WX11114), .SDIN(n6202), .SSEL(test_se), .CLK(
        CK), .Q(n6198) );
  sdffs1 \DFF_1630/Q_reg  ( .DIN(WX11112), .SDIN(n6206), .SSEL(test_se), .CLK(
        CK), .Q(n6202) );
  sdffs1 \DFF_1629/Q_reg  ( .DIN(WX11110), .SDIN(n6210), .SSEL(test_se), .CLK(
        CK), .Q(n6206) );
  sdffs1 \DFF_1628/Q_reg  ( .DIN(WX11108), .SDIN(n6214), .SSEL(test_se), .CLK(
        CK), .Q(n6210) );
  sdffs1 \DFF_1627/Q_reg  ( .DIN(WX11106), .SDIN(n6218), .SSEL(test_se), .CLK(
        CK), .Q(n6214) );
  sdffs1 \DFF_1626/Q_reg  ( .DIN(WX11104), .SDIN(n6222), .SSEL(test_se), .CLK(
        CK), .Q(n6218) );
  sdffs1 \DFF_1625/Q_reg  ( .DIN(WX11102), .SDIN(n6226), .SSEL(test_se), .CLK(
        CK), .Q(n6222) );
  sdffs1 \DFF_1624/Q_reg  ( .DIN(WX11100), .SDIN(n6230), .SSEL(test_se), .CLK(
        CK), .Q(n6226) );
  sdffs1 \DFF_1623/Q_reg  ( .DIN(WX11098), .SDIN(n6234), .SSEL(test_se), .CLK(
        CK), .Q(n6230) );
  sdffs1 \DFF_1622/Q_reg  ( .DIN(WX11096), .SDIN(n6238), .SSEL(test_se), .CLK(
        CK), .Q(n6234) );
  sdffs1 \DFF_1621/Q_reg  ( .DIN(WX11094), .SDIN(n6242), .SSEL(test_se), .CLK(
        CK), .Q(n6238) );
  sdffs1 \DFF_1620/Q_reg  ( .DIN(WX11092), .SDIN(n6246), .SSEL(test_se), .CLK(
        CK), .Q(n6242) );
  sdffs1 \DFF_1619/Q_reg  ( .DIN(WX11090), .SDIN(n6250), .SSEL(test_se), .CLK(
        CK), .Q(n6246) );
  sdffs1 \DFF_1618/Q_reg  ( .DIN(WX11088), .SDIN(n6254), .SSEL(test_se), .CLK(
        CK), .Q(n6250) );
  sdffs1 \DFF_1617/Q_reg  ( .DIN(WX11086), .SDIN(n6258), .SSEL(test_se), .CLK(
        CK), .Q(n6254) );
  sdffs1 \DFF_1616/Q_reg  ( .DIN(WX11084), .SDIN(n6262), .SSEL(test_se), .CLK(
        CK), .Q(n6258) );
  sdffs1 \DFF_1615/Q_reg  ( .DIN(WX11082), .SDIN(n6267), .SSEL(test_se), .CLK(
        CK), .Q(n6262) );
  sdffs1 \DFF_1614/Q_reg  ( .DIN(WX11080), .SDIN(n6272), .SSEL(test_se), .CLK(
        CK), .Q(n6267) );
  sdffs1 \DFF_1613/Q_reg  ( .DIN(WX11078), .SDIN(n6277), .SSEL(test_se), .CLK(
        CK), .Q(n6272) );
  sdffs1 \DFF_1612/Q_reg  ( .DIN(WX11076), .SDIN(n6282), .SSEL(test_se), .CLK(
        CK), .Q(n6277) );
  sdffs1 \DFF_1611/Q_reg  ( .DIN(WX11074), .SDIN(n6288), .SSEL(test_se), .CLK(
        CK), .Q(n6282) );
  sdffs1 \DFF_1610/Q_reg  ( .DIN(WX11072), .SDIN(n6293), .SSEL(test_se), .CLK(
        CK), .Q(n6288) );
  sdffs1 \DFF_1609/Q_reg  ( .DIN(WX11070), .SDIN(n6298), .SSEL(test_se), .CLK(
        CK), .Q(n6293) );
  sdffs1 \DFF_1608/Q_reg  ( .DIN(WX11068), .SDIN(n6303), .SSEL(test_se), .CLK(
        CK), .Q(n6298) );
  sdffs1 \DFF_1607/Q_reg  ( .DIN(WX11066), .SDIN(n6308), .SSEL(test_se), .CLK(
        CK), .Q(n6303) );
  sdffs1 \DFF_1606/Q_reg  ( .DIN(WX11064), .SDIN(n6313), .SSEL(test_se), .CLK(
        CK), .Q(n6308) );
  sdffs1 \DFF_1605/Q_reg  ( .DIN(WX11062), .SDIN(n6318), .SSEL(test_se), .CLK(
        CK), .Q(n6313) );
  sdffs1 \DFF_1604/Q_reg  ( .DIN(WX11060), .SDIN(n6323), .SSEL(test_se), .CLK(
        CK), .Q(n6318) );
  sdffs1 \DFF_1603/Q_reg  ( .DIN(WX11058), .SDIN(n6328), .SSEL(test_se), .CLK(
        CK), .Q(n6323) );
  sdffs1 \DFF_1602/Q_reg  ( .DIN(WX11056), .SDIN(n6333), .SSEL(test_se), .CLK(
        CK), .Q(n6328) );
  sdffs1 \DFF_1601/Q_reg  ( .DIN(WX11054), .SDIN(n6339), .SSEL(test_se), .CLK(
        CK), .Q(n6333) );
  sdffs1 \DFF_1600/Q_reg  ( .DIN(WX11052), .SDIN(n7930), .SSEL(test_se), .CLK(
        CK), .Q(n6339) );
  sdffs1 \DFF_1599/Q_reg  ( .DIN(WX11050), .SDIN(n7929), .SSEL(test_se), .CLK(
        CK), .Q(n7930), .QN(n6197) );
  sdffs1 \DFF_1598/Q_reg  ( .DIN(WX11048), .SDIN(n7928), .SSEL(test_se), .CLK(
        CK), .Q(n7929), .QN(n6201) );
  sdffs1 \DFF_1597/Q_reg  ( .DIN(WX11046), .SDIN(n7927), .SSEL(test_se), .CLK(
        CK), .Q(n7928), .QN(n6205) );
  sdffs1 \DFF_1596/Q_reg  ( .DIN(WX11044), .SDIN(n7926), .SSEL(test_se), .CLK(
        CK), .Q(n7927), .QN(n6209) );
  sdffs1 \DFF_1595/Q_reg  ( .DIN(WX11042), .SDIN(n7925), .SSEL(test_se), .CLK(
        CK), .Q(n7926), .QN(n6213) );
  sdffs1 \DFF_1594/Q_reg  ( .DIN(WX11040), .SDIN(n7924), .SSEL(test_se), .CLK(
        CK), .Q(n7925), .QN(n6217) );
  sdffs1 \DFF_1593/Q_reg  ( .DIN(WX11038), .SDIN(n7923), .SSEL(test_se), .CLK(
        CK), .Q(n7924), .QN(n6221) );
  sdffs1 \DFF_1592/Q_reg  ( .DIN(WX11036), .SDIN(n7922), .SSEL(test_se), .CLK(
        CK), .Q(n7923), .QN(n6225) );
  sdffs1 \DFF_1591/Q_reg  ( .DIN(WX11034), .SDIN(n7921), .SSEL(test_se), .CLK(
        CK), .Q(n7922), .QN(n6229) );
  sdffs1 \DFF_1590/Q_reg  ( .DIN(WX11032), .SDIN(n7920), .SSEL(test_se), .CLK(
        CK), .Q(n7921), .QN(n6233) );
  sdffs1 \DFF_1589/Q_reg  ( .DIN(WX11030), .SDIN(n7919), .SSEL(test_se), .CLK(
        CK), .Q(n7920), .QN(n6237) );
  sdffs1 \DFF_1588/Q_reg  ( .DIN(WX11028), .SDIN(n7918), .SSEL(test_se), .CLK(
        CK), .Q(n7919), .QN(n6241) );
  sdffs1 \DFF_1587/Q_reg  ( .DIN(WX11026), .SDIN(n7917), .SSEL(test_se), .CLK(
        CK), .Q(n7918), .QN(n6245) );
  sdffs1 \DFF_1586/Q_reg  ( .DIN(WX11024), .SDIN(n7916), .SSEL(test_se), .CLK(
        CK), .Q(n7917), .QN(n6249) );
  sdffs1 \DFF_1585/Q_reg  ( .DIN(WX11022), .SDIN(n7915), .SSEL(test_se), .CLK(
        CK), .Q(n7916), .QN(n6253) );
  sdffs1 \DFF_1584/Q_reg  ( .DIN(WX11020), .SDIN(n7914), .SSEL(test_se), .CLK(
        CK), .Q(n7915), .QN(n6257) );
  sdffs1 \DFF_1583/Q_reg  ( .DIN(WX11018), .SDIN(n7913), .SSEL(test_se), .CLK(
        CK), .Q(n7914), .QN(n6261) );
  sdffs1 \DFF_1582/Q_reg  ( .DIN(WX11016), .SDIN(n7912), .SSEL(test_se), .CLK(
        CK), .Q(n7913), .QN(n6266) );
  sdffs1 \DFF_1581/Q_reg  ( .DIN(WX11014), .SDIN(n7911), .SSEL(test_se), .CLK(
        CK), .Q(n7912), .QN(n6271) );
  sdffs1 \DFF_1580/Q_reg  ( .DIN(WX11012), .SDIN(n7910), .SSEL(test_se), .CLK(
        CK), .Q(n7911), .QN(n6276) );
  sdffs1 \DFF_1579/Q_reg  ( .DIN(WX11010), .SDIN(n7909), .SSEL(test_se), .CLK(
        CK), .Q(n7910), .QN(n6281) );
  sdffs1 \DFF_1578/Q_reg  ( .DIN(WX11008), .SDIN(n7908), .SSEL(test_se), .CLK(
        CK), .Q(n7909), .QN(n6287) );
  sdffs1 \DFF_1577/Q_reg  ( .DIN(WX11006), .SDIN(n7907), .SSEL(test_se), .CLK(
        CK), .Q(n7908), .QN(n6292) );
  sdffs1 \DFF_1576/Q_reg  ( .DIN(WX11004), .SDIN(n7906), .SSEL(test_se), .CLK(
        CK), .Q(n7907), .QN(n6297) );
  sdffs1 \DFF_1575/Q_reg  ( .DIN(WX11002), .SDIN(n7905), .SSEL(test_se), .CLK(
        CK), .Q(n7906), .QN(n6302) );
  sdffs1 \DFF_1574/Q_reg  ( .DIN(WX11000), .SDIN(n7904), .SSEL(test_se), .CLK(
        CK), .Q(n7905), .QN(n6307) );
  sdffs1 \DFF_1573/Q_reg  ( .DIN(WX10998), .SDIN(n7903), .SSEL(test_se), .CLK(
        CK), .Q(n7904), .QN(n6312) );
  sdffs1 \DFF_1572/Q_reg  ( .DIN(WX10996), .SDIN(n7902), .SSEL(test_se), .CLK(
        CK), .Q(n7903), .QN(n6317) );
  sdffs1 \DFF_1571/Q_reg  ( .DIN(WX10994), .SDIN(n7901), .SSEL(test_se), .CLK(
        CK), .Q(n7902), .QN(n6322) );
  sdffs1 \DFF_1570/Q_reg  ( .DIN(WX10992), .SDIN(n7900), .SSEL(test_se), .CLK(
        CK), .Q(n7901), .QN(n6327) );
  sdffs1 \DFF_1569/Q_reg  ( .DIN(WX10990), .SDIN(n7899), .SSEL(test_se), .CLK(
        CK), .Q(n7900), .QN(n6332) );
  sdffs1 \DFF_1568/Q_reg  ( .DIN(WX10988), .SDIN(n7898), .SSEL(test_se), .CLK(
        CK), .Q(n7899), .QN(n6338) );
  sdffs1 \DFF_1567/Q_reg  ( .DIN(WX10890), .SDIN(n7897), .SSEL(test_se), .CLK(
        CK), .Q(n7898), .QN(n6344) );
  sdffs1 \DFF_1566/Q_reg  ( .DIN(WX10888), .SDIN(n7896), .SSEL(test_se), .CLK(
        CK), .Q(n7897), .QN(n6345) );
  sdffs1 \DFF_1565/Q_reg  ( .DIN(WX10886), .SDIN(n7895), .SSEL(test_se), .CLK(
        CK), .Q(n7896), .QN(n6346) );
  sdffs1 \DFF_1564/Q_reg  ( .DIN(WX10884), .SDIN(n7894), .SSEL(test_se), .CLK(
        CK), .Q(n7895), .QN(n6347) );
  sdffs1 \DFF_1563/Q_reg  ( .DIN(WX10882), .SDIN(n7893), .SSEL(test_se), .CLK(
        CK), .Q(n7894), .QN(n6348) );
  sdffs1 \DFF_1562/Q_reg  ( .DIN(WX10880), .SDIN(n7892), .SSEL(test_se), .CLK(
        CK), .Q(n7893), .QN(n6349) );
  sdffs1 \DFF_1561/Q_reg  ( .DIN(WX10878), .SDIN(n7891), .SSEL(test_se), .CLK(
        CK), .Q(n7892), .QN(n6350) );
  sdffs1 \DFF_1560/Q_reg  ( .DIN(WX10876), .SDIN(n7890), .SSEL(test_se), .CLK(
        CK), .Q(n7891), .QN(n6351) );
  sdffs1 \DFF_1559/Q_reg  ( .DIN(WX10874), .SDIN(n7889), .SSEL(test_se), .CLK(
        CK), .Q(n7890), .QN(n6352) );
  sdffs1 \DFF_1558/Q_reg  ( .DIN(WX10872), .SDIN(n7888), .SSEL(test_se), .CLK(
        CK), .Q(n7889), .QN(n6353) );
  sdffs1 \DFF_1557/Q_reg  ( .DIN(WX10870), .SDIN(n7887), .SSEL(test_se), .CLK(
        CK), .Q(n7888), .QN(n6355) );
  sdffs1 \DFF_1556/Q_reg  ( .DIN(WX10868), .SDIN(n7886), .SSEL(test_se), .CLK(
        CK), .Q(n7887), .QN(n6356) );
  sdffs1 \DFF_1555/Q_reg  ( .DIN(WX10866), .SDIN(n7885), .SSEL(test_se), .CLK(
        CK), .Q(n7886), .QN(n6357) );
  sdffs1 \DFF_1554/Q_reg  ( .DIN(WX10864), .SDIN(n7884), .SSEL(test_se), .CLK(
        CK), .Q(n7885), .QN(n6358) );
  sdffs1 \DFF_1553/Q_reg  ( .DIN(WX10862), .SDIN(n7883), .SSEL(test_se), .CLK(
        CK), .Q(n7884), .QN(n6359) );
  sdffs1 \DFF_1552/Q_reg  ( .DIN(WX10860), .SDIN(n7882), .SSEL(test_se), .CLK(
        CK), .Q(n7883), .QN(n6360) );
  sdffs1 \DFF_1551/Q_reg  ( .DIN(WX10858), .SDIN(n7881), .SSEL(test_se), .CLK(
        CK), .Q(n7882), .QN(n6361) );
  sdffs1 \DFF_1550/Q_reg  ( .DIN(WX10856), .SDIN(n7880), .SSEL(test_se), .CLK(
        CK), .Q(n7881), .QN(n6362) );
  sdffs1 \DFF_1549/Q_reg  ( .DIN(WX10854), .SDIN(n7879), .SSEL(test_se), .CLK(
        CK), .Q(n7880), .QN(n6363) );
  sdffs1 \DFF_1548/Q_reg  ( .DIN(WX10852), .SDIN(n7878), .SSEL(test_se), .CLK(
        CK), .Q(n7879), .QN(n6364) );
  sdffs1 \DFF_1547/Q_reg  ( .DIN(WX10850), .SDIN(n7877), .SSEL(test_se), .CLK(
        CK), .Q(n7878), .QN(n6365) );
  sdffs1 \DFF_1546/Q_reg  ( .DIN(WX10848), .SDIN(n7876), .SSEL(test_se), .CLK(
        CK), .Q(n7877), .QN(n6366) );
  sdffs1 \DFF_1545/Q_reg  ( .DIN(WX10846), .SDIN(n7875), .SSEL(test_se), .CLK(
        CK), .Q(n7876), .QN(n6367) );
  sdffs1 \DFF_1544/Q_reg  ( .DIN(WX10844), .SDIN(n7874), .SSEL(test_se), .CLK(
        CK), .Q(n7875), .QN(n6368) );
  sdffs1 \DFF_1543/Q_reg  ( .DIN(WX10842), .SDIN(n7873), .SSEL(test_se), .CLK(
        CK), .Q(n7874), .QN(n6369) );
  sdffs1 \DFF_1542/Q_reg  ( .DIN(WX10840), .SDIN(n7872), .SSEL(test_se), .CLK(
        CK), .Q(n7873), .QN(n6370) );
  sdffs1 \DFF_1541/Q_reg  ( .DIN(WX10838), .SDIN(n7871), .SSEL(test_se), .CLK(
        CK), .Q(n7872), .QN(n6371) );
  sdffs1 \DFF_1540/Q_reg  ( .DIN(WX10836), .SDIN(n7870), .SSEL(test_se), .CLK(
        CK), .Q(n7871), .QN(n6372) );
  sdffs1 \DFF_1539/Q_reg  ( .DIN(WX10834), .SDIN(n7869), .SSEL(test_se), .CLK(
        CK), .Q(n7870), .QN(n6373) );
  sdffs1 \DFF_1538/Q_reg  ( .DIN(WX10832), .SDIN(n7868), .SSEL(test_se), .CLK(
        CK), .Q(n7869), .QN(n6374) );
  sdffs1 \DFF_1537/Q_reg  ( .DIN(WX10830), .SDIN(n7867), .SSEL(test_se), .CLK(
        CK), .Q(n7868), .QN(n6375) );
  sdffs1 \DFF_1536/Q_reg  ( .DIN(WX10828), .SDIN(CRC_OUT_2_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7867), .QN(n6343) );
  sdffs1 \DFF_1535/Q_reg  ( .DIN(WX10377), .SDIN(CRC_OUT_2_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_31), .QN(n6430) );
  sdffs1 \DFF_1534/Q_reg  ( .DIN(WX10375), .SDIN(CRC_OUT_2_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_30), .QN(n6383) );
  sdffs1 \DFF_1533/Q_reg  ( .DIN(WX10373), .SDIN(CRC_OUT_2_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_29), .QN(n6385) );
  sdffs1 \DFF_1532/Q_reg  ( .DIN(WX10371), .SDIN(CRC_OUT_2_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_28), .QN(n6387) );
  sdffs1 \DFF_1531/Q_reg  ( .DIN(WX10369), .SDIN(CRC_OUT_2_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_27), .QN(n6389) );
  sdffs1 \DFF_1530/Q_reg  ( .DIN(WX10367), .SDIN(CRC_OUT_2_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_26), .QN(n6391) );
  sdffs1 \DFF_1529/Q_reg  ( .DIN(WX10365), .SDIN(CRC_OUT_2_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_25), .QN(n6393) );
  sdffs1 \DFF_1528/Q_reg  ( .DIN(WX10363), .SDIN(CRC_OUT_2_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_24), .QN(n6395) );
  sdffs1 \DFF_1527/Q_reg  ( .DIN(WX10361), .SDIN(CRC_OUT_2_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_23), .QN(n6397) );
  sdffs1 \DFF_1526/Q_reg  ( .DIN(WX10359), .SDIN(CRC_OUT_2_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_22), .QN(n6399) );
  sdffs1 \DFF_1525/Q_reg  ( .DIN(WX10357), .SDIN(CRC_OUT_2_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_21), .QN(n6401) );
  sdffs1 \DFF_1524/Q_reg  ( .DIN(WX10355), .SDIN(CRC_OUT_2_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_20), .QN(n6403) );
  sdffs1 \DFF_1523/Q_reg  ( .DIN(WX10353), .SDIN(CRC_OUT_2_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_19), .QN(n6405) );
  sdffs1 \DFF_1522/Q_reg  ( .DIN(WX10351), .SDIN(CRC_OUT_2_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_18), .QN(n6407) );
  sdffs1 \DFF_1521/Q_reg  ( .DIN(WX10349), .SDIN(CRC_OUT_2_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_17), .QN(n6409) );
  sdffs1 \DFF_1520/Q_reg  ( .DIN(WX10347), .SDIN(CRC_OUT_2_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_16), .QN(n6411) );
  sdffs1 \DFF_1519/Q_reg  ( .DIN(WX10345), .SDIN(CRC_OUT_2_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_15), .QN(n6413) );
  sdffs1 \DFF_1518/Q_reg  ( .DIN(WX10343), .SDIN(CRC_OUT_2_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_14), .QN(n6415) );
  sdffs1 \DFF_1517/Q_reg  ( .DIN(WX10341), .SDIN(CRC_OUT_2_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_13), .QN(n6416) );
  sdffs1 \DFF_1516/Q_reg  ( .DIN(WX10339), .SDIN(CRC_OUT_2_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_12), .QN(n6417) );
  sdffs1 \DFF_1515/Q_reg  ( .DIN(WX10337), .SDIN(CRC_OUT_2_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_11), .QN(n6418) );
  sdffs1 \DFF_1514/Q_reg  ( .DIN(WX10335), .SDIN(CRC_OUT_2_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_10), .QN(n6419) );
  sdffs1 \DFF_1513/Q_reg  ( .DIN(WX10333), .SDIN(CRC_OUT_2_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_9), .QN(n6420) );
  sdffs1 \DFF_1512/Q_reg  ( .DIN(WX10331), .SDIN(CRC_OUT_2_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_8), .QN(n6421) );
  sdffs1 \DFF_1511/Q_reg  ( .DIN(WX10329), .SDIN(CRC_OUT_2_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_7), .QN(n6422) );
  sdffs1 \DFF_1510/Q_reg  ( .DIN(WX10327), .SDIN(CRC_OUT_2_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_6), .QN(n6423) );
  sdffs1 \DFF_1509/Q_reg  ( .DIN(WX10325), .SDIN(CRC_OUT_2_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_5), .QN(n6424) );
  sdffs1 \DFF_1508/Q_reg  ( .DIN(WX10323), .SDIN(CRC_OUT_2_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_4), .QN(n6425) );
  sdffs1 \DFF_1507/Q_reg  ( .DIN(WX10321), .SDIN(CRC_OUT_2_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_3), .QN(n6426) );
  sdffs1 \DFF_1506/Q_reg  ( .DIN(WX10319), .SDIN(CRC_OUT_2_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_2), .QN(n6427) );
  sdffs1 \DFF_1505/Q_reg  ( .DIN(WX10317), .SDIN(CRC_OUT_2_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_2_1), .QN(n6428) );
  sdffs1 \DFF_1504/Q_reg  ( .DIN(WX10315), .SDIN(n7866), .SSEL(test_se), .CLK(
        CK), .Q(CRC_OUT_2_0), .QN(n6429) );
  sdffs1 \DFF_1503/Q_reg  ( .DIN(WX9949), .SDIN(n7865), .SSEL(test_se), .CLK(
        CK), .Q(n7866), .QN(n3205) );
  sdffs1 \DFF_1502/Q_reg  ( .DIN(WX9947), .SDIN(n7864), .SSEL(test_se), .CLK(
        CK), .Q(n7865), .QN(n3206) );
  sdffs1 \DFF_1501/Q_reg  ( .DIN(WX9945), .SDIN(n7863), .SSEL(test_se), .CLK(
        CK), .Q(n7864), .QN(n3207) );
  sdffs1 \DFF_1500/Q_reg  ( .DIN(WX9943), .SDIN(n7862), .SSEL(test_se), .CLK(
        CK), .Q(n7863), .QN(n3208) );
  sdffs1 \DFF_1499/Q_reg  ( .DIN(WX9941), .SDIN(n7861), .SSEL(test_se), .CLK(
        CK), .Q(n7862), .QN(n3209) );
  sdffs1 \DFF_1498/Q_reg  ( .DIN(WX9939), .SDIN(n7860), .SSEL(test_se), .CLK(
        CK), .Q(n7861), .QN(n3210) );
  sdffs1 \DFF_1497/Q_reg  ( .DIN(WX9937), .SDIN(n7859), .SSEL(test_se), .CLK(
        CK), .Q(n7860), .QN(n3211) );
  sdffs1 \DFF_1496/Q_reg  ( .DIN(WX9935), .SDIN(n7858), .SSEL(test_se), .CLK(
        CK), .Q(n7859), .QN(n3212) );
  sdffs1 \DFF_1495/Q_reg  ( .DIN(WX9933), .SDIN(n7857), .SSEL(test_se), .CLK(
        CK), .Q(n7858), .QN(n3213) );
  sdffs1 \DFF_1494/Q_reg  ( .DIN(WX9931), .SDIN(n7856), .SSEL(test_se), .CLK(
        CK), .Q(n7857), .QN(n3214) );
  sdffs1 \DFF_1493/Q_reg  ( .DIN(WX9929), .SDIN(n7855), .SSEL(test_se), .CLK(
        CK), .Q(n7856), .QN(n3215) );
  sdffs1 \DFF_1492/Q_reg  ( .DIN(WX9927), .SDIN(n7854), .SSEL(test_se), .CLK(
        CK), .Q(n7855), .QN(n3216) );
  sdffs1 \DFF_1491/Q_reg  ( .DIN(WX9925), .SDIN(n7853), .SSEL(test_se), .CLK(
        CK), .Q(n7854), .QN(n3217) );
  sdffs1 \DFF_1490/Q_reg  ( .DIN(WX9923), .SDIN(n7852), .SSEL(test_se), .CLK(
        CK), .Q(n7853), .QN(n3218) );
  sdffs1 \DFF_1489/Q_reg  ( .DIN(WX9921), .SDIN(n7851), .SSEL(test_se), .CLK(
        CK), .Q(n7852), .QN(n3219) );
  sdffs1 \DFF_1488/Q_reg  ( .DIN(WX9919), .SDIN(n7850), .SSEL(test_se), .CLK(
        CK), .Q(n7851), .QN(n3220) );
  sdffs1 \DFF_1487/Q_reg  ( .DIN(WX9917), .SDIN(n7849), .SSEL(test_se), .CLK(
        CK), .Q(n7850), .QN(n6414) );
  sdffs1 \DFF_1486/Q_reg  ( .DIN(WX9915), .SDIN(n7848), .SSEL(test_se), .CLK(
        CK), .Q(n7849), .QN(n6412) );
  sdffs1 \DFF_1485/Q_reg  ( .DIN(WX9913), .SDIN(n7847), .SSEL(test_se), .CLK(
        CK), .Q(n7848), .QN(n6410) );
  sdffs1 \DFF_1484/Q_reg  ( .DIN(WX9911), .SDIN(n7846), .SSEL(test_se), .CLK(
        CK), .Q(n7847), .QN(n6408) );
  sdffs1 \DFF_1483/Q_reg  ( .DIN(WX9909), .SDIN(n7845), .SSEL(test_se), .CLK(
        CK), .Q(n7846), .QN(n6406) );
  sdffs1 \DFF_1482/Q_reg  ( .DIN(WX9907), .SDIN(n7844), .SSEL(test_se), .CLK(
        CK), .Q(n7845), .QN(n6404) );
  sdffs1 \DFF_1481/Q_reg  ( .DIN(WX9905), .SDIN(n7843), .SSEL(test_se), .CLK(
        CK), .Q(n7844), .QN(n6402) );
  sdffs1 \DFF_1480/Q_reg  ( .DIN(WX9903), .SDIN(n7842), .SSEL(test_se), .CLK(
        CK), .Q(n7843), .QN(n6400) );
  sdffs1 \DFF_1479/Q_reg  ( .DIN(WX9901), .SDIN(n7841), .SSEL(test_se), .CLK(
        CK), .Q(n7842), .QN(n6398) );
  sdffs1 \DFF_1478/Q_reg  ( .DIN(WX9899), .SDIN(n7840), .SSEL(test_se), .CLK(
        CK), .Q(n7841), .QN(n6396) );
  sdffs1 \DFF_1477/Q_reg  ( .DIN(WX9897), .SDIN(n7839), .SSEL(test_se), .CLK(
        CK), .Q(n7840), .QN(n6394) );
  sdffs1 \DFF_1476/Q_reg  ( .DIN(WX9895), .SDIN(n7838), .SSEL(test_se), .CLK(
        CK), .Q(n7839), .QN(n6392) );
  sdffs1 \DFF_1475/Q_reg  ( .DIN(WX9893), .SDIN(n7837), .SSEL(test_se), .CLK(
        CK), .Q(n7838), .QN(n6390) );
  sdffs1 \DFF_1474/Q_reg  ( .DIN(WX9891), .SDIN(n7836), .SSEL(test_se), .CLK(
        CK), .Q(n7837), .QN(n6388) );
  sdffs1 \DFF_1473/Q_reg  ( .DIN(WX9889), .SDIN(n7835), .SSEL(test_se), .CLK(
        CK), .Q(n7836), .QN(n6386) );
  sdffs1 \DFF_1472/Q_reg  ( .DIN(WX9887), .SDIN(n7834), .SSEL(test_se), .CLK(
        CK), .Q(n7835), .QN(n6384) );
  sdffs1 \DFF_1471/Q_reg  ( .DIN(WX9885), .SDIN(n7833), .SSEL(test_se), .CLK(
        CK), .Q(n7834), .QN(n4997) );
  sdffs1 \DFF_1470/Q_reg  ( .DIN(WX9883), .SDIN(n7832), .SSEL(test_se), .CLK(
        CK), .Q(n7833), .QN(n5001) );
  sdffs1 \DFF_1469/Q_reg  ( .DIN(WX9881), .SDIN(n7831), .SSEL(test_se), .CLK(
        CK), .Q(n7832), .QN(n5005) );
  sdffs1 \DFF_1468/Q_reg  ( .DIN(WX9879), .SDIN(n7830), .SSEL(test_se), .CLK(
        CK), .Q(n7831), .QN(n5009) );
  sdffs1 \DFF_1467/Q_reg  ( .DIN(WX9877), .SDIN(n7829), .SSEL(test_se), .CLK(
        CK), .Q(n7830), .QN(n5013) );
  sdffs1 \DFF_1466/Q_reg  ( .DIN(WX9875), .SDIN(n7828), .SSEL(test_se), .CLK(
        CK), .Q(n7829), .QN(n5017) );
  sdffs1 \DFF_1465/Q_reg  ( .DIN(WX9873), .SDIN(n7827), .SSEL(test_se), .CLK(
        CK), .Q(n7828), .QN(n5021) );
  sdffs1 \DFF_1464/Q_reg  ( .DIN(WX9871), .SDIN(n7826), .SSEL(test_se), .CLK(
        CK), .Q(n7827), .QN(n5025) );
  sdffs1 \DFF_1463/Q_reg  ( .DIN(WX9869), .SDIN(n7825), .SSEL(test_se), .CLK(
        CK), .Q(n7826), .QN(n5029) );
  sdffs1 \DFF_1462/Q_reg  ( .DIN(WX9867), .SDIN(n7824), .SSEL(test_se), .CLK(
        CK), .Q(n7825), .QN(n5033) );
  sdffs1 \DFF_1461/Q_reg  ( .DIN(WX9865), .SDIN(n7823), .SSEL(test_se), .CLK(
        CK), .Q(n7824), .QN(n5037) );
  sdffs1 \DFF_1460/Q_reg  ( .DIN(WX9863), .SDIN(n7822), .SSEL(test_se), .CLK(
        CK), .Q(n7823), .QN(n5041) );
  sdffs1 \DFF_1459/Q_reg  ( .DIN(WX9861), .SDIN(n7821), .SSEL(test_se), .CLK(
        CK), .Q(n7822), .QN(n5045) );
  sdffs1 \DFF_1458/Q_reg  ( .DIN(WX9859), .SDIN(n7820), .SSEL(test_se), .CLK(
        CK), .Q(n7821), .QN(n5049) );
  sdffs1 \DFF_1457/Q_reg  ( .DIN(WX9857), .SDIN(n7819), .SSEL(test_se), .CLK(
        CK), .Q(n7820), .QN(n5053) );
  sdffs1 \DFF_1456/Q_reg  ( .DIN(WX9855), .SDIN(n7818), .SSEL(test_se), .CLK(
        CK), .Q(n7819), .QN(n5057) );
  sdffs1 \DFF_1455/Q_reg  ( .DIN(WX9853), .SDIN(n7817), .SSEL(test_se), .CLK(
        CK), .Q(n7818), .QN(n5061) );
  sdffs1 \DFF_1454/Q_reg  ( .DIN(WX9851), .SDIN(n7816), .SSEL(test_se), .CLK(
        CK), .Q(n7817), .QN(n5065) );
  sdffs1 \DFF_1453/Q_reg  ( .DIN(WX9849), .SDIN(n7815), .SSEL(test_se), .CLK(
        CK), .Q(n7816), .QN(n5069) );
  sdffs1 \DFF_1452/Q_reg  ( .DIN(WX9847), .SDIN(n7814), .SSEL(test_se), .CLK(
        CK), .Q(n7815), .QN(n5073) );
  sdffs1 \DFF_1451/Q_reg  ( .DIN(WX9845), .SDIN(n7813), .SSEL(test_se), .CLK(
        CK), .Q(n7814), .QN(n5077) );
  sdffs1 \DFF_1450/Q_reg  ( .DIN(WX9843), .SDIN(n7812), .SSEL(test_se), .CLK(
        CK), .Q(n7813), .QN(n5081) );
  sdffs1 \DFF_1449/Q_reg  ( .DIN(WX9841), .SDIN(n7811), .SSEL(test_se), .CLK(
        CK), .Q(n7812), .QN(n5085) );
  sdffs1 \DFF_1448/Q_reg  ( .DIN(WX9839), .SDIN(n7810), .SSEL(test_se), .CLK(
        CK), .Q(n7811), .QN(n5089) );
  sdffs1 \DFF_1447/Q_reg  ( .DIN(WX9837), .SDIN(n7809), .SSEL(test_se), .CLK(
        CK), .Q(n7810), .QN(n5093) );
  sdffs1 \DFF_1446/Q_reg  ( .DIN(WX9835), .SDIN(n7808), .SSEL(test_se), .CLK(
        CK), .Q(n7809), .QN(n5097) );
  sdffs1 \DFF_1445/Q_reg  ( .DIN(WX9833), .SDIN(n7807), .SSEL(test_se), .CLK(
        CK), .Q(n7808), .QN(n5101) );
  sdffs1 \DFF_1444/Q_reg  ( .DIN(WX9831), .SDIN(n7806), .SSEL(test_se), .CLK(
        CK), .Q(n7807), .QN(n5105) );
  sdffs1 \DFF_1443/Q_reg  ( .DIN(WX9829), .SDIN(n7805), .SSEL(test_se), .CLK(
        CK), .Q(n7806), .QN(n5109) );
  sdffs1 \DFF_1442/Q_reg  ( .DIN(WX9827), .SDIN(n7804), .SSEL(test_se), .CLK(
        CK), .Q(n7805), .QN(n5113) );
  sdffs1 \DFF_1441/Q_reg  ( .DIN(WX9825), .SDIN(n7803), .SSEL(test_se), .CLK(
        CK), .Q(n7804), .QN(n5117) );
  sdffs1 \DFF_1440/Q_reg  ( .DIN(WX9823), .SDIN(n7802), .SSEL(test_se), .CLK(
        CK), .Q(n7803), .QN(n5121) );
  sdffs1 \DFF_1439/Q_reg  ( .DIN(WX9821), .SDIN(n7801), .SSEL(test_se), .CLK(
        CK), .Q(n7802), .QN(n4996) );
  sdffs1 \DFF_1438/Q_reg  ( .DIN(WX9819), .SDIN(n7800), .SSEL(test_se), .CLK(
        CK), .Q(n7801), .QN(n5000) );
  sdffs1 \DFF_1437/Q_reg  ( .DIN(WX9817), .SDIN(n7799), .SSEL(test_se), .CLK(
        CK), .Q(n7800), .QN(n5004) );
  sdffs1 \DFF_1436/Q_reg  ( .DIN(WX9815), .SDIN(n7798), .SSEL(test_se), .CLK(
        CK), .Q(n7799), .QN(n5008) );
  sdffs1 \DFF_1435/Q_reg  ( .DIN(WX9813), .SDIN(n7797), .SSEL(test_se), .CLK(
        CK), .Q(n7798), .QN(n5012) );
  sdffs1 \DFF_1434/Q_reg  ( .DIN(WX9811), .SDIN(n7796), .SSEL(test_se), .CLK(
        CK), .Q(n7797), .QN(n5016) );
  sdffs1 \DFF_1433/Q_reg  ( .DIN(WX9809), .SDIN(n7795), .SSEL(test_se), .CLK(
        CK), .Q(n7796), .QN(n5020) );
  sdffs1 \DFF_1432/Q_reg  ( .DIN(WX9807), .SDIN(n7794), .SSEL(test_se), .CLK(
        CK), .Q(n7795), .QN(n5024) );
  sdffs1 \DFF_1431/Q_reg  ( .DIN(WX9805), .SDIN(n7793), .SSEL(test_se), .CLK(
        CK), .Q(n7794), .QN(n5028) );
  sdffs1 \DFF_1430/Q_reg  ( .DIN(WX9803), .SDIN(n7792), .SSEL(test_se), .CLK(
        CK), .Q(n7793), .QN(n5032) );
  sdffs1 \DFF_1429/Q_reg  ( .DIN(WX9801), .SDIN(n7791), .SSEL(test_se), .CLK(
        CK), .Q(n7792), .QN(n5036) );
  sdffs1 \DFF_1428/Q_reg  ( .DIN(WX9799), .SDIN(n7790), .SSEL(test_se), .CLK(
        CK), .Q(n7791), .QN(n5040) );
  sdffs1 \DFF_1427/Q_reg  ( .DIN(WX9797), .SDIN(n7789), .SSEL(test_se), .CLK(
        CK), .Q(n7790), .QN(n5044) );
  sdffs1 \DFF_1426/Q_reg  ( .DIN(WX9795), .SDIN(n7788), .SSEL(test_se), .CLK(
        CK), .Q(n7789), .QN(n5048) );
  sdffs1 \DFF_1425/Q_reg  ( .DIN(WX9793), .SDIN(n7787), .SSEL(test_se), .CLK(
        CK), .Q(n7788), .QN(n5052) );
  sdffs1 \DFF_1424/Q_reg  ( .DIN(WX9791), .SDIN(n5060), .SSEL(test_se), .CLK(
        CK), .Q(n7787), .QN(n5056) );
  sdffs1 \DFF_1423/Q_reg  ( .DIN(WX9789), .SDIN(n5064), .SSEL(test_se), .CLK(
        CK), .Q(n5060) );
  sdffs1 \DFF_1422/Q_reg  ( .DIN(WX9787), .SDIN(n5068), .SSEL(test_se), .CLK(
        CK), .Q(n5064) );
  sdffs1 \DFF_1421/Q_reg  ( .DIN(WX9785), .SDIN(n5072), .SSEL(test_se), .CLK(
        CK), .Q(n5068) );
  sdffs1 \DFF_1420/Q_reg  ( .DIN(WX9783), .SDIN(n5076), .SSEL(test_se), .CLK(
        CK), .Q(n5072) );
  sdffs1 \DFF_1419/Q_reg  ( .DIN(WX9781), .SDIN(n5080), .SSEL(test_se), .CLK(
        CK), .Q(n5076) );
  sdffs1 \DFF_1418/Q_reg  ( .DIN(WX9779), .SDIN(n5084), .SSEL(test_se), .CLK(
        CK), .Q(n5080) );
  sdffs1 \DFF_1417/Q_reg  ( .DIN(WX9777), .SDIN(n5088), .SSEL(test_se), .CLK(
        CK), .Q(n5084) );
  sdffs1 \DFF_1416/Q_reg  ( .DIN(WX9775), .SDIN(n5092), .SSEL(test_se), .CLK(
        CK), .Q(n5088) );
  sdffs1 \DFF_1415/Q_reg  ( .DIN(WX9773), .SDIN(n5096), .SSEL(test_se), .CLK(
        CK), .Q(n5092) );
  sdffs1 \DFF_1414/Q_reg  ( .DIN(WX9771), .SDIN(n5100), .SSEL(test_se), .CLK(
        CK), .Q(n5096) );
  sdffs1 \DFF_1413/Q_reg  ( .DIN(WX9769), .SDIN(n5104), .SSEL(test_se), .CLK(
        CK), .Q(n5100) );
  sdffs1 \DFF_1412/Q_reg  ( .DIN(WX9767), .SDIN(n5108), .SSEL(test_se), .CLK(
        CK), .Q(n5104) );
  sdffs1 \DFF_1411/Q_reg  ( .DIN(WX9765), .SDIN(n5112), .SSEL(test_se), .CLK(
        CK), .Q(n5108) );
  sdffs1 \DFF_1410/Q_reg  ( .DIN(WX9763), .SDIN(n5116), .SSEL(test_se), .CLK(
        CK), .Q(n5112) );
  sdffs1 \DFF_1409/Q_reg  ( .DIN(WX9761), .SDIN(n5120), .SSEL(test_se), .CLK(
        CK), .Q(n5116) );
  sdffs1 \DFF_1408/Q_reg  ( .DIN(WX9759), .SDIN(n4995), .SSEL(test_se), .CLK(
        CK), .Q(n5120) );
  sdffs1 \DFF_1407/Q_reg  ( .DIN(WX9757), .SDIN(n4999), .SSEL(test_se), .CLK(
        CK), .Q(n4995) );
  sdffs1 \DFF_1406/Q_reg  ( .DIN(WX9755), .SDIN(n5003), .SSEL(test_se), .CLK(
        CK), .Q(n4999) );
  sdffs1 \DFF_1405/Q_reg  ( .DIN(WX9753), .SDIN(n5007), .SSEL(test_se), .CLK(
        CK), .Q(n5003) );
  sdffs1 \DFF_1404/Q_reg  ( .DIN(WX9751), .SDIN(n5011), .SSEL(test_se), .CLK(
        CK), .Q(n5007) );
  sdffs1 \DFF_1403/Q_reg  ( .DIN(WX9749), .SDIN(n5015), .SSEL(test_se), .CLK(
        CK), .Q(n5011) );
  sdffs1 \DFF_1402/Q_reg  ( .DIN(WX9747), .SDIN(n5019), .SSEL(test_se), .CLK(
        CK), .Q(n5015) );
  sdffs1 \DFF_1401/Q_reg  ( .DIN(WX9745), .SDIN(n5023), .SSEL(test_se), .CLK(
        CK), .Q(n5019) );
  sdffs1 \DFF_1400/Q_reg  ( .DIN(WX9743), .SDIN(n5027), .SSEL(test_se), .CLK(
        CK), .Q(n5023) );
  sdffs1 \DFF_1399/Q_reg  ( .DIN(WX9741), .SDIN(n5031), .SSEL(test_se), .CLK(
        CK), .Q(n5027) );
  sdffs1 \DFF_1398/Q_reg  ( .DIN(WX9739), .SDIN(n5035), .SSEL(test_se), .CLK(
        CK), .Q(n5031) );
  sdffs1 \DFF_1397/Q_reg  ( .DIN(WX9737), .SDIN(n5039), .SSEL(test_se), .CLK(
        CK), .Q(n5035) );
  sdffs1 \DFF_1396/Q_reg  ( .DIN(WX9735), .SDIN(n5043), .SSEL(test_se), .CLK(
        CK), .Q(n5039) );
  sdffs1 \DFF_1395/Q_reg  ( .DIN(WX9733), .SDIN(n5047), .SSEL(test_se), .CLK(
        CK), .Q(n5043) );
  sdffs1 \DFF_1394/Q_reg  ( .DIN(WX9731), .SDIN(n5051), .SSEL(test_se), .CLK(
        CK), .Q(n5047) );
  sdffs1 \DFF_1393/Q_reg  ( .DIN(WX9729), .SDIN(n5055), .SSEL(test_se), .CLK(
        CK), .Q(n5051) );
  sdffs1 \DFF_1392/Q_reg  ( .DIN(WX9727), .SDIN(n7786), .SSEL(test_se), .CLK(
        CK), .Q(n5055) );
  sdffs1 \DFF_1391/Q_reg  ( .DIN(WX9725), .SDIN(n7785), .SSEL(test_se), .CLK(
        CK), .Q(n7786), .QN(n5059) );
  sdffs1 \DFF_1390/Q_reg  ( .DIN(WX9723), .SDIN(n7784), .SSEL(test_se), .CLK(
        CK), .Q(n7785), .QN(n5063) );
  sdffs1 \DFF_1389/Q_reg  ( .DIN(WX9721), .SDIN(n7783), .SSEL(test_se), .CLK(
        CK), .Q(n7784), .QN(n5067) );
  sdffs1 \DFF_1388/Q_reg  ( .DIN(WX9719), .SDIN(n7782), .SSEL(test_se), .CLK(
        CK), .Q(n7783), .QN(n5071) );
  sdffs1 \DFF_1387/Q_reg  ( .DIN(WX9717), .SDIN(n7781), .SSEL(test_se), .CLK(
        CK), .Q(n7782), .QN(n5075) );
  sdffs1 \DFF_1386/Q_reg  ( .DIN(WX9715), .SDIN(n7780), .SSEL(test_se), .CLK(
        CK), .Q(n7781), .QN(n5079) );
  sdffs1 \DFF_1385/Q_reg  ( .DIN(WX9713), .SDIN(n7779), .SSEL(test_se), .CLK(
        CK), .Q(n7780), .QN(n5083) );
  sdffs1 \DFF_1384/Q_reg  ( .DIN(WX9711), .SDIN(n7778), .SSEL(test_se), .CLK(
        CK), .Q(n7779), .QN(n5087) );
  sdffs1 \DFF_1383/Q_reg  ( .DIN(WX9709), .SDIN(n7777), .SSEL(test_se), .CLK(
        CK), .Q(n7778), .QN(n5091) );
  sdffs1 \DFF_1382/Q_reg  ( .DIN(WX9707), .SDIN(n7776), .SSEL(test_se), .CLK(
        CK), .Q(n7777), .QN(n5095) );
  sdffs1 \DFF_1381/Q_reg  ( .DIN(WX9705), .SDIN(n7775), .SSEL(test_se), .CLK(
        CK), .Q(n7776), .QN(n5099) );
  sdffs1 \DFF_1380/Q_reg  ( .DIN(WX9703), .SDIN(n7774), .SSEL(test_se), .CLK(
        CK), .Q(n7775), .QN(n5103) );
  sdffs1 \DFF_1379/Q_reg  ( .DIN(WX9701), .SDIN(n7773), .SSEL(test_se), .CLK(
        CK), .Q(n7774), .QN(n5107) );
  sdffs1 \DFF_1378/Q_reg  ( .DIN(WX9699), .SDIN(n7772), .SSEL(test_se), .CLK(
        CK), .Q(n7773), .QN(n5111) );
  sdffs1 \DFF_1377/Q_reg  ( .DIN(WX9697), .SDIN(n7771), .SSEL(test_se), .CLK(
        CK), .Q(n7772), .QN(n5115) );
  sdffs1 \DFF_1376/Q_reg  ( .DIN(WX9695), .SDIN(n7770), .SSEL(test_se), .CLK(
        CK), .Q(n7771), .QN(n5119) );
  sdffs1 \DFF_1375/Q_reg  ( .DIN(WX9597), .SDIN(n7769), .SSEL(test_se), .CLK(
        CK), .Q(n7770), .QN(n4964) );
  sdffs1 \DFF_1374/Q_reg  ( .DIN(WX9595), .SDIN(n7768), .SSEL(test_se), .CLK(
        CK), .Q(n7769), .QN(n4965) );
  sdffs1 \DFF_1373/Q_reg  ( .DIN(WX9593), .SDIN(n7767), .SSEL(test_se), .CLK(
        CK), .Q(n7768), .QN(n4966) );
  sdffs1 \DFF_1372/Q_reg  ( .DIN(WX9591), .SDIN(n7766), .SSEL(test_se), .CLK(
        CK), .Q(n7767), .QN(n4967) );
  sdffs1 \DFF_1371/Q_reg  ( .DIN(WX9589), .SDIN(n7765), .SSEL(test_se), .CLK(
        CK), .Q(n7766), .QN(n4968) );
  sdffs1 \DFF_1370/Q_reg  ( .DIN(WX9587), .SDIN(n7764), .SSEL(test_se), .CLK(
        CK), .Q(n7765), .QN(n4969) );
  sdffs1 \DFF_1369/Q_reg  ( .DIN(WX9585), .SDIN(n7763), .SSEL(test_se), .CLK(
        CK), .Q(n7764), .QN(n4970) );
  sdffs1 \DFF_1368/Q_reg  ( .DIN(WX9583), .SDIN(n7762), .SSEL(test_se), .CLK(
        CK), .Q(n7763), .QN(n4971) );
  sdffs1 \DFF_1367/Q_reg  ( .DIN(WX9581), .SDIN(n7761), .SSEL(test_se), .CLK(
        CK), .Q(n7762), .QN(n4972) );
  sdffs1 \DFF_1366/Q_reg  ( .DIN(WX9579), .SDIN(n7760), .SSEL(test_se), .CLK(
        CK), .Q(n7761), .QN(n4973) );
  sdffs1 \DFF_1365/Q_reg  ( .DIN(WX9577), .SDIN(n7759), .SSEL(test_se), .CLK(
        CK), .Q(n7760), .QN(n4974) );
  sdffs1 \DFF_1364/Q_reg  ( .DIN(WX9575), .SDIN(n7758), .SSEL(test_se), .CLK(
        CK), .Q(n7759), .QN(n4975) );
  sdffs1 \DFF_1363/Q_reg  ( .DIN(WX9573), .SDIN(n7757), .SSEL(test_se), .CLK(
        CK), .Q(n7758), .QN(n4976) );
  sdffs1 \DFF_1362/Q_reg  ( .DIN(WX9571), .SDIN(n7756), .SSEL(test_se), .CLK(
        CK), .Q(n7757), .QN(n4977) );
  sdffs1 \DFF_1361/Q_reg  ( .DIN(WX9569), .SDIN(n7755), .SSEL(test_se), .CLK(
        CK), .Q(n7756), .QN(n4978) );
  sdffs1 \DFF_1360/Q_reg  ( .DIN(WX9567), .SDIN(n7754), .SSEL(test_se), .CLK(
        CK), .Q(n7755), .QN(n4979) );
  sdffs1 \DFF_1359/Q_reg  ( .DIN(WX9565), .SDIN(n7753), .SSEL(test_se), .CLK(
        CK), .Q(n7754), .QN(n4980) );
  sdffs1 \DFF_1358/Q_reg  ( .DIN(WX9563), .SDIN(n7752), .SSEL(test_se), .CLK(
        CK), .Q(n7753), .QN(n4981) );
  sdffs1 \DFF_1357/Q_reg  ( .DIN(WX9561), .SDIN(n7751), .SSEL(test_se), .CLK(
        CK), .Q(n7752), .QN(n4982) );
  sdffs1 \DFF_1356/Q_reg  ( .DIN(WX9559), .SDIN(n7750), .SSEL(test_se), .CLK(
        CK), .Q(n7751), .QN(n4983) );
  sdffs1 \DFF_1355/Q_reg  ( .DIN(WX9557), .SDIN(n7749), .SSEL(test_se), .CLK(
        CK), .Q(n7750), .QN(n4984) );
  sdffs1 \DFF_1354/Q_reg  ( .DIN(WX9555), .SDIN(n7748), .SSEL(test_se), .CLK(
        CK), .Q(n7749), .QN(n4985) );
  sdffs1 \DFF_1353/Q_reg  ( .DIN(WX9553), .SDIN(n7747), .SSEL(test_se), .CLK(
        CK), .Q(n7748), .QN(n4986) );
  sdffs1 \DFF_1352/Q_reg  ( .DIN(WX9551), .SDIN(n7746), .SSEL(test_se), .CLK(
        CK), .Q(n7747), .QN(n4987) );
  sdffs1 \DFF_1351/Q_reg  ( .DIN(WX9549), .SDIN(n7745), .SSEL(test_se), .CLK(
        CK), .Q(n7746), .QN(n4988) );
  sdffs1 \DFF_1350/Q_reg  ( .DIN(WX9547), .SDIN(n7744), .SSEL(test_se), .CLK(
        CK), .Q(n7745), .QN(n4989) );
  sdffs1 \DFF_1349/Q_reg  ( .DIN(WX9545), .SDIN(n7743), .SSEL(test_se), .CLK(
        CK), .Q(n7744), .QN(n4990) );
  sdffs1 \DFF_1348/Q_reg  ( .DIN(WX9543), .SDIN(n7742), .SSEL(test_se), .CLK(
        CK), .Q(n7743), .QN(n4991) );
  sdffs1 \DFF_1347/Q_reg  ( .DIN(WX9541), .SDIN(n7741), .SSEL(test_se), .CLK(
        CK), .Q(n7742), .QN(n4992) );
  sdffs1 \DFF_1346/Q_reg  ( .DIN(WX9539), .SDIN(n7740), .SSEL(test_se), .CLK(
        CK), .Q(n7741), .QN(n4993) );
  sdffs1 \DFF_1345/Q_reg  ( .DIN(WX9537), .SDIN(n7739), .SSEL(test_se), .CLK(
        CK), .Q(n7740), .QN(n4994) );
  sdffs1 \DFF_1344/Q_reg  ( .DIN(WX9535), .SDIN(CRC_OUT_3_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7739), .QN(n4963) );
  sdffs1 \DFF_1343/Q_reg  ( .DIN(WX9084), .SDIN(CRC_OUT_3_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_31), .QN(n5122) );
  sdffs1 \DFF_1342/Q_reg  ( .DIN(WX9082), .SDIN(CRC_OUT_3_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_30), .QN(n5118) );
  sdffs1 \DFF_1341/Q_reg  ( .DIN(WX9080), .SDIN(CRC_OUT_3_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_29), .QN(n5114) );
  sdffs1 \DFF_1340/Q_reg  ( .DIN(WX9078), .SDIN(CRC_OUT_3_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_28), .QN(n5110) );
  sdffs1 \DFF_1339/Q_reg  ( .DIN(WX9076), .SDIN(CRC_OUT_3_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_27), .QN(n5106) );
  sdffs1 \DFF_1338/Q_reg  ( .DIN(WX9074), .SDIN(CRC_OUT_3_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_26), .QN(n5102) );
  sdffs1 \DFF_1337/Q_reg  ( .DIN(WX9072), .SDIN(CRC_OUT_3_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_25), .QN(n5098) );
  sdffs1 \DFF_1336/Q_reg  ( .DIN(WX9070), .SDIN(CRC_OUT_3_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_24), .QN(n5094) );
  sdffs1 \DFF_1335/Q_reg  ( .DIN(WX9068), .SDIN(CRC_OUT_3_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_23), .QN(n5090) );
  sdffs1 \DFF_1334/Q_reg  ( .DIN(WX9066), .SDIN(CRC_OUT_3_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_22), .QN(n5086) );
  sdffs1 \DFF_1333/Q_reg  ( .DIN(WX9064), .SDIN(CRC_OUT_3_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_21), .QN(n5082) );
  sdffs1 \DFF_1332/Q_reg  ( .DIN(WX9062), .SDIN(CRC_OUT_3_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_20), .QN(n5078) );
  sdffs1 \DFF_1331/Q_reg  ( .DIN(WX9060), .SDIN(CRC_OUT_3_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_19), .QN(n5074) );
  sdffs1 \DFF_1330/Q_reg  ( .DIN(WX9058), .SDIN(CRC_OUT_3_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_18), .QN(n5070) );
  sdffs1 \DFF_1329/Q_reg  ( .DIN(WX9056), .SDIN(CRC_OUT_3_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_17), .QN(n5066) );
  sdffs1 \DFF_1328/Q_reg  ( .DIN(WX9054), .SDIN(CRC_OUT_3_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_16), .QN(n5062) );
  sdffs1 \DFF_1327/Q_reg  ( .DIN(WX9052), .SDIN(CRC_OUT_3_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_15), .QN(n5058) );
  sdffs1 \DFF_1326/Q_reg  ( .DIN(WX9050), .SDIN(CRC_OUT_3_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_14), .QN(n5054) );
  sdffs1 \DFF_1325/Q_reg  ( .DIN(WX9048), .SDIN(CRC_OUT_3_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_13), .QN(n5050) );
  sdffs1 \DFF_1324/Q_reg  ( .DIN(WX9046), .SDIN(CRC_OUT_3_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_12), .QN(n5046) );
  sdffs1 \DFF_1323/Q_reg  ( .DIN(WX9044), .SDIN(CRC_OUT_3_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_11), .QN(n5042) );
  sdffs1 \DFF_1322/Q_reg  ( .DIN(WX9042), .SDIN(CRC_OUT_3_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_10), .QN(n5038) );
  sdffs1 \DFF_1321/Q_reg  ( .DIN(WX9040), .SDIN(CRC_OUT_3_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_9), .QN(n5034) );
  sdffs1 \DFF_1320/Q_reg  ( .DIN(WX9038), .SDIN(CRC_OUT_3_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_8), .QN(n5030) );
  sdffs1 \DFF_1319/Q_reg  ( .DIN(WX9036), .SDIN(CRC_OUT_3_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_7), .QN(n5026) );
  sdffs1 \DFF_1318/Q_reg  ( .DIN(WX9034), .SDIN(CRC_OUT_3_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_6), .QN(n5022) );
  sdffs1 \DFF_1317/Q_reg  ( .DIN(WX9032), .SDIN(CRC_OUT_3_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_5), .QN(n5018) );
  sdffs1 \DFF_1316/Q_reg  ( .DIN(WX9030), .SDIN(CRC_OUT_3_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_4), .QN(n5014) );
  sdffs1 \DFF_1315/Q_reg  ( .DIN(WX9028), .SDIN(CRC_OUT_3_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_3), .QN(n5010) );
  sdffs1 \DFF_1314/Q_reg  ( .DIN(WX9026), .SDIN(CRC_OUT_3_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_2), .QN(n5006) );
  sdffs1 \DFF_1313/Q_reg  ( .DIN(WX9024), .SDIN(CRC_OUT_3_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_3_1), .QN(n5002) );
  sdffs1 \DFF_1312/Q_reg  ( .DIN(WX9022), .SDIN(n7738), .SSEL(test_se), .CLK(
        CK), .Q(CRC_OUT_3_0), .QN(n4998) );
  sdffs1 \DFF_1311/Q_reg  ( .DIN(WX8656), .SDIN(n7737), .SSEL(test_se), .CLK(
        CK), .Q(n7738), .QN(n3221) );
  sdffs1 \DFF_1310/Q_reg  ( .DIN(WX8654), .SDIN(n7736), .SSEL(test_se), .CLK(
        CK), .Q(n7737), .QN(n3222) );
  sdffs1 \DFF_1309/Q_reg  ( .DIN(WX8652), .SDIN(n7735), .SSEL(test_se), .CLK(
        CK), .Q(n7736), .QN(n3223) );
  sdffs1 \DFF_1308/Q_reg  ( .DIN(WX8650), .SDIN(n7734), .SSEL(test_se), .CLK(
        CK), .Q(n7735), .QN(n3224) );
  sdffs1 \DFF_1307/Q_reg  ( .DIN(WX8648), .SDIN(n7733), .SSEL(test_se), .CLK(
        CK), .Q(n7734), .QN(n3225) );
  sdffs1 \DFF_1306/Q_reg  ( .DIN(WX8646), .SDIN(n7732), .SSEL(test_se), .CLK(
        CK), .Q(n7733), .QN(n3226) );
  sdffs1 \DFF_1305/Q_reg  ( .DIN(WX8644), .SDIN(n7731), .SSEL(test_se), .CLK(
        CK), .Q(n7732), .QN(n3227) );
  sdffs1 \DFF_1304/Q_reg  ( .DIN(WX8642), .SDIN(n7730), .SSEL(test_se), .CLK(
        CK), .Q(n7731), .QN(n3228) );
  sdffs1 \DFF_1303/Q_reg  ( .DIN(WX8640), .SDIN(n7729), .SSEL(test_se), .CLK(
        CK), .Q(n7730), .QN(n3229) );
  sdffs1 \DFF_1302/Q_reg  ( .DIN(WX8638), .SDIN(n7728), .SSEL(test_se), .CLK(
        CK), .Q(n7729), .QN(n3230) );
  sdffs1 \DFF_1301/Q_reg  ( .DIN(WX8636), .SDIN(n7727), .SSEL(test_se), .CLK(
        CK), .Q(n7728), .QN(n3231) );
  sdffs1 \DFF_1300/Q_reg  ( .DIN(WX8634), .SDIN(n7726), .SSEL(test_se), .CLK(
        CK), .Q(n7727), .QN(n3232) );
  sdffs1 \DFF_1299/Q_reg  ( .DIN(WX8632), .SDIN(n7725), .SSEL(test_se), .CLK(
        CK), .Q(n7726), .QN(n3233) );
  sdffs1 \DFF_1298/Q_reg  ( .DIN(WX8630), .SDIN(n7724), .SSEL(test_se), .CLK(
        CK), .Q(n7725), .QN(n3234) );
  sdffs1 \DFF_1297/Q_reg  ( .DIN(WX8628), .SDIN(n7723), .SSEL(test_se), .CLK(
        CK), .Q(n7724), .QN(n3235) );
  sdffs1 \DFF_1296/Q_reg  ( .DIN(WX8626), .SDIN(n7722), .SSEL(test_se), .CLK(
        CK), .Q(n7723), .QN(n3236) );
  sdffs1 \DFF_1295/Q_reg  ( .DIN(WX8624), .SDIN(n7721), .SSEL(test_se), .CLK(
        CK), .Q(n7722), .QN(n5222) );
  sdffs1 \DFF_1294/Q_reg  ( .DIN(WX8622), .SDIN(n7720), .SSEL(test_se), .CLK(
        CK), .Q(n7721), .QN(n5227) );
  sdffs1 \DFF_1293/Q_reg  ( .DIN(WX8620), .SDIN(n7719), .SSEL(test_se), .CLK(
        CK), .Q(n7720), .QN(n5232) );
  sdffs1 \DFF_1292/Q_reg  ( .DIN(WX8618), .SDIN(n7718), .SSEL(test_se), .CLK(
        CK), .Q(n7719), .QN(n5237) );
  sdffs1 \DFF_1291/Q_reg  ( .DIN(WX8616), .SDIN(n7717), .SSEL(test_se), .CLK(
        CK), .Q(n7718), .QN(n5242) );
  sdffs1 \DFF_1290/Q_reg  ( .DIN(WX8614), .SDIN(n7716), .SSEL(test_se), .CLK(
        CK), .Q(n7717), .QN(n5247) );
  sdffs1 \DFF_1289/Q_reg  ( .DIN(WX8612), .SDIN(n7715), .SSEL(test_se), .CLK(
        CK), .Q(n7716), .QN(n5252) );
  sdffs1 \DFF_1288/Q_reg  ( .DIN(WX8610), .SDIN(n7714), .SSEL(test_se), .CLK(
        CK), .Q(n7715), .QN(n5257) );
  sdffs1 \DFF_1287/Q_reg  ( .DIN(WX8608), .SDIN(n7713), .SSEL(test_se), .CLK(
        CK), .Q(n7714), .QN(n5262) );
  sdffs1 \DFF_1286/Q_reg  ( .DIN(WX8606), .SDIN(n7712), .SSEL(test_se), .CLK(
        CK), .Q(n7713), .QN(n5267) );
  sdffs1 \DFF_1285/Q_reg  ( .DIN(WX8604), .SDIN(n7711), .SSEL(test_se), .CLK(
        CK), .Q(n7712), .QN(n5272) );
  sdffs1 \DFF_1284/Q_reg  ( .DIN(WX8602), .SDIN(n7710), .SSEL(test_se), .CLK(
        CK), .Q(n7711), .QN(n5277) );
  sdffs1 \DFF_1283/Q_reg  ( .DIN(WX8600), .SDIN(n7709), .SSEL(test_se), .CLK(
        CK), .Q(n7710), .QN(n5282) );
  sdffs1 \DFF_1282/Q_reg  ( .DIN(WX8598), .SDIN(n7708), .SSEL(test_se), .CLK(
        CK), .Q(n7709), .QN(n5287) );
  sdffs1 \DFF_1281/Q_reg  ( .DIN(WX8596), .SDIN(n7707), .SSEL(test_se), .CLK(
        CK), .Q(n7708), .QN(n5292) );
  sdffs1 \DFF_1280/Q_reg  ( .DIN(WX8594), .SDIN(n7706), .SSEL(test_se), .CLK(
        CK), .Q(n7707), .QN(n5297) );
  sdffs1 \DFF_1279/Q_reg  ( .DIN(WX8592), .SDIN(n7705), .SSEL(test_se), .CLK(
        CK), .Q(n7706), .QN(n5157) );
  sdffs1 \DFF_1278/Q_reg  ( .DIN(WX8590), .SDIN(n7704), .SSEL(test_se), .CLK(
        CK), .Q(n7705), .QN(n5161) );
  sdffs1 \DFF_1277/Q_reg  ( .DIN(WX8588), .SDIN(n7703), .SSEL(test_se), .CLK(
        CK), .Q(n7704), .QN(n5165) );
  sdffs1 \DFF_1276/Q_reg  ( .DIN(WX8586), .SDIN(n7702), .SSEL(test_se), .CLK(
        CK), .Q(n7703), .QN(n5169) );
  sdffs1 \DFF_1275/Q_reg  ( .DIN(WX8584), .SDIN(n7701), .SSEL(test_se), .CLK(
        CK), .Q(n7702), .QN(n5173) );
  sdffs1 \DFF_1274/Q_reg  ( .DIN(WX8582), .SDIN(n7700), .SSEL(test_se), .CLK(
        CK), .Q(n7701), .QN(n5177) );
  sdffs1 \DFF_1273/Q_reg  ( .DIN(WX8580), .SDIN(n7699), .SSEL(test_se), .CLK(
        CK), .Q(n7700), .QN(n5181) );
  sdffs1 \DFF_1272/Q_reg  ( .DIN(WX8578), .SDIN(n7698), .SSEL(test_se), .CLK(
        CK), .Q(n7699), .QN(n5185) );
  sdffs1 \DFF_1271/Q_reg  ( .DIN(WX8576), .SDIN(n7697), .SSEL(test_se), .CLK(
        CK), .Q(n7698), .QN(n5189) );
  sdffs1 \DFF_1270/Q_reg  ( .DIN(WX8574), .SDIN(n7696), .SSEL(test_se), .CLK(
        CK), .Q(n7697), .QN(n5193) );
  sdffs1 \DFF_1269/Q_reg  ( .DIN(WX8572), .SDIN(n7695), .SSEL(test_se), .CLK(
        CK), .Q(n7696), .QN(n5197) );
  sdffs1 \DFF_1268/Q_reg  ( .DIN(WX8570), .SDIN(n7694), .SSEL(test_se), .CLK(
        CK), .Q(n7695), .QN(n5201) );
  sdffs1 \DFF_1267/Q_reg  ( .DIN(WX8568), .SDIN(n7693), .SSEL(test_se), .CLK(
        CK), .Q(n7694), .QN(n5205) );
  sdffs1 \DFF_1266/Q_reg  ( .DIN(WX8566), .SDIN(n7692), .SSEL(test_se), .CLK(
        CK), .Q(n7693), .QN(n5209) );
  sdffs1 \DFF_1265/Q_reg  ( .DIN(WX8564), .SDIN(n7691), .SSEL(test_se), .CLK(
        CK), .Q(n7692), .QN(n5213) );
  sdffs1 \DFF_1264/Q_reg  ( .DIN(WX8562), .SDIN(n7690), .SSEL(test_se), .CLK(
        CK), .Q(n7691), .QN(n5217) );
  sdffs1 \DFF_1263/Q_reg  ( .DIN(WX8560), .SDIN(n7689), .SSEL(test_se), .CLK(
        CK), .Q(n7690), .QN(n5221) );
  sdffs1 \DFF_1262/Q_reg  ( .DIN(WX8558), .SDIN(n7688), .SSEL(test_se), .CLK(
        CK), .Q(n7689), .QN(n5226) );
  sdffs1 \DFF_1261/Q_reg  ( .DIN(WX8556), .SDIN(n7687), .SSEL(test_se), .CLK(
        CK), .Q(n7688), .QN(n5231) );
  sdffs1 \DFF_1260/Q_reg  ( .DIN(WX8554), .SDIN(n7686), .SSEL(test_se), .CLK(
        CK), .Q(n7687), .QN(n5236) );
  sdffs1 \DFF_1259/Q_reg  ( .DIN(WX8552), .SDIN(n7685), .SSEL(test_se), .CLK(
        CK), .Q(n7686), .QN(n5241) );
  sdffs1 \DFF_1258/Q_reg  ( .DIN(WX8550), .SDIN(n7684), .SSEL(test_se), .CLK(
        CK), .Q(n7685), .QN(n5246) );
  sdffs1 \DFF_1257/Q_reg  ( .DIN(WX8548), .SDIN(n7683), .SSEL(test_se), .CLK(
        CK), .Q(n7684), .QN(n5251) );
  sdffs1 \DFF_1256/Q_reg  ( .DIN(WX8546), .SDIN(n7682), .SSEL(test_se), .CLK(
        CK), .Q(n7683), .QN(n5256) );
  sdffs1 \DFF_1255/Q_reg  ( .DIN(WX8544), .SDIN(n7681), .SSEL(test_se), .CLK(
        CK), .Q(n7682), .QN(n5261) );
  sdffs1 \DFF_1254/Q_reg  ( .DIN(WX8542), .SDIN(n7680), .SSEL(test_se), .CLK(
        CK), .Q(n7681), .QN(n5266) );
  sdffs1 \DFF_1253/Q_reg  ( .DIN(WX8540), .SDIN(n7679), .SSEL(test_se), .CLK(
        CK), .Q(n7680), .QN(n5271) );
  sdffs1 \DFF_1252/Q_reg  ( .DIN(WX8538), .SDIN(n7678), .SSEL(test_se), .CLK(
        CK), .Q(n7679), .QN(n5276) );
  sdffs1 \DFF_1251/Q_reg  ( .DIN(WX8536), .SDIN(n7677), .SSEL(test_se), .CLK(
        CK), .Q(n7678), .QN(n5281) );
  sdffs1 \DFF_1250/Q_reg  ( .DIN(WX8534), .SDIN(n7676), .SSEL(test_se), .CLK(
        CK), .Q(n7677), .QN(n5286) );
  sdffs1 \DFF_1249/Q_reg  ( .DIN(WX8532), .SDIN(n7675), .SSEL(test_se), .CLK(
        CK), .Q(n7676), .QN(n5291) );
  sdffs1 \DFF_1248/Q_reg  ( .DIN(WX8530), .SDIN(n7674), .SSEL(test_se), .CLK(
        CK), .Q(n7675), .QN(n5296) );
  sdffs1 \DFF_1247/Q_reg  ( .DIN(WX8528), .SDIN(n7673), .SSEL(test_se), .CLK(
        CK), .Q(n7674), .QN(n5156) );
  sdffs1 \DFF_1246/Q_reg  ( .DIN(WX8526), .SDIN(n7672), .SSEL(test_se), .CLK(
        CK), .Q(n7673), .QN(n5160) );
  sdffs1 \DFF_1245/Q_reg  ( .DIN(WX8524), .SDIN(n7671), .SSEL(test_se), .CLK(
        CK), .Q(n7672), .QN(n5164) );
  sdffs1 \DFF_1244/Q_reg  ( .DIN(WX8522), .SDIN(n7670), .SSEL(test_se), .CLK(
        CK), .Q(n7671), .QN(n5168) );
  sdffs1 \DFF_1243/Q_reg  ( .DIN(WX8520), .SDIN(n7669), .SSEL(test_se), .CLK(
        CK), .Q(n7670), .QN(n5172) );
  sdffs1 \DFF_1242/Q_reg  ( .DIN(WX8518), .SDIN(n7668), .SSEL(test_se), .CLK(
        CK), .Q(n7669), .QN(n5176) );
  sdffs1 \DFF_1241/Q_reg  ( .DIN(WX8516), .SDIN(n7667), .SSEL(test_se), .CLK(
        CK), .Q(n7668), .QN(n5180) );
  sdffs1 \DFF_1240/Q_reg  ( .DIN(WX8514), .SDIN(n7666), .SSEL(test_se), .CLK(
        CK), .Q(n7667), .QN(n5184) );
  sdffs1 \DFF_1239/Q_reg  ( .DIN(WX8512), .SDIN(n7665), .SSEL(test_se), .CLK(
        CK), .Q(n7666), .QN(n5188) );
  sdffs1 \DFF_1238/Q_reg  ( .DIN(WX8510), .SDIN(n7664), .SSEL(test_se), .CLK(
        CK), .Q(n7665), .QN(n5192) );
  sdffs1 \DFF_1237/Q_reg  ( .DIN(WX8508), .SDIN(n7663), .SSEL(test_se), .CLK(
        CK), .Q(n7664), .QN(n5196) );
  sdffs1 \DFF_1236/Q_reg  ( .DIN(WX8506), .SDIN(n7662), .SSEL(test_se), .CLK(
        CK), .Q(n7663), .QN(n5200) );
  sdffs1 \DFF_1235/Q_reg  ( .DIN(WX8504), .SDIN(n7661), .SSEL(test_se), .CLK(
        CK), .Q(n7662), .QN(n5204) );
  sdffs1 \DFF_1234/Q_reg  ( .DIN(WX8502), .SDIN(n7660), .SSEL(test_se), .CLK(
        CK), .Q(n7661), .QN(n5208) );
  sdffs1 \DFF_1233/Q_reg  ( .DIN(WX8500), .SDIN(n7659), .SSEL(test_se), .CLK(
        CK), .Q(n7660), .QN(n5212) );
  sdffs1 \DFF_1232/Q_reg  ( .DIN(WX8498), .SDIN(n5220), .SSEL(test_se), .CLK(
        CK), .Q(n7659), .QN(n5216) );
  sdffs1 \DFF_1231/Q_reg  ( .DIN(WX8496), .SDIN(n5225), .SSEL(test_se), .CLK(
        CK), .Q(n5220) );
  sdffs1 \DFF_1230/Q_reg  ( .DIN(WX8494), .SDIN(n5230), .SSEL(test_se), .CLK(
        CK), .Q(n5225) );
  sdffs1 \DFF_1229/Q_reg  ( .DIN(WX8492), .SDIN(n5235), .SSEL(test_se), .CLK(
        CK), .Q(n5230) );
  sdffs1 \DFF_1228/Q_reg  ( .DIN(WX8490), .SDIN(n5240), .SSEL(test_se), .CLK(
        CK), .Q(n5235) );
  sdffs1 \DFF_1227/Q_reg  ( .DIN(WX8488), .SDIN(n5245), .SSEL(test_se), .CLK(
        CK), .Q(n5240) );
  sdffs1 \DFF_1226/Q_reg  ( .DIN(WX8486), .SDIN(n5250), .SSEL(test_se), .CLK(
        CK), .Q(n5245) );
  sdffs1 \DFF_1225/Q_reg  ( .DIN(WX8484), .SDIN(n5255), .SSEL(test_se), .CLK(
        CK), .Q(n5250) );
  sdffs1 \DFF_1224/Q_reg  ( .DIN(WX8482), .SDIN(n5260), .SSEL(test_se), .CLK(
        CK), .Q(n5255) );
  sdffs1 \DFF_1223/Q_reg  ( .DIN(WX8480), .SDIN(n5265), .SSEL(test_se), .CLK(
        CK), .Q(n5260) );
  sdffs1 \DFF_1222/Q_reg  ( .DIN(WX8478), .SDIN(n5270), .SSEL(test_se), .CLK(
        CK), .Q(n5265) );
  sdffs1 \DFF_1221/Q_reg  ( .DIN(WX8476), .SDIN(n5275), .SSEL(test_se), .CLK(
        CK), .Q(n5270) );
  sdffs1 \DFF_1220/Q_reg  ( .DIN(WX8474), .SDIN(n5280), .SSEL(test_se), .CLK(
        CK), .Q(n5275) );
  sdffs1 \DFF_1219/Q_reg  ( .DIN(WX8472), .SDIN(n5285), .SSEL(test_se), .CLK(
        CK), .Q(n5280) );
  sdffs1 \DFF_1218/Q_reg  ( .DIN(WX8470), .SDIN(n5290), .SSEL(test_se), .CLK(
        CK), .Q(n5285) );
  sdffs1 \DFF_1217/Q_reg  ( .DIN(WX8468), .SDIN(n5295), .SSEL(test_se), .CLK(
        CK), .Q(n5290) );
  sdffs1 \DFF_1216/Q_reg  ( .DIN(WX8466), .SDIN(n5155), .SSEL(test_se), .CLK(
        CK), .Q(n5295) );
  sdffs1 \DFF_1215/Q_reg  ( .DIN(WX8464), .SDIN(n5159), .SSEL(test_se), .CLK(
        CK), .Q(n5155) );
  sdffs1 \DFF_1214/Q_reg  ( .DIN(WX8462), .SDIN(n5163), .SSEL(test_se), .CLK(
        CK), .Q(n5159) );
  sdffs1 \DFF_1213/Q_reg  ( .DIN(WX8460), .SDIN(n5167), .SSEL(test_se), .CLK(
        CK), .Q(n5163) );
  sdffs1 \DFF_1212/Q_reg  ( .DIN(WX8458), .SDIN(n5171), .SSEL(test_se), .CLK(
        CK), .Q(n5167) );
  sdffs1 \DFF_1211/Q_reg  ( .DIN(WX8456), .SDIN(n5175), .SSEL(test_se), .CLK(
        CK), .Q(n5171) );
  sdffs1 \DFF_1210/Q_reg  ( .DIN(WX8454), .SDIN(n5179), .SSEL(test_se), .CLK(
        CK), .Q(n5175) );
  sdffs1 \DFF_1209/Q_reg  ( .DIN(WX8452), .SDIN(n5183), .SSEL(test_se), .CLK(
        CK), .Q(n5179) );
  sdffs1 \DFF_1208/Q_reg  ( .DIN(WX8450), .SDIN(n5187), .SSEL(test_se), .CLK(
        CK), .Q(n5183) );
  sdffs1 \DFF_1207/Q_reg  ( .DIN(WX8448), .SDIN(n5191), .SSEL(test_se), .CLK(
        CK), .Q(n5187) );
  sdffs1 \DFF_1206/Q_reg  ( .DIN(WX8446), .SDIN(n5195), .SSEL(test_se), .CLK(
        CK), .Q(n5191) );
  sdffs1 \DFF_1205/Q_reg  ( .DIN(WX8444), .SDIN(n5199), .SSEL(test_se), .CLK(
        CK), .Q(n5195) );
  sdffs1 \DFF_1204/Q_reg  ( .DIN(WX8442), .SDIN(n5203), .SSEL(test_se), .CLK(
        CK), .Q(n5199) );
  sdffs1 \DFF_1203/Q_reg  ( .DIN(WX8440), .SDIN(n5207), .SSEL(test_se), .CLK(
        CK), .Q(n5203) );
  sdffs1 \DFF_1202/Q_reg  ( .DIN(WX8438), .SDIN(n5211), .SSEL(test_se), .CLK(
        CK), .Q(n5207) );
  sdffs1 \DFF_1201/Q_reg  ( .DIN(WX8436), .SDIN(n5215), .SSEL(test_se), .CLK(
        CK), .Q(n5211) );
  sdffs1 \DFF_1200/Q_reg  ( .DIN(WX8434), .SDIN(n7658), .SSEL(test_se), .CLK(
        CK), .Q(n5215) );
  sdffs1 \DFF_1199/Q_reg  ( .DIN(WX8432), .SDIN(n7657), .SSEL(test_se), .CLK(
        CK), .Q(n7658), .QN(n5219) );
  sdffs1 \DFF_1198/Q_reg  ( .DIN(WX8430), .SDIN(n7656), .SSEL(test_se), .CLK(
        CK), .Q(n7657), .QN(n5224) );
  sdffs1 \DFF_1197/Q_reg  ( .DIN(WX8428), .SDIN(n7655), .SSEL(test_se), .CLK(
        CK), .Q(n7656), .QN(n5229) );
  sdffs1 \DFF_1196/Q_reg  ( .DIN(WX8426), .SDIN(n7654), .SSEL(test_se), .CLK(
        CK), .Q(n7655), .QN(n5234) );
  sdffs1 \DFF_1195/Q_reg  ( .DIN(WX8424), .SDIN(n7653), .SSEL(test_se), .CLK(
        CK), .Q(n7654), .QN(n5239) );
  sdffs1 \DFF_1194/Q_reg  ( .DIN(WX8422), .SDIN(n7652), .SSEL(test_se), .CLK(
        CK), .Q(n7653), .QN(n5244) );
  sdffs1 \DFF_1193/Q_reg  ( .DIN(WX8420), .SDIN(n7651), .SSEL(test_se), .CLK(
        CK), .Q(n7652), .QN(n5249) );
  sdffs1 \DFF_1192/Q_reg  ( .DIN(WX8418), .SDIN(n7650), .SSEL(test_se), .CLK(
        CK), .Q(n7651), .QN(n5254) );
  sdffs1 \DFF_1191/Q_reg  ( .DIN(WX8416), .SDIN(n7649), .SSEL(test_se), .CLK(
        CK), .Q(n7650), .QN(n5259) );
  sdffs1 \DFF_1190/Q_reg  ( .DIN(WX8414), .SDIN(n7648), .SSEL(test_se), .CLK(
        CK), .Q(n7649), .QN(n5264) );
  sdffs1 \DFF_1189/Q_reg  ( .DIN(WX8412), .SDIN(n7647), .SSEL(test_se), .CLK(
        CK), .Q(n7648), .QN(n5269) );
  sdffs1 \DFF_1188/Q_reg  ( .DIN(WX8410), .SDIN(n7646), .SSEL(test_se), .CLK(
        CK), .Q(n7647), .QN(n5274) );
  sdffs1 \DFF_1187/Q_reg  ( .DIN(WX8408), .SDIN(n7645), .SSEL(test_se), .CLK(
        CK), .Q(n7646), .QN(n5279) );
  sdffs1 \DFF_1186/Q_reg  ( .DIN(WX8406), .SDIN(n7644), .SSEL(test_se), .CLK(
        CK), .Q(n7645), .QN(n5284) );
  sdffs1 \DFF_1185/Q_reg  ( .DIN(WX8404), .SDIN(n7643), .SSEL(test_se), .CLK(
        CK), .Q(n7644), .QN(n5289) );
  sdffs1 \DFF_1184/Q_reg  ( .DIN(WX8402), .SDIN(n7642), .SSEL(test_se), .CLK(
        CK), .Q(n7643), .QN(n5294) );
  sdffs1 \DFF_1183/Q_reg  ( .DIN(WX8304), .SDIN(n7641), .SSEL(test_se), .CLK(
        CK), .Q(n7642), .QN(n5124) );
  sdffs1 \DFF_1182/Q_reg  ( .DIN(WX8302), .SDIN(n7640), .SSEL(test_se), .CLK(
        CK), .Q(n7641), .QN(n5125) );
  sdffs1 \DFF_1181/Q_reg  ( .DIN(WX8300), .SDIN(n7639), .SSEL(test_se), .CLK(
        CK), .Q(n7640), .QN(n5126) );
  sdffs1 \DFF_1180/Q_reg  ( .DIN(WX8298), .SDIN(n7638), .SSEL(test_se), .CLK(
        CK), .Q(n7639), .QN(n5127) );
  sdffs1 \DFF_1179/Q_reg  ( .DIN(WX8296), .SDIN(n7637), .SSEL(test_se), .CLK(
        CK), .Q(n7638), .QN(n5128) );
  sdffs1 \DFF_1178/Q_reg  ( .DIN(WX8294), .SDIN(n7636), .SSEL(test_se), .CLK(
        CK), .Q(n7637), .QN(n5129) );
  sdffs1 \DFF_1177/Q_reg  ( .DIN(WX8292), .SDIN(n7635), .SSEL(test_se), .CLK(
        CK), .Q(n7636), .QN(n5130) );
  sdffs1 \DFF_1176/Q_reg  ( .DIN(WX8290), .SDIN(n7634), .SSEL(test_se), .CLK(
        CK), .Q(n7635), .QN(n5131) );
  sdffs1 \DFF_1175/Q_reg  ( .DIN(WX8288), .SDIN(n7633), .SSEL(test_se), .CLK(
        CK), .Q(n7634), .QN(n5132) );
  sdffs1 \DFF_1174/Q_reg  ( .DIN(WX8286), .SDIN(n7632), .SSEL(test_se), .CLK(
        CK), .Q(n7633), .QN(n5133) );
  sdffs1 \DFF_1173/Q_reg  ( .DIN(WX8284), .SDIN(n7631), .SSEL(test_se), .CLK(
        CK), .Q(n7632), .QN(n5134) );
  sdffs1 \DFF_1172/Q_reg  ( .DIN(WX8282), .SDIN(n7630), .SSEL(test_se), .CLK(
        CK), .Q(n7631), .QN(n5135) );
  sdffs1 \DFF_1171/Q_reg  ( .DIN(WX8280), .SDIN(n7629), .SSEL(test_se), .CLK(
        CK), .Q(n7630), .QN(n5136) );
  sdffs1 \DFF_1170/Q_reg  ( .DIN(WX8278), .SDIN(n7628), .SSEL(test_se), .CLK(
        CK), .Q(n7629), .QN(n5137) );
  sdffs1 \DFF_1169/Q_reg  ( .DIN(WX8276), .SDIN(n7627), .SSEL(test_se), .CLK(
        CK), .Q(n7628), .QN(n5138) );
  sdffs1 \DFF_1168/Q_reg  ( .DIN(WX8274), .SDIN(n7626), .SSEL(test_se), .CLK(
        CK), .Q(n7627), .QN(n5139) );
  sdffs1 \DFF_1167/Q_reg  ( .DIN(WX8272), .SDIN(n7625), .SSEL(test_se), .CLK(
        CK), .Q(n7626), .QN(n5140) );
  sdffs1 \DFF_1166/Q_reg  ( .DIN(WX8270), .SDIN(n7624), .SSEL(test_se), .CLK(
        CK), .Q(n7625), .QN(n5141) );
  sdffs1 \DFF_1165/Q_reg  ( .DIN(WX8268), .SDIN(n7623), .SSEL(test_se), .CLK(
        CK), .Q(n7624), .QN(n5142) );
  sdffs1 \DFF_1164/Q_reg  ( .DIN(WX8266), .SDIN(n7622), .SSEL(test_se), .CLK(
        CK), .Q(n7623), .QN(n5143) );
  sdffs1 \DFF_1163/Q_reg  ( .DIN(WX8264), .SDIN(n7621), .SSEL(test_se), .CLK(
        CK), .Q(n7622), .QN(n5144) );
  sdffs1 \DFF_1162/Q_reg  ( .DIN(WX8262), .SDIN(n7620), .SSEL(test_se), .CLK(
        CK), .Q(n7621), .QN(n5145) );
  sdffs1 \DFF_1161/Q_reg  ( .DIN(WX8260), .SDIN(n7619), .SSEL(test_se), .CLK(
        CK), .Q(n7620), .QN(n5146) );
  sdffs1 \DFF_1160/Q_reg  ( .DIN(WX8258), .SDIN(n7618), .SSEL(test_se), .CLK(
        CK), .Q(n7619), .QN(n5147) );
  sdffs1 \DFF_1159/Q_reg  ( .DIN(WX8256), .SDIN(n7617), .SSEL(test_se), .CLK(
        CK), .Q(n7618), .QN(n5148) );
  sdffs1 \DFF_1158/Q_reg  ( .DIN(WX8254), .SDIN(n7616), .SSEL(test_se), .CLK(
        CK), .Q(n7617), .QN(n5149) );
  sdffs1 \DFF_1157/Q_reg  ( .DIN(WX8252), .SDIN(n7615), .SSEL(test_se), .CLK(
        CK), .Q(n7616), .QN(n5150) );
  sdffs1 \DFF_1156/Q_reg  ( .DIN(WX8250), .SDIN(n7614), .SSEL(test_se), .CLK(
        CK), .Q(n7615), .QN(n5151) );
  sdffs1 \DFF_1155/Q_reg  ( .DIN(WX8248), .SDIN(n7613), .SSEL(test_se), .CLK(
        CK), .Q(n7614), .QN(n5152) );
  sdffs1 \DFF_1154/Q_reg  ( .DIN(WX8246), .SDIN(n7612), .SSEL(test_se), .CLK(
        CK), .Q(n7613), .QN(n5153) );
  sdffs1 \DFF_1153/Q_reg  ( .DIN(WX8244), .SDIN(n7611), .SSEL(test_se), .CLK(
        CK), .Q(n7612), .QN(n5154) );
  sdffs1 \DFF_1152/Q_reg  ( .DIN(WX8242), .SDIN(CRC_OUT_4_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7611), .QN(n5123) );
  sdffs1 \DFF_1151/Q_reg  ( .DIN(WX7791), .SDIN(CRC_OUT_4_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_31), .QN(n5298) );
  sdffs1 \DFF_1150/Q_reg  ( .DIN(WX7789), .SDIN(CRC_OUT_4_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_30), .QN(n5293) );
  sdffs1 \DFF_1149/Q_reg  ( .DIN(WX7787), .SDIN(CRC_OUT_4_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_29), .QN(n5288) );
  sdffs1 \DFF_1148/Q_reg  ( .DIN(WX7785), .SDIN(CRC_OUT_4_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_28), .QN(n5283) );
  sdffs1 \DFF_1147/Q_reg  ( .DIN(WX7783), .SDIN(CRC_OUT_4_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_27), .QN(n5278) );
  sdffs1 \DFF_1146/Q_reg  ( .DIN(WX7781), .SDIN(CRC_OUT_4_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_26), .QN(n5273) );
  sdffs1 \DFF_1145/Q_reg  ( .DIN(WX7779), .SDIN(CRC_OUT_4_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_25), .QN(n5268) );
  sdffs1 \DFF_1144/Q_reg  ( .DIN(WX7777), .SDIN(CRC_OUT_4_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_24), .QN(n5263) );
  sdffs1 \DFF_1143/Q_reg  ( .DIN(WX7775), .SDIN(CRC_OUT_4_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_23), .QN(n5258) );
  sdffs1 \DFF_1142/Q_reg  ( .DIN(WX7773), .SDIN(CRC_OUT_4_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_22), .QN(n5253) );
  sdffs1 \DFF_1141/Q_reg  ( .DIN(WX7771), .SDIN(CRC_OUT_4_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_21), .QN(n5248) );
  sdffs1 \DFF_1140/Q_reg  ( .DIN(WX7769), .SDIN(CRC_OUT_4_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_20), .QN(n5243) );
  sdffs1 \DFF_1139/Q_reg  ( .DIN(WX7767), .SDIN(CRC_OUT_4_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_19), .QN(n5238) );
  sdffs1 \DFF_1138/Q_reg  ( .DIN(WX7765), .SDIN(CRC_OUT_4_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_18), .QN(n5233) );
  sdffs1 \DFF_1137/Q_reg  ( .DIN(WX7763), .SDIN(CRC_OUT_4_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_17), .QN(n5228) );
  sdffs1 \DFF_1136/Q_reg  ( .DIN(WX7761), .SDIN(CRC_OUT_4_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_16), .QN(n5223) );
  sdffs1 \DFF_1135/Q_reg  ( .DIN(WX7759), .SDIN(CRC_OUT_4_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_15), .QN(n5218) );
  sdffs1 \DFF_1134/Q_reg  ( .DIN(WX7757), .SDIN(CRC_OUT_4_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_14), .QN(n5214) );
  sdffs1 \DFF_1133/Q_reg  ( .DIN(WX7755), .SDIN(CRC_OUT_4_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_13), .QN(n5210) );
  sdffs1 \DFF_1132/Q_reg  ( .DIN(WX7753), .SDIN(CRC_OUT_4_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_12), .QN(n5206) );
  sdffs1 \DFF_1131/Q_reg  ( .DIN(WX7751), .SDIN(CRC_OUT_4_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_11), .QN(n5202) );
  sdffs1 \DFF_1130/Q_reg  ( .DIN(WX7749), .SDIN(CRC_OUT_4_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_10), .QN(n5198) );
  sdffs1 \DFF_1129/Q_reg  ( .DIN(WX7747), .SDIN(CRC_OUT_4_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_9), .QN(n5194) );
  sdffs1 \DFF_1128/Q_reg  ( .DIN(WX7745), .SDIN(CRC_OUT_4_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_8), .QN(n5190) );
  sdffs1 \DFF_1127/Q_reg  ( .DIN(WX7743), .SDIN(CRC_OUT_4_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_7), .QN(n5186) );
  sdffs1 \DFF_1126/Q_reg  ( .DIN(WX7741), .SDIN(CRC_OUT_4_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_6), .QN(n5182) );
  sdffs1 \DFF_1125/Q_reg  ( .DIN(WX7739), .SDIN(CRC_OUT_4_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_5), .QN(n5178) );
  sdffs1 \DFF_1124/Q_reg  ( .DIN(WX7737), .SDIN(CRC_OUT_4_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_4), .QN(n5174) );
  sdffs1 \DFF_1123/Q_reg  ( .DIN(WX7735), .SDIN(CRC_OUT_4_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_3), .QN(n5170) );
  sdffs1 \DFF_1122/Q_reg  ( .DIN(WX7733), .SDIN(CRC_OUT_4_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_2), .QN(n5166) );
  sdffs1 \DFF_1121/Q_reg  ( .DIN(WX7731), .SDIN(CRC_OUT_4_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_4_1), .QN(n5162) );
  sdffs1 \DFF_1120/Q_reg  ( .DIN(WX7729), .SDIN(n7610), .SSEL(test_se), .CLK(
        CK), .Q(CRC_OUT_4_0), .QN(n5158) );
  sdffs1 \DFF_1119/Q_reg  ( .DIN(WX7363), .SDIN(n7609), .SSEL(test_se), .CLK(
        CK), .Q(n7610), .QN(n3237) );
  sdffs1 \DFF_1118/Q_reg  ( .DIN(WX7361), .SDIN(n7608), .SSEL(test_se), .CLK(
        CK), .Q(n7609), .QN(n3238) );
  sdffs1 \DFF_1117/Q_reg  ( .DIN(WX7359), .SDIN(n7607), .SSEL(test_se), .CLK(
        CK), .Q(n7608), .QN(n3239) );
  sdffs1 \DFF_1116/Q_reg  ( .DIN(WX7357), .SDIN(n7606), .SSEL(test_se), .CLK(
        CK), .Q(n7607), .QN(n3240) );
  sdffs1 \DFF_1115/Q_reg  ( .DIN(WX7355), .SDIN(n7605), .SSEL(test_se), .CLK(
        CK), .Q(n7606), .QN(n3241) );
  sdffs1 \DFF_1114/Q_reg  ( .DIN(WX7353), .SDIN(n7604), .SSEL(test_se), .CLK(
        CK), .Q(n7605), .QN(n3242) );
  sdffs1 \DFF_1113/Q_reg  ( .DIN(WX7351), .SDIN(n7603), .SSEL(test_se), .CLK(
        CK), .Q(n7604), .QN(n3243) );
  sdffs1 \DFF_1112/Q_reg  ( .DIN(WX7349), .SDIN(n7602), .SSEL(test_se), .CLK(
        CK), .Q(n7603), .QN(n3244) );
  sdffs1 \DFF_1111/Q_reg  ( .DIN(WX7347), .SDIN(n7601), .SSEL(test_se), .CLK(
        CK), .Q(n7602), .QN(n3245) );
  sdffs1 \DFF_1110/Q_reg  ( .DIN(WX7345), .SDIN(n7600), .SSEL(test_se), .CLK(
        CK), .Q(n7601), .QN(n3246) );
  sdffs1 \DFF_1109/Q_reg  ( .DIN(WX7343), .SDIN(n7599), .SSEL(test_se), .CLK(
        CK), .Q(n7600), .QN(n3247) );
  sdffs1 \DFF_1108/Q_reg  ( .DIN(WX7341), .SDIN(n7598), .SSEL(test_se), .CLK(
        CK), .Q(n7599), .QN(n3248) );
  sdffs1 \DFF_1107/Q_reg  ( .DIN(WX7339), .SDIN(n7597), .SSEL(test_se), .CLK(
        CK), .Q(n7598), .QN(n3249) );
  sdffs1 \DFF_1106/Q_reg  ( .DIN(WX7337), .SDIN(n7596), .SSEL(test_se), .CLK(
        CK), .Q(n7597), .QN(n3250) );
  sdffs1 \DFF_1105/Q_reg  ( .DIN(WX7335), .SDIN(n7595), .SSEL(test_se), .CLK(
        CK), .Q(n7596), .QN(n3251) );
  sdffs1 \DFF_1104/Q_reg  ( .DIN(WX7333), .SDIN(n7594), .SSEL(test_se), .CLK(
        CK), .Q(n7595), .QN(n3252) );
  sdffs1 \DFF_1103/Q_reg  ( .DIN(WX7331), .SDIN(n7593), .SSEL(test_se), .CLK(
        CK), .Q(n7594), .QN(n5398) );
  sdffs1 \DFF_1102/Q_reg  ( .DIN(WX7329), .SDIN(n7592), .SSEL(test_se), .CLK(
        CK), .Q(n7593), .QN(n5403) );
  sdffs1 \DFF_1101/Q_reg  ( .DIN(WX7327), .SDIN(n7591), .SSEL(test_se), .CLK(
        CK), .Q(n7592), .QN(n5408) );
  sdffs1 \DFF_1100/Q_reg  ( .DIN(WX7325), .SDIN(n7590), .SSEL(test_se), .CLK(
        CK), .Q(n7591), .QN(n5413) );
  sdffs1 \DFF_1099/Q_reg  ( .DIN(WX7323), .SDIN(n7589), .SSEL(test_se), .CLK(
        CK), .Q(n7590), .QN(n5418) );
  sdffs1 \DFF_1098/Q_reg  ( .DIN(WX7321), .SDIN(n7588), .SSEL(test_se), .CLK(
        CK), .Q(n7589), .QN(n5423) );
  sdffs1 \DFF_1097/Q_reg  ( .DIN(WX7319), .SDIN(n7587), .SSEL(test_se), .CLK(
        CK), .Q(n7588), .QN(n5428) );
  sdffs1 \DFF_1096/Q_reg  ( .DIN(WX7317), .SDIN(n7586), .SSEL(test_se), .CLK(
        CK), .Q(n7587), .QN(n5433) );
  sdffs1 \DFF_1095/Q_reg  ( .DIN(WX7315), .SDIN(n7585), .SSEL(test_se), .CLK(
        CK), .Q(n7586), .QN(n5438) );
  sdffs1 \DFF_1094/Q_reg  ( .DIN(WX7313), .SDIN(n7584), .SSEL(test_se), .CLK(
        CK), .Q(n7585), .QN(n5443) );
  sdffs1 \DFF_1093/Q_reg  ( .DIN(WX7311), .SDIN(n7583), .SSEL(test_se), .CLK(
        CK), .Q(n7584), .QN(n5448) );
  sdffs1 \DFF_1092/Q_reg  ( .DIN(WX7309), .SDIN(n7582), .SSEL(test_se), .CLK(
        CK), .Q(n7583), .QN(n5453) );
  sdffs1 \DFF_1091/Q_reg  ( .DIN(WX7307), .SDIN(n7581), .SSEL(test_se), .CLK(
        CK), .Q(n7582), .QN(n5458) );
  sdffs1 \DFF_1090/Q_reg  ( .DIN(WX7305), .SDIN(n7580), .SSEL(test_se), .CLK(
        CK), .Q(n7581), .QN(n5463) );
  sdffs1 \DFF_1089/Q_reg  ( .DIN(WX7303), .SDIN(n7579), .SSEL(test_se), .CLK(
        CK), .Q(n7580), .QN(n5468) );
  sdffs1 \DFF_1088/Q_reg  ( .DIN(WX7301), .SDIN(n7578), .SSEL(test_se), .CLK(
        CK), .Q(n7579), .QN(n5473) );
  sdffs1 \DFF_1087/Q_reg  ( .DIN(WX7299), .SDIN(n7577), .SSEL(test_se), .CLK(
        CK), .Q(n7578), .QN(n5333) );
  sdffs1 \DFF_1086/Q_reg  ( .DIN(WX7297), .SDIN(n7576), .SSEL(test_se), .CLK(
        CK), .Q(n7577), .QN(n5337) );
  sdffs1 \DFF_1085/Q_reg  ( .DIN(WX7295), .SDIN(n7575), .SSEL(test_se), .CLK(
        CK), .Q(n7576), .QN(n5341) );
  sdffs1 \DFF_1084/Q_reg  ( .DIN(WX7293), .SDIN(n7574), .SSEL(test_se), .CLK(
        CK), .Q(n7575), .QN(n5345) );
  sdffs1 \DFF_1083/Q_reg  ( .DIN(WX7291), .SDIN(n7573), .SSEL(test_se), .CLK(
        CK), .Q(n7574), .QN(n5349) );
  sdffs1 \DFF_1082/Q_reg  ( .DIN(WX7289), .SDIN(n7572), .SSEL(test_se), .CLK(
        CK), .Q(n7573), .QN(n5353) );
  sdffs1 \DFF_1081/Q_reg  ( .DIN(WX7287), .SDIN(n7571), .SSEL(test_se), .CLK(
        CK), .Q(n7572), .QN(n5357) );
  sdffs1 \DFF_1080/Q_reg  ( .DIN(WX7285), .SDIN(n7570), .SSEL(test_se), .CLK(
        CK), .Q(n7571), .QN(n5361) );
  sdffs1 \DFF_1079/Q_reg  ( .DIN(WX7283), .SDIN(n7569), .SSEL(test_se), .CLK(
        CK), .Q(n7570), .QN(n5365) );
  sdffs1 \DFF_1078/Q_reg  ( .DIN(WX7281), .SDIN(n7568), .SSEL(test_se), .CLK(
        CK), .Q(n7569), .QN(n5369) );
  sdffs1 \DFF_1077/Q_reg  ( .DIN(WX7279), .SDIN(n7567), .SSEL(test_se), .CLK(
        CK), .Q(n7568), .QN(n5373) );
  sdffs1 \DFF_1076/Q_reg  ( .DIN(WX7277), .SDIN(n7566), .SSEL(test_se), .CLK(
        CK), .Q(n7567), .QN(n5377) );
  sdffs1 \DFF_1075/Q_reg  ( .DIN(WX7275), .SDIN(n7565), .SSEL(test_se), .CLK(
        CK), .Q(n7566), .QN(n5381) );
  sdffs1 \DFF_1074/Q_reg  ( .DIN(WX7273), .SDIN(n7564), .SSEL(test_se), .CLK(
        CK), .Q(n7565), .QN(n5385) );
  sdffs1 \DFF_1073/Q_reg  ( .DIN(WX7271), .SDIN(n7563), .SSEL(test_se), .CLK(
        CK), .Q(n7564), .QN(n5389) );
  sdffs1 \DFF_1072/Q_reg  ( .DIN(WX7269), .SDIN(n7562), .SSEL(test_se), .CLK(
        CK), .Q(n7563), .QN(n5393) );
  sdffs1 \DFF_1071/Q_reg  ( .DIN(WX7267), .SDIN(n7561), .SSEL(test_se), .CLK(
        CK), .Q(n7562), .QN(n5397) );
  sdffs1 \DFF_1070/Q_reg  ( .DIN(WX7265), .SDIN(n7560), .SSEL(test_se), .CLK(
        CK), .Q(n7561), .QN(n5402) );
  sdffs1 \DFF_1069/Q_reg  ( .DIN(WX7263), .SDIN(n7559), .SSEL(test_se), .CLK(
        CK), .Q(n7560), .QN(n5407) );
  sdffs1 \DFF_1068/Q_reg  ( .DIN(WX7261), .SDIN(n7558), .SSEL(test_se), .CLK(
        CK), .Q(n7559), .QN(n5412) );
  sdffs1 \DFF_1067/Q_reg  ( .DIN(WX7259), .SDIN(n7557), .SSEL(test_se), .CLK(
        CK), .Q(n7558), .QN(n5417) );
  sdffs1 \DFF_1066/Q_reg  ( .DIN(WX7257), .SDIN(n7556), .SSEL(test_se), .CLK(
        CK), .Q(n7557), .QN(n5422) );
  sdffs1 \DFF_1065/Q_reg  ( .DIN(WX7255), .SDIN(n7555), .SSEL(test_se), .CLK(
        CK), .Q(n7556), .QN(n5427) );
  sdffs1 \DFF_1064/Q_reg  ( .DIN(WX7253), .SDIN(n7554), .SSEL(test_se), .CLK(
        CK), .Q(n7555), .QN(n5432) );
  sdffs1 \DFF_1063/Q_reg  ( .DIN(WX7251), .SDIN(n7553), .SSEL(test_se), .CLK(
        CK), .Q(n7554), .QN(n5437) );
  sdffs1 \DFF_1062/Q_reg  ( .DIN(WX7249), .SDIN(n7552), .SSEL(test_se), .CLK(
        CK), .Q(n7553), .QN(n5442) );
  sdffs1 \DFF_1061/Q_reg  ( .DIN(WX7247), .SDIN(n7551), .SSEL(test_se), .CLK(
        CK), .Q(n7552), .QN(n5447) );
  sdffs1 \DFF_1060/Q_reg  ( .DIN(WX7245), .SDIN(n7550), .SSEL(test_se), .CLK(
        CK), .Q(n7551), .QN(n5452) );
  sdffs1 \DFF_1059/Q_reg  ( .DIN(WX7243), .SDIN(n7549), .SSEL(test_se), .CLK(
        CK), .Q(n7550), .QN(n5457) );
  sdffs1 \DFF_1058/Q_reg  ( .DIN(WX7241), .SDIN(n7548), .SSEL(test_se), .CLK(
        CK), .Q(n7549), .QN(n5462) );
  sdffs1 \DFF_1057/Q_reg  ( .DIN(WX7239), .SDIN(n7547), .SSEL(test_se), .CLK(
        CK), .Q(n7548), .QN(n5467) );
  sdffs1 \DFF_1056/Q_reg  ( .DIN(WX7237), .SDIN(n7546), .SSEL(test_se), .CLK(
        CK), .Q(n7547), .QN(n5472) );
  sdffs1 \DFF_1055/Q_reg  ( .DIN(WX7235), .SDIN(n7545), .SSEL(test_se), .CLK(
        CK), .Q(n7546), .QN(n5332) );
  sdffs1 \DFF_1054/Q_reg  ( .DIN(WX7233), .SDIN(n7544), .SSEL(test_se), .CLK(
        CK), .Q(n7545), .QN(n5336) );
  sdffs1 \DFF_1053/Q_reg  ( .DIN(WX7231), .SDIN(n7543), .SSEL(test_se), .CLK(
        CK), .Q(n7544), .QN(n5340) );
  sdffs1 \DFF_1052/Q_reg  ( .DIN(WX7229), .SDIN(n7542), .SSEL(test_se), .CLK(
        CK), .Q(n7543), .QN(n5344) );
  sdffs1 \DFF_1051/Q_reg  ( .DIN(WX7227), .SDIN(n7541), .SSEL(test_se), .CLK(
        CK), .Q(n7542), .QN(n5348) );
  sdffs1 \DFF_1050/Q_reg  ( .DIN(WX7225), .SDIN(n7540), .SSEL(test_se), .CLK(
        CK), .Q(n7541), .QN(n5352) );
  sdffs1 \DFF_1049/Q_reg  ( .DIN(WX7223), .SDIN(n7539), .SSEL(test_se), .CLK(
        CK), .Q(n7540), .QN(n5356) );
  sdffs1 \DFF_1048/Q_reg  ( .DIN(WX7221), .SDIN(n7538), .SSEL(test_se), .CLK(
        CK), .Q(n7539), .QN(n5360) );
  sdffs1 \DFF_1047/Q_reg  ( .DIN(WX7219), .SDIN(n7537), .SSEL(test_se), .CLK(
        CK), .Q(n7538), .QN(n5364) );
  sdffs1 \DFF_1046/Q_reg  ( .DIN(WX7217), .SDIN(n7536), .SSEL(test_se), .CLK(
        CK), .Q(n7537), .QN(n5368) );
  sdffs1 \DFF_1045/Q_reg  ( .DIN(WX7215), .SDIN(n7535), .SSEL(test_se), .CLK(
        CK), .Q(n7536), .QN(n5372) );
  sdffs1 \DFF_1044/Q_reg  ( .DIN(WX7213), .SDIN(n7534), .SSEL(test_se), .CLK(
        CK), .Q(n7535), .QN(n5376) );
  sdffs1 \DFF_1043/Q_reg  ( .DIN(WX7211), .SDIN(n7533), .SSEL(test_se), .CLK(
        CK), .Q(n7534), .QN(n5380) );
  sdffs1 \DFF_1042/Q_reg  ( .DIN(WX7209), .SDIN(n7532), .SSEL(test_se), .CLK(
        CK), .Q(n7533), .QN(n5384) );
  sdffs1 \DFF_1041/Q_reg  ( .DIN(WX7207), .SDIN(n7531), .SSEL(test_se), .CLK(
        CK), .Q(n7532), .QN(n5388) );
  sdffs1 \DFF_1040/Q_reg  ( .DIN(WX7205), .SDIN(n5396), .SSEL(test_se), .CLK(
        CK), .Q(n7531), .QN(n5392) );
  sdffs1 \DFF_1039/Q_reg  ( .DIN(WX7203), .SDIN(n5401), .SSEL(test_se), .CLK(
        CK), .Q(n5396) );
  sdffs1 \DFF_1038/Q_reg  ( .DIN(WX7201), .SDIN(n5406), .SSEL(test_se), .CLK(
        CK), .Q(n5401) );
  sdffs1 \DFF_1037/Q_reg  ( .DIN(WX7199), .SDIN(n5411), .SSEL(test_se), .CLK(
        CK), .Q(n5406) );
  sdffs1 \DFF_1036/Q_reg  ( .DIN(WX7197), .SDIN(n5416), .SSEL(test_se), .CLK(
        CK), .Q(n5411) );
  sdffs1 \DFF_1035/Q_reg  ( .DIN(WX7195), .SDIN(n5421), .SSEL(test_se), .CLK(
        CK), .Q(n5416) );
  sdffs1 \DFF_1034/Q_reg  ( .DIN(WX7193), .SDIN(n5426), .SSEL(test_se), .CLK(
        CK), .Q(n5421) );
  sdffs1 \DFF_1033/Q_reg  ( .DIN(WX7191), .SDIN(n5431), .SSEL(test_se), .CLK(
        CK), .Q(n5426) );
  sdffs1 \DFF_1032/Q_reg  ( .DIN(WX7189), .SDIN(n5436), .SSEL(test_se), .CLK(
        CK), .Q(n5431) );
  sdffs1 \DFF_1031/Q_reg  ( .DIN(WX7187), .SDIN(n5441), .SSEL(test_se), .CLK(
        CK), .Q(n5436) );
  sdffs1 \DFF_1030/Q_reg  ( .DIN(WX7185), .SDIN(n5446), .SSEL(test_se), .CLK(
        CK), .Q(n5441) );
  sdffs1 \DFF_1029/Q_reg  ( .DIN(WX7183), .SDIN(n5451), .SSEL(test_se), .CLK(
        CK), .Q(n5446) );
  sdffs1 \DFF_1028/Q_reg  ( .DIN(WX7181), .SDIN(n5456), .SSEL(test_se), .CLK(
        CK), .Q(n5451) );
  sdffs1 \DFF_1027/Q_reg  ( .DIN(WX7179), .SDIN(n5461), .SSEL(test_se), .CLK(
        CK), .Q(n5456) );
  sdffs1 \DFF_1026/Q_reg  ( .DIN(WX7177), .SDIN(n5466), .SSEL(test_se), .CLK(
        CK), .Q(n5461) );
  sdffs1 \DFF_1025/Q_reg  ( .DIN(WX7175), .SDIN(n5471), .SSEL(test_se), .CLK(
        CK), .Q(n5466) );
  sdffs1 \DFF_1024/Q_reg  ( .DIN(WX7173), .SDIN(n5331), .SSEL(test_se), .CLK(
        CK), .Q(n5471) );
  sdffs1 \DFF_1023/Q_reg  ( .DIN(WX7171), .SDIN(n5335), .SSEL(test_se), .CLK(
        CK), .Q(n5331) );
  sdffs1 \DFF_1022/Q_reg  ( .DIN(WX7169), .SDIN(n5339), .SSEL(test_se), .CLK(
        CK), .Q(n5335) );
  sdffs1 \DFF_1021/Q_reg  ( .DIN(WX7167), .SDIN(n5343), .SSEL(test_se), .CLK(
        CK), .Q(n5339) );
  sdffs1 \DFF_1020/Q_reg  ( .DIN(WX7165), .SDIN(n5347), .SSEL(test_se), .CLK(
        CK), .Q(n5343) );
  sdffs1 \DFF_1019/Q_reg  ( .DIN(WX7163), .SDIN(n5351), .SSEL(test_se), .CLK(
        CK), .Q(n5347) );
  sdffs1 \DFF_1018/Q_reg  ( .DIN(WX7161), .SDIN(n5355), .SSEL(test_se), .CLK(
        CK), .Q(n5351) );
  sdffs1 \DFF_1017/Q_reg  ( .DIN(WX7159), .SDIN(n5359), .SSEL(test_se), .CLK(
        CK), .Q(n5355) );
  sdffs1 \DFF_1016/Q_reg  ( .DIN(WX7157), .SDIN(n5363), .SSEL(test_se), .CLK(
        CK), .Q(n5359) );
  sdffs1 \DFF_1015/Q_reg  ( .DIN(WX7155), .SDIN(n5367), .SSEL(test_se), .CLK(
        CK), .Q(n5363) );
  sdffs1 \DFF_1014/Q_reg  ( .DIN(WX7153), .SDIN(n5371), .SSEL(test_se), .CLK(
        CK), .Q(n5367) );
  sdffs1 \DFF_1013/Q_reg  ( .DIN(WX7151), .SDIN(n5375), .SSEL(test_se), .CLK(
        CK), .Q(n5371) );
  sdffs1 \DFF_1012/Q_reg  ( .DIN(WX7149), .SDIN(n5379), .SSEL(test_se), .CLK(
        CK), .Q(n5375) );
  sdffs1 \DFF_1011/Q_reg  ( .DIN(WX7147), .SDIN(n5383), .SSEL(test_se), .CLK(
        CK), .Q(n5379) );
  sdffs1 \DFF_1010/Q_reg  ( .DIN(WX7145), .SDIN(n5387), .SSEL(test_se), .CLK(
        CK), .Q(n5383) );
  sdffs1 \DFF_1009/Q_reg  ( .DIN(WX7143), .SDIN(n5391), .SSEL(test_se), .CLK(
        CK), .Q(n5387) );
  sdffs1 \DFF_1008/Q_reg  ( .DIN(WX7141), .SDIN(n7530), .SSEL(test_se), .CLK(
        CK), .Q(n5391) );
  sdffs1 \DFF_1007/Q_reg  ( .DIN(WX7139), .SDIN(n7529), .SSEL(test_se), .CLK(
        CK), .Q(n7530), .QN(n5395) );
  sdffs1 \DFF_1006/Q_reg  ( .DIN(WX7137), .SDIN(n7528), .SSEL(test_se), .CLK(
        CK), .Q(n7529), .QN(n5400) );
  sdffs1 \DFF_1005/Q_reg  ( .DIN(WX7135), .SDIN(n7527), .SSEL(test_se), .CLK(
        CK), .Q(n7528), .QN(n5405) );
  sdffs1 \DFF_1004/Q_reg  ( .DIN(WX7133), .SDIN(n7526), .SSEL(test_se), .CLK(
        CK), .Q(n7527), .QN(n5410) );
  sdffs1 \DFF_1003/Q_reg  ( .DIN(WX7131), .SDIN(n7525), .SSEL(test_se), .CLK(
        CK), .Q(n7526), .QN(n5415) );
  sdffs1 \DFF_1002/Q_reg  ( .DIN(WX7129), .SDIN(n7524), .SSEL(test_se), .CLK(
        CK), .Q(n7525), .QN(n5420) );
  sdffs1 \DFF_1001/Q_reg  ( .DIN(WX7127), .SDIN(n7523), .SSEL(test_se), .CLK(
        CK), .Q(n7524), .QN(n5425) );
  sdffs1 \DFF_1000/Q_reg  ( .DIN(WX7125), .SDIN(n7522), .SSEL(test_se), .CLK(
        CK), .Q(n7523), .QN(n5430) );
  sdffs1 \DFF_999/Q_reg  ( .DIN(WX7123), .SDIN(n7521), .SSEL(test_se), .CLK(CK), .Q(n7522), .QN(n5435) );
  sdffs1 \DFF_998/Q_reg  ( .DIN(WX7121), .SDIN(n7520), .SSEL(test_se), .CLK(CK), .Q(n7521), .QN(n5440) );
  sdffs1 \DFF_997/Q_reg  ( .DIN(WX7119), .SDIN(n7519), .SSEL(test_se), .CLK(CK), .Q(n7520), .QN(n5445) );
  sdffs1 \DFF_996/Q_reg  ( .DIN(WX7117), .SDIN(n7518), .SSEL(test_se), .CLK(CK), .Q(n7519), .QN(n5450) );
  sdffs1 \DFF_995/Q_reg  ( .DIN(WX7115), .SDIN(n7517), .SSEL(test_se), .CLK(CK), .Q(n7518), .QN(n5455) );
  sdffs1 \DFF_994/Q_reg  ( .DIN(WX7113), .SDIN(n7516), .SSEL(test_se), .CLK(CK), .Q(n7517), .QN(n5460) );
  sdffs1 \DFF_993/Q_reg  ( .DIN(WX7111), .SDIN(n7515), .SSEL(test_se), .CLK(CK), .Q(n7516), .QN(n5465) );
  sdffs1 \DFF_992/Q_reg  ( .DIN(WX7109), .SDIN(n7514), .SSEL(test_se), .CLK(CK), .Q(n7515), .QN(n5470) );
  sdffs1 \DFF_991/Q_reg  ( .DIN(WX7011), .SDIN(n7513), .SSEL(test_se), .CLK(CK), .Q(n7514), .QN(n5300) );
  sdffs1 \DFF_990/Q_reg  ( .DIN(WX7009), .SDIN(n7512), .SSEL(test_se), .CLK(CK), .Q(n7513), .QN(n5301) );
  sdffs1 \DFF_989/Q_reg  ( .DIN(WX7007), .SDIN(n7511), .SSEL(test_se), .CLK(CK), .Q(n7512), .QN(n5302) );
  sdffs1 \DFF_988/Q_reg  ( .DIN(WX7005), .SDIN(n7510), .SSEL(test_se), .CLK(CK), .Q(n7511), .QN(n5303) );
  sdffs1 \DFF_987/Q_reg  ( .DIN(WX7003), .SDIN(n7509), .SSEL(test_se), .CLK(CK), .Q(n7510), .QN(n5304) );
  sdffs1 \DFF_986/Q_reg  ( .DIN(WX7001), .SDIN(n7508), .SSEL(test_se), .CLK(CK), .Q(n7509), .QN(n5305) );
  sdffs1 \DFF_985/Q_reg  ( .DIN(WX6999), .SDIN(n7507), .SSEL(test_se), .CLK(CK), .Q(n7508), .QN(n5306) );
  sdffs1 \DFF_984/Q_reg  ( .DIN(WX6997), .SDIN(n7506), .SSEL(test_se), .CLK(CK), .Q(n7507), .QN(n5307) );
  sdffs1 \DFF_983/Q_reg  ( .DIN(WX6995), .SDIN(n7505), .SSEL(test_se), .CLK(CK), .Q(n7506), .QN(n5308) );
  sdffs1 \DFF_982/Q_reg  ( .DIN(WX6993), .SDIN(n7504), .SSEL(test_se), .CLK(CK), .Q(n7505), .QN(n5309) );
  sdffs1 \DFF_981/Q_reg  ( .DIN(WX6991), .SDIN(n7503), .SSEL(test_se), .CLK(CK), .Q(n7504), .QN(n5310) );
  sdffs1 \DFF_980/Q_reg  ( .DIN(WX6989), .SDIN(n7502), .SSEL(test_se), .CLK(CK), .Q(n7503), .QN(n5311) );
  sdffs1 \DFF_979/Q_reg  ( .DIN(WX6987), .SDIN(n7501), .SSEL(test_se), .CLK(CK), .Q(n7502), .QN(n5312) );
  sdffs1 \DFF_978/Q_reg  ( .DIN(WX6985), .SDIN(n7500), .SSEL(test_se), .CLK(CK), .Q(n7501), .QN(n5313) );
  sdffs1 \DFF_977/Q_reg  ( .DIN(WX6983), .SDIN(n7499), .SSEL(test_se), .CLK(CK), .Q(n7500), .QN(n5314) );
  sdffs1 \DFF_976/Q_reg  ( .DIN(WX6981), .SDIN(n7498), .SSEL(test_se), .CLK(CK), .Q(n7499), .QN(n5315) );
  sdffs1 \DFF_975/Q_reg  ( .DIN(WX6979), .SDIN(n7497), .SSEL(test_se), .CLK(CK), .Q(n7498), .QN(n5316) );
  sdffs1 \DFF_974/Q_reg  ( .DIN(WX6977), .SDIN(n7496), .SSEL(test_se), .CLK(CK), .Q(n7497), .QN(n5317) );
  sdffs1 \DFF_973/Q_reg  ( .DIN(WX6975), .SDIN(n7495), .SSEL(test_se), .CLK(CK), .Q(n7496), .QN(n5318) );
  sdffs1 \DFF_972/Q_reg  ( .DIN(WX6973), .SDIN(n7494), .SSEL(test_se), .CLK(CK), .Q(n7495), .QN(n5319) );
  sdffs1 \DFF_971/Q_reg  ( .DIN(WX6971), .SDIN(n7493), .SSEL(test_se), .CLK(CK), .Q(n7494), .QN(n5320) );
  sdffs1 \DFF_970/Q_reg  ( .DIN(WX6969), .SDIN(n7492), .SSEL(test_se), .CLK(CK), .Q(n7493), .QN(n5321) );
  sdffs1 \DFF_969/Q_reg  ( .DIN(WX6967), .SDIN(n7491), .SSEL(test_se), .CLK(CK), .Q(n7492), .QN(n5322) );
  sdffs1 \DFF_968/Q_reg  ( .DIN(WX6965), .SDIN(n7490), .SSEL(test_se), .CLK(CK), .Q(n7491), .QN(n5323) );
  sdffs1 \DFF_967/Q_reg  ( .DIN(WX6963), .SDIN(n7489), .SSEL(test_se), .CLK(CK), .Q(n7490), .QN(n5324) );
  sdffs1 \DFF_966/Q_reg  ( .DIN(WX6961), .SDIN(n7488), .SSEL(test_se), .CLK(CK), .Q(n7489), .QN(n5325) );
  sdffs1 \DFF_965/Q_reg  ( .DIN(WX6959), .SDIN(n7487), .SSEL(test_se), .CLK(CK), .Q(n7488), .QN(n5326) );
  sdffs1 \DFF_964/Q_reg  ( .DIN(WX6957), .SDIN(n7486), .SSEL(test_se), .CLK(CK), .Q(n7487), .QN(n5327) );
  sdffs1 \DFF_963/Q_reg  ( .DIN(WX6955), .SDIN(n7485), .SSEL(test_se), .CLK(CK), .Q(n7486), .QN(n5328) );
  sdffs1 \DFF_962/Q_reg  ( .DIN(WX6953), .SDIN(n7484), .SSEL(test_se), .CLK(CK), .Q(n7485), .QN(n5329) );
  sdffs1 \DFF_961/Q_reg  ( .DIN(WX6951), .SDIN(n7483), .SSEL(test_se), .CLK(CK), .Q(n7484), .QN(n5330) );
  sdffs1 \DFF_960/Q_reg  ( .DIN(WX6949), .SDIN(CRC_OUT_5_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7483), .QN(n5299) );
  sdffs1 \DFF_959/Q_reg  ( .DIN(WX6498), .SDIN(CRC_OUT_5_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_31), .QN(n5474) );
  sdffs1 \DFF_958/Q_reg  ( .DIN(WX6496), .SDIN(CRC_OUT_5_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_30), .QN(n5469) );
  sdffs1 \DFF_957/Q_reg  ( .DIN(WX6494), .SDIN(CRC_OUT_5_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_29), .QN(n5464) );
  sdffs1 \DFF_956/Q_reg  ( .DIN(WX6492), .SDIN(CRC_OUT_5_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_28), .QN(n5459) );
  sdffs1 \DFF_955/Q_reg  ( .DIN(WX6490), .SDIN(CRC_OUT_5_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_27), .QN(n5454) );
  sdffs1 \DFF_954/Q_reg  ( .DIN(WX6488), .SDIN(CRC_OUT_5_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_26), .QN(n5449) );
  sdffs1 \DFF_953/Q_reg  ( .DIN(WX6486), .SDIN(CRC_OUT_5_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_25), .QN(n5444) );
  sdffs1 \DFF_952/Q_reg  ( .DIN(WX6484), .SDIN(CRC_OUT_5_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_24), .QN(n5439) );
  sdffs1 \DFF_951/Q_reg  ( .DIN(WX6482), .SDIN(CRC_OUT_5_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_23), .QN(n5434) );
  sdffs1 \DFF_950/Q_reg  ( .DIN(WX6480), .SDIN(CRC_OUT_5_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_22), .QN(n5429) );
  sdffs1 \DFF_949/Q_reg  ( .DIN(WX6478), .SDIN(CRC_OUT_5_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_21), .QN(n5424) );
  sdffs1 \DFF_948/Q_reg  ( .DIN(WX6476), .SDIN(CRC_OUT_5_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_20), .QN(n5419) );
  sdffs1 \DFF_947/Q_reg  ( .DIN(WX6474), .SDIN(CRC_OUT_5_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_19), .QN(n5414) );
  sdffs1 \DFF_946/Q_reg  ( .DIN(WX6472), .SDIN(CRC_OUT_5_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_18), .QN(n5409) );
  sdffs1 \DFF_945/Q_reg  ( .DIN(WX6470), .SDIN(CRC_OUT_5_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_17), .QN(n5404) );
  sdffs1 \DFF_944/Q_reg  ( .DIN(WX6468), .SDIN(CRC_OUT_5_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_16), .QN(n5399) );
  sdffs1 \DFF_943/Q_reg  ( .DIN(WX6466), .SDIN(CRC_OUT_5_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_15), .QN(n5394) );
  sdffs1 \DFF_942/Q_reg  ( .DIN(WX6464), .SDIN(CRC_OUT_5_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_14), .QN(n5390) );
  sdffs1 \DFF_941/Q_reg  ( .DIN(WX6462), .SDIN(CRC_OUT_5_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_13), .QN(n5386) );
  sdffs1 \DFF_940/Q_reg  ( .DIN(WX6460), .SDIN(CRC_OUT_5_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_12), .QN(n5382) );
  sdffs1 \DFF_939/Q_reg  ( .DIN(WX6458), .SDIN(CRC_OUT_5_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_11), .QN(n5378) );
  sdffs1 \DFF_938/Q_reg  ( .DIN(WX6456), .SDIN(CRC_OUT_5_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_10), .QN(n5374) );
  sdffs1 \DFF_937/Q_reg  ( .DIN(WX6454), .SDIN(CRC_OUT_5_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_9), .QN(n5370) );
  sdffs1 \DFF_936/Q_reg  ( .DIN(WX6452), .SDIN(CRC_OUT_5_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_8), .QN(n5366) );
  sdffs1 \DFF_935/Q_reg  ( .DIN(WX6450), .SDIN(CRC_OUT_5_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_7), .QN(n5362) );
  sdffs1 \DFF_934/Q_reg  ( .DIN(WX6448), .SDIN(CRC_OUT_5_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_6), .QN(n5358) );
  sdffs1 \DFF_933/Q_reg  ( .DIN(WX6446), .SDIN(CRC_OUT_5_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_5), .QN(n5354) );
  sdffs1 \DFF_932/Q_reg  ( .DIN(WX6444), .SDIN(CRC_OUT_5_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_4), .QN(n5350) );
  sdffs1 \DFF_931/Q_reg  ( .DIN(WX6442), .SDIN(CRC_OUT_5_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_3), .QN(n5346) );
  sdffs1 \DFF_930/Q_reg  ( .DIN(WX6440), .SDIN(CRC_OUT_5_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_2), .QN(n5342) );
  sdffs1 \DFF_929/Q_reg  ( .DIN(WX6438), .SDIN(CRC_OUT_5_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_5_1), .QN(n5338) );
  sdffs1 \DFF_928/Q_reg  ( .DIN(WX6436), .SDIN(n7482), .SSEL(test_se), .CLK(CK), .Q(CRC_OUT_5_0), .QN(n5334) );
  sdffs1 \DFF_927/Q_reg  ( .DIN(WX6070), .SDIN(n7481), .SSEL(test_se), .CLK(CK), .Q(n7482), .QN(n3253) );
  sdffs1 \DFF_926/Q_reg  ( .DIN(WX6068), .SDIN(n7480), .SSEL(test_se), .CLK(CK), .Q(n7481), .QN(n3254) );
  sdffs1 \DFF_925/Q_reg  ( .DIN(WX6066), .SDIN(n7479), .SSEL(test_se), .CLK(CK), .Q(n7480), .QN(n3255) );
  sdffs1 \DFF_924/Q_reg  ( .DIN(WX6064), .SDIN(n7478), .SSEL(test_se), .CLK(CK), .Q(n7479), .QN(n3256) );
  sdffs1 \DFF_923/Q_reg  ( .DIN(WX6062), .SDIN(n7477), .SSEL(test_se), .CLK(CK), .Q(n7478), .QN(n3257) );
  sdffs1 \DFF_922/Q_reg  ( .DIN(WX6060), .SDIN(n7476), .SSEL(test_se), .CLK(CK), .Q(n7477), .QN(n3258) );
  sdffs1 \DFF_921/Q_reg  ( .DIN(WX6058), .SDIN(n7475), .SSEL(test_se), .CLK(CK), .Q(n7476), .QN(n3259) );
  sdffs1 \DFF_920/Q_reg  ( .DIN(WX6056), .SDIN(n7474), .SSEL(test_se), .CLK(CK), .Q(n7475), .QN(n3260) );
  sdffs1 \DFF_919/Q_reg  ( .DIN(WX6054), .SDIN(n7473), .SSEL(test_se), .CLK(CK), .Q(n7474), .QN(n3261) );
  sdffs1 \DFF_918/Q_reg  ( .DIN(WX6052), .SDIN(n7472), .SSEL(test_se), .CLK(CK), .Q(n7473), .QN(n3262) );
  sdffs1 \DFF_917/Q_reg  ( .DIN(WX6050), .SDIN(n7471), .SSEL(test_se), .CLK(CK), .Q(n7472), .QN(n3263) );
  sdffs1 \DFF_916/Q_reg  ( .DIN(WX6048), .SDIN(n7470), .SSEL(test_se), .CLK(CK), .Q(n7471), .QN(n3264) );
  sdffs1 \DFF_915/Q_reg  ( .DIN(WX6046), .SDIN(n7469), .SSEL(test_se), .CLK(CK), .Q(n7470), .QN(n3265) );
  sdffs1 \DFF_914/Q_reg  ( .DIN(WX6044), .SDIN(n7468), .SSEL(test_se), .CLK(CK), .Q(n7469), .QN(n3266) );
  sdffs1 \DFF_913/Q_reg  ( .DIN(WX6042), .SDIN(n7467), .SSEL(test_se), .CLK(CK), .Q(n7468), .QN(n3267) );
  sdffs1 \DFF_912/Q_reg  ( .DIN(WX6040), .SDIN(n7466), .SSEL(test_se), .CLK(CK), .Q(n7467), .QN(n3268) );
  sdffs1 \DFF_911/Q_reg  ( .DIN(WX6038), .SDIN(n7465), .SSEL(test_se), .CLK(CK), .Q(n7466), .QN(n5574) );
  sdffs1 \DFF_910/Q_reg  ( .DIN(WX6036), .SDIN(n7464), .SSEL(test_se), .CLK(CK), .Q(n7465), .QN(n5579) );
  sdffs1 \DFF_909/Q_reg  ( .DIN(WX6034), .SDIN(n7463), .SSEL(test_se), .CLK(CK), .Q(n7464), .QN(n5584) );
  sdffs1 \DFF_908/Q_reg  ( .DIN(WX6032), .SDIN(n7462), .SSEL(test_se), .CLK(CK), .Q(n7463), .QN(n5589) );
  sdffs1 \DFF_907/Q_reg  ( .DIN(WX6030), .SDIN(n7461), .SSEL(test_se), .CLK(CK), .Q(n7462), .QN(n5594) );
  sdffs1 \DFF_906/Q_reg  ( .DIN(WX6028), .SDIN(n7460), .SSEL(test_se), .CLK(CK), .Q(n7461), .QN(n5599) );
  sdffs1 \DFF_905/Q_reg  ( .DIN(WX6026), .SDIN(n7459), .SSEL(test_se), .CLK(CK), .Q(n7460), .QN(n5604) );
  sdffs1 \DFF_904/Q_reg  ( .DIN(WX6024), .SDIN(n7458), .SSEL(test_se), .CLK(CK), .Q(n7459), .QN(n5609) );
  sdffs1 \DFF_903/Q_reg  ( .DIN(WX6022), .SDIN(n7457), .SSEL(test_se), .CLK(CK), .Q(n7458), .QN(n5614) );
  sdffs1 \DFF_902/Q_reg  ( .DIN(WX6020), .SDIN(n7456), .SSEL(test_se), .CLK(CK), .Q(n7457), .QN(n5619) );
  sdffs1 \DFF_901/Q_reg  ( .DIN(WX6018), .SDIN(n7455), .SSEL(test_se), .CLK(CK), .Q(n7456), .QN(n5624) );
  sdffs1 \DFF_900/Q_reg  ( .DIN(WX6016), .SDIN(n7454), .SSEL(test_se), .CLK(CK), .Q(n7455), .QN(n5629) );
  sdffs1 \DFF_899/Q_reg  ( .DIN(WX6014), .SDIN(n7453), .SSEL(test_se), .CLK(CK), .Q(n7454), .QN(n5634) );
  sdffs1 \DFF_898/Q_reg  ( .DIN(WX6012), .SDIN(n7452), .SSEL(test_se), .CLK(CK), .Q(n7453), .QN(n5639) );
  sdffs1 \DFF_897/Q_reg  ( .DIN(WX6010), .SDIN(n7451), .SSEL(test_se), .CLK(CK), .Q(n7452), .QN(n5644) );
  sdffs1 \DFF_896/Q_reg  ( .DIN(WX6008), .SDIN(n7450), .SSEL(test_se), .CLK(CK), .Q(n7451), .QN(n5649) );
  sdffs1 \DFF_895/Q_reg  ( .DIN(WX6006), .SDIN(n7449), .SSEL(test_se), .CLK(CK), .Q(n7450), .QN(n5509) );
  sdffs1 \DFF_894/Q_reg  ( .DIN(WX6004), .SDIN(n7448), .SSEL(test_se), .CLK(CK), .Q(n7449), .QN(n5513) );
  sdffs1 \DFF_893/Q_reg  ( .DIN(WX6002), .SDIN(n7447), .SSEL(test_se), .CLK(CK), .Q(n7448), .QN(n5517) );
  sdffs1 \DFF_892/Q_reg  ( .DIN(WX6000), .SDIN(n7446), .SSEL(test_se), .CLK(CK), .Q(n7447), .QN(n5521) );
  sdffs1 \DFF_891/Q_reg  ( .DIN(WX5998), .SDIN(n7445), .SSEL(test_se), .CLK(CK), .Q(n7446), .QN(n5525) );
  sdffs1 \DFF_890/Q_reg  ( .DIN(WX5996), .SDIN(n7444), .SSEL(test_se), .CLK(CK), .Q(n7445), .QN(n5529) );
  sdffs1 \DFF_889/Q_reg  ( .DIN(WX5994), .SDIN(n7443), .SSEL(test_se), .CLK(CK), .Q(n7444), .QN(n5533) );
  sdffs1 \DFF_888/Q_reg  ( .DIN(WX5992), .SDIN(n7442), .SSEL(test_se), .CLK(CK), .Q(n7443), .QN(n5537) );
  sdffs1 \DFF_887/Q_reg  ( .DIN(WX5990), .SDIN(n7441), .SSEL(test_se), .CLK(CK), .Q(n7442), .QN(n5541) );
  sdffs1 \DFF_886/Q_reg  ( .DIN(WX5988), .SDIN(n7440), .SSEL(test_se), .CLK(CK), .Q(n7441), .QN(n5545) );
  sdffs1 \DFF_885/Q_reg  ( .DIN(WX5986), .SDIN(n7439), .SSEL(test_se), .CLK(CK), .Q(n7440), .QN(n5549) );
  sdffs1 \DFF_884/Q_reg  ( .DIN(WX5984), .SDIN(n7438), .SSEL(test_se), .CLK(CK), .Q(n7439), .QN(n5553) );
  sdffs1 \DFF_883/Q_reg  ( .DIN(WX5982), .SDIN(n7437), .SSEL(test_se), .CLK(CK), .Q(n7438), .QN(n5557) );
  sdffs1 \DFF_882/Q_reg  ( .DIN(WX5980), .SDIN(n7436), .SSEL(test_se), .CLK(CK), .Q(n7437), .QN(n5561) );
  sdffs1 \DFF_881/Q_reg  ( .DIN(WX5978), .SDIN(n7435), .SSEL(test_se), .CLK(CK), .Q(n7436), .QN(n5565) );
  sdffs1 \DFF_880/Q_reg  ( .DIN(WX5976), .SDIN(n7434), .SSEL(test_se), .CLK(CK), .Q(n7435), .QN(n5569) );
  sdffs1 \DFF_879/Q_reg  ( .DIN(WX5974), .SDIN(n7433), .SSEL(test_se), .CLK(CK), .Q(n7434), .QN(n5573) );
  sdffs1 \DFF_878/Q_reg  ( .DIN(WX5972), .SDIN(n7432), .SSEL(test_se), .CLK(CK), .Q(n7433), .QN(n5578) );
  sdffs1 \DFF_877/Q_reg  ( .DIN(WX5970), .SDIN(n7431), .SSEL(test_se), .CLK(CK), .Q(n7432), .QN(n5583) );
  sdffs1 \DFF_876/Q_reg  ( .DIN(WX5968), .SDIN(n7430), .SSEL(test_se), .CLK(CK), .Q(n7431), .QN(n5588) );
  sdffs1 \DFF_875/Q_reg  ( .DIN(WX5966), .SDIN(n7429), .SSEL(test_se), .CLK(CK), .Q(n7430), .QN(n5593) );
  sdffs1 \DFF_874/Q_reg  ( .DIN(WX5964), .SDIN(n7428), .SSEL(test_se), .CLK(CK), .Q(n7429), .QN(n5598) );
  sdffs1 \DFF_873/Q_reg  ( .DIN(WX5962), .SDIN(n7427), .SSEL(test_se), .CLK(CK), .Q(n7428), .QN(n5603) );
  sdffs1 \DFF_872/Q_reg  ( .DIN(WX5960), .SDIN(n7426), .SSEL(test_se), .CLK(CK), .Q(n7427), .QN(n5608) );
  sdffs1 \DFF_871/Q_reg  ( .DIN(WX5958), .SDIN(n7425), .SSEL(test_se), .CLK(CK), .Q(n7426), .QN(n5613) );
  sdffs1 \DFF_870/Q_reg  ( .DIN(WX5956), .SDIN(n7424), .SSEL(test_se), .CLK(CK), .Q(n7425), .QN(n5618) );
  sdffs1 \DFF_869/Q_reg  ( .DIN(WX5954), .SDIN(n7423), .SSEL(test_se), .CLK(CK), .Q(n7424), .QN(n5623) );
  sdffs1 \DFF_868/Q_reg  ( .DIN(WX5952), .SDIN(n7422), .SSEL(test_se), .CLK(CK), .Q(n7423), .QN(n5628) );
  sdffs1 \DFF_867/Q_reg  ( .DIN(WX5950), .SDIN(n7421), .SSEL(test_se), .CLK(CK), .Q(n7422), .QN(n5633) );
  sdffs1 \DFF_866/Q_reg  ( .DIN(WX5948), .SDIN(n7420), .SSEL(test_se), .CLK(CK), .Q(n7421), .QN(n5638) );
  sdffs1 \DFF_865/Q_reg  ( .DIN(WX5946), .SDIN(n7419), .SSEL(test_se), .CLK(CK), .Q(n7420), .QN(n5643) );
  sdffs1 \DFF_864/Q_reg  ( .DIN(WX5944), .SDIN(n7418), .SSEL(test_se), .CLK(CK), .Q(n7419), .QN(n5648) );
  sdffs1 \DFF_863/Q_reg  ( .DIN(WX5942), .SDIN(n7417), .SSEL(test_se), .CLK(CK), .Q(n7418), .QN(n5508) );
  sdffs1 \DFF_862/Q_reg  ( .DIN(WX5940), .SDIN(n7416), .SSEL(test_se), .CLK(CK), .Q(n7417), .QN(n5512) );
  sdffs1 \DFF_861/Q_reg  ( .DIN(WX5938), .SDIN(n7415), .SSEL(test_se), .CLK(CK), .Q(n7416), .QN(n5516) );
  sdffs1 \DFF_860/Q_reg  ( .DIN(WX5936), .SDIN(n7414), .SSEL(test_se), .CLK(CK), .Q(n7415), .QN(n5520) );
  sdffs1 \DFF_859/Q_reg  ( .DIN(WX5934), .SDIN(n7413), .SSEL(test_se), .CLK(CK), .Q(n7414), .QN(n5524) );
  sdffs1 \DFF_858/Q_reg  ( .DIN(WX5932), .SDIN(n7412), .SSEL(test_se), .CLK(CK), .Q(n7413), .QN(n5528) );
  sdffs1 \DFF_857/Q_reg  ( .DIN(WX5930), .SDIN(n7411), .SSEL(test_se), .CLK(CK), .Q(n7412), .QN(n5532) );
  sdffs1 \DFF_856/Q_reg  ( .DIN(WX5928), .SDIN(n7410), .SSEL(test_se), .CLK(CK), .Q(n7411), .QN(n5536) );
  sdffs1 \DFF_855/Q_reg  ( .DIN(WX5926), .SDIN(n7409), .SSEL(test_se), .CLK(CK), .Q(n7410), .QN(n5540) );
  sdffs1 \DFF_854/Q_reg  ( .DIN(WX5924), .SDIN(n7408), .SSEL(test_se), .CLK(CK), .Q(n7409), .QN(n5544) );
  sdffs1 \DFF_853/Q_reg  ( .DIN(WX5922), .SDIN(n7407), .SSEL(test_se), .CLK(CK), .Q(n7408), .QN(n5548) );
  sdffs1 \DFF_852/Q_reg  ( .DIN(WX5920), .SDIN(n7406), .SSEL(test_se), .CLK(CK), .Q(n7407), .QN(n5552) );
  sdffs1 \DFF_851/Q_reg  ( .DIN(WX5918), .SDIN(n7405), .SSEL(test_se), .CLK(CK), .Q(n7406), .QN(n5556) );
  sdffs1 \DFF_850/Q_reg  ( .DIN(WX5916), .SDIN(n7404), .SSEL(test_se), .CLK(CK), .Q(n7405), .QN(n5560) );
  sdffs1 \DFF_849/Q_reg  ( .DIN(WX5914), .SDIN(n7403), .SSEL(test_se), .CLK(CK), .Q(n7404), .QN(n5564) );
  sdffs1 \DFF_848/Q_reg  ( .DIN(WX5912), .SDIN(n5572), .SSEL(test_se), .CLK(CK), .Q(n7403), .QN(n5568) );
  sdffs1 \DFF_847/Q_reg  ( .DIN(WX5910), .SDIN(n5577), .SSEL(test_se), .CLK(CK), .Q(n5572) );
  sdffs1 \DFF_846/Q_reg  ( .DIN(WX5908), .SDIN(n5582), .SSEL(test_se), .CLK(CK), .Q(n5577) );
  sdffs1 \DFF_845/Q_reg  ( .DIN(WX5906), .SDIN(n5587), .SSEL(test_se), .CLK(CK), .Q(n5582) );
  sdffs1 \DFF_844/Q_reg  ( .DIN(WX5904), .SDIN(n5592), .SSEL(test_se), .CLK(CK), .Q(n5587) );
  sdffs1 \DFF_843/Q_reg  ( .DIN(WX5902), .SDIN(n5597), .SSEL(test_se), .CLK(CK), .Q(n5592) );
  sdffs1 \DFF_842/Q_reg  ( .DIN(WX5900), .SDIN(n5602), .SSEL(test_se), .CLK(CK), .Q(n5597) );
  sdffs1 \DFF_841/Q_reg  ( .DIN(WX5898), .SDIN(n5607), .SSEL(test_se), .CLK(CK), .Q(n5602) );
  sdffs1 \DFF_840/Q_reg  ( .DIN(WX5896), .SDIN(n5612), .SSEL(test_se), .CLK(CK), .Q(n5607) );
  sdffs1 \DFF_839/Q_reg  ( .DIN(WX5894), .SDIN(n5617), .SSEL(test_se), .CLK(CK), .Q(n5612) );
  sdffs1 \DFF_838/Q_reg  ( .DIN(WX5892), .SDIN(n5622), .SSEL(test_se), .CLK(CK), .Q(n5617) );
  sdffs1 \DFF_837/Q_reg  ( .DIN(WX5890), .SDIN(n5627), .SSEL(test_se), .CLK(CK), .Q(n5622) );
  sdffs1 \DFF_836/Q_reg  ( .DIN(WX5888), .SDIN(n5632), .SSEL(test_se), .CLK(CK), .Q(n5627) );
  sdffs1 \DFF_835/Q_reg  ( .DIN(WX5886), .SDIN(n5637), .SSEL(test_se), .CLK(CK), .Q(n5632) );
  sdffs1 \DFF_834/Q_reg  ( .DIN(WX5884), .SDIN(n5642), .SSEL(test_se), .CLK(CK), .Q(n5637) );
  sdffs1 \DFF_833/Q_reg  ( .DIN(WX5882), .SDIN(n5647), .SSEL(test_se), .CLK(CK), .Q(n5642) );
  sdffs1 \DFF_832/Q_reg  ( .DIN(WX5880), .SDIN(n5507), .SSEL(test_se), .CLK(CK), .Q(n5647) );
  sdffs1 \DFF_831/Q_reg  ( .DIN(WX5878), .SDIN(n5511), .SSEL(test_se), .CLK(CK), .Q(n5507) );
  sdffs1 \DFF_830/Q_reg  ( .DIN(WX5876), .SDIN(n5515), .SSEL(test_se), .CLK(CK), .Q(n5511) );
  sdffs1 \DFF_829/Q_reg  ( .DIN(WX5874), .SDIN(n5519), .SSEL(test_se), .CLK(CK), .Q(n5515) );
  sdffs1 \DFF_828/Q_reg  ( .DIN(WX5872), .SDIN(n5523), .SSEL(test_se), .CLK(CK), .Q(n5519) );
  sdffs1 \DFF_827/Q_reg  ( .DIN(WX5870), .SDIN(n5527), .SSEL(test_se), .CLK(CK), .Q(n5523) );
  sdffs1 \DFF_826/Q_reg  ( .DIN(WX5868), .SDIN(n5531), .SSEL(test_se), .CLK(CK), .Q(n5527) );
  sdffs1 \DFF_825/Q_reg  ( .DIN(WX5866), .SDIN(n5535), .SSEL(test_se), .CLK(CK), .Q(n5531) );
  sdffs1 \DFF_824/Q_reg  ( .DIN(WX5864), .SDIN(n5539), .SSEL(test_se), .CLK(CK), .Q(n5535) );
  sdffs1 \DFF_823/Q_reg  ( .DIN(WX5862), .SDIN(n5543), .SSEL(test_se), .CLK(CK), .Q(n5539) );
  sdffs1 \DFF_822/Q_reg  ( .DIN(WX5860), .SDIN(n5547), .SSEL(test_se), .CLK(CK), .Q(n5543) );
  sdffs1 \DFF_821/Q_reg  ( .DIN(WX5858), .SDIN(n5551), .SSEL(test_se), .CLK(CK), .Q(n5547) );
  sdffs1 \DFF_820/Q_reg  ( .DIN(WX5856), .SDIN(n5555), .SSEL(test_se), .CLK(CK), .Q(n5551) );
  sdffs1 \DFF_819/Q_reg  ( .DIN(WX5854), .SDIN(n5559), .SSEL(test_se), .CLK(CK), .Q(n5555) );
  sdffs1 \DFF_818/Q_reg  ( .DIN(WX5852), .SDIN(n5563), .SSEL(test_se), .CLK(CK), .Q(n5559) );
  sdffs1 \DFF_817/Q_reg  ( .DIN(WX5850), .SDIN(n5567), .SSEL(test_se), .CLK(CK), .Q(n5563) );
  sdffs1 \DFF_816/Q_reg  ( .DIN(WX5848), .SDIN(n7402), .SSEL(test_se), .CLK(CK), .Q(n5567) );
  sdffs1 \DFF_815/Q_reg  ( .DIN(WX5846), .SDIN(n7401), .SSEL(test_se), .CLK(CK), .Q(n7402), .QN(n5571) );
  sdffs1 \DFF_814/Q_reg  ( .DIN(WX5844), .SDIN(n7400), .SSEL(test_se), .CLK(CK), .Q(n7401), .QN(n5576) );
  sdffs1 \DFF_813/Q_reg  ( .DIN(WX5842), .SDIN(n7399), .SSEL(test_se), .CLK(CK), .Q(n7400), .QN(n5581) );
  sdffs1 \DFF_812/Q_reg  ( .DIN(WX5840), .SDIN(n7398), .SSEL(test_se), .CLK(CK), .Q(n7399), .QN(n5586) );
  sdffs1 \DFF_811/Q_reg  ( .DIN(WX5838), .SDIN(n7397), .SSEL(test_se), .CLK(CK), .Q(n7398), .QN(n5591) );
  sdffs1 \DFF_810/Q_reg  ( .DIN(WX5836), .SDIN(n7396), .SSEL(test_se), .CLK(CK), .Q(n7397), .QN(n5596) );
  sdffs1 \DFF_809/Q_reg  ( .DIN(WX5834), .SDIN(n7395), .SSEL(test_se), .CLK(CK), .Q(n7396), .QN(n5601) );
  sdffs1 \DFF_808/Q_reg  ( .DIN(WX5832), .SDIN(n7394), .SSEL(test_se), .CLK(CK), .Q(n7395), .QN(n5606) );
  sdffs1 \DFF_807/Q_reg  ( .DIN(WX5830), .SDIN(n7393), .SSEL(test_se), .CLK(CK), .Q(n7394), .QN(n5611) );
  sdffs1 \DFF_806/Q_reg  ( .DIN(WX5828), .SDIN(n7392), .SSEL(test_se), .CLK(CK), .Q(n7393), .QN(n5616) );
  sdffs1 \DFF_805/Q_reg  ( .DIN(WX5826), .SDIN(n7391), .SSEL(test_se), .CLK(CK), .Q(n7392), .QN(n5621) );
  sdffs1 \DFF_804/Q_reg  ( .DIN(WX5824), .SDIN(n7390), .SSEL(test_se), .CLK(CK), .Q(n7391), .QN(n5626) );
  sdffs1 \DFF_803/Q_reg  ( .DIN(WX5822), .SDIN(n7389), .SSEL(test_se), .CLK(CK), .Q(n7390), .QN(n5631) );
  sdffs1 \DFF_802/Q_reg  ( .DIN(WX5820), .SDIN(n7388), .SSEL(test_se), .CLK(CK), .Q(n7389), .QN(n5636) );
  sdffs1 \DFF_801/Q_reg  ( .DIN(WX5818), .SDIN(n7387), .SSEL(test_se), .CLK(CK), .Q(n7388), .QN(n5641) );
  sdffs1 \DFF_800/Q_reg  ( .DIN(WX5816), .SDIN(n7386), .SSEL(test_se), .CLK(CK), .Q(n7387), .QN(n5646) );
  sdffs1 \DFF_799/Q_reg  ( .DIN(WX5718), .SDIN(n7385), .SSEL(test_se), .CLK(CK), .Q(n7386), .QN(n5476) );
  sdffs1 \DFF_798/Q_reg  ( .DIN(WX5716), .SDIN(n7384), .SSEL(test_se), .CLK(CK), .Q(n7385), .QN(n5477) );
  sdffs1 \DFF_797/Q_reg  ( .DIN(WX5714), .SDIN(n7383), .SSEL(test_se), .CLK(CK), .Q(n7384), .QN(n5478) );
  sdffs1 \DFF_796/Q_reg  ( .DIN(WX5712), .SDIN(n7382), .SSEL(test_se), .CLK(CK), .Q(n7383), .QN(n5479) );
  sdffs1 \DFF_795/Q_reg  ( .DIN(WX5710), .SDIN(n7381), .SSEL(test_se), .CLK(CK), .Q(n7382), .QN(n5480) );
  sdffs1 \DFF_794/Q_reg  ( .DIN(WX5708), .SDIN(n7380), .SSEL(test_se), .CLK(CK), .Q(n7381), .QN(n5481) );
  sdffs1 \DFF_793/Q_reg  ( .DIN(WX5706), .SDIN(n7379), .SSEL(test_se), .CLK(CK), .Q(n7380), .QN(n5482) );
  sdffs1 \DFF_792/Q_reg  ( .DIN(WX5704), .SDIN(n7378), .SSEL(test_se), .CLK(CK), .Q(n7379), .QN(n5483) );
  sdffs1 \DFF_791/Q_reg  ( .DIN(WX5702), .SDIN(n7377), .SSEL(test_se), .CLK(CK), .Q(n7378), .QN(n5484) );
  sdffs1 \DFF_790/Q_reg  ( .DIN(WX5700), .SDIN(n7376), .SSEL(test_se), .CLK(CK), .Q(n7377), .QN(n5485) );
  sdffs1 \DFF_789/Q_reg  ( .DIN(WX5698), .SDIN(n7375), .SSEL(test_se), .CLK(CK), .Q(n7376), .QN(n5486) );
  sdffs1 \DFF_788/Q_reg  ( .DIN(WX5696), .SDIN(n7374), .SSEL(test_se), .CLK(CK), .Q(n7375), .QN(n5487) );
  sdffs1 \DFF_787/Q_reg  ( .DIN(WX5694), .SDIN(n7373), .SSEL(test_se), .CLK(CK), .Q(n7374), .QN(n5488) );
  sdffs1 \DFF_786/Q_reg  ( .DIN(WX5692), .SDIN(n7372), .SSEL(test_se), .CLK(CK), .Q(n7373), .QN(n5489) );
  sdffs1 \DFF_785/Q_reg  ( .DIN(WX5690), .SDIN(n7371), .SSEL(test_se), .CLK(CK), .Q(n7372), .QN(n5490) );
  sdffs1 \DFF_784/Q_reg  ( .DIN(WX5688), .SDIN(n7370), .SSEL(test_se), .CLK(CK), .Q(n7371), .QN(n5491) );
  sdffs1 \DFF_783/Q_reg  ( .DIN(WX5686), .SDIN(n7369), .SSEL(test_se), .CLK(CK), .Q(n7370), .QN(n5492) );
  sdffs1 \DFF_782/Q_reg  ( .DIN(WX5684), .SDIN(n7368), .SSEL(test_se), .CLK(CK), .Q(n7369), .QN(n5493) );
  sdffs1 \DFF_781/Q_reg  ( .DIN(WX5682), .SDIN(n7367), .SSEL(test_se), .CLK(CK), .Q(n7368), .QN(n5494) );
  sdffs1 \DFF_780/Q_reg  ( .DIN(WX5680), .SDIN(n7366), .SSEL(test_se), .CLK(CK), .Q(n7367), .QN(n5495) );
  sdffs1 \DFF_779/Q_reg  ( .DIN(WX5678), .SDIN(n7365), .SSEL(test_se), .CLK(CK), .Q(n7366), .QN(n5496) );
  sdffs1 \DFF_778/Q_reg  ( .DIN(WX5676), .SDIN(n7364), .SSEL(test_se), .CLK(CK), .Q(n7365), .QN(n5497) );
  sdffs1 \DFF_777/Q_reg  ( .DIN(WX5674), .SDIN(n7363), .SSEL(test_se), .CLK(CK), .Q(n7364), .QN(n5498) );
  sdffs1 \DFF_776/Q_reg  ( .DIN(WX5672), .SDIN(n7362), .SSEL(test_se), .CLK(CK), .Q(n7363), .QN(n5499) );
  sdffs1 \DFF_775/Q_reg  ( .DIN(WX5670), .SDIN(n7361), .SSEL(test_se), .CLK(CK), .Q(n7362), .QN(n5500) );
  sdffs1 \DFF_774/Q_reg  ( .DIN(WX5668), .SDIN(n7360), .SSEL(test_se), .CLK(CK), .Q(n7361), .QN(n5501) );
  sdffs1 \DFF_773/Q_reg  ( .DIN(WX5666), .SDIN(n7359), .SSEL(test_se), .CLK(CK), .Q(n7360), .QN(n5502) );
  sdffs1 \DFF_772/Q_reg  ( .DIN(WX5664), .SDIN(n7358), .SSEL(test_se), .CLK(CK), .Q(n7359), .QN(n5503) );
  sdffs1 \DFF_771/Q_reg  ( .DIN(WX5662), .SDIN(n7357), .SSEL(test_se), .CLK(CK), .Q(n7358), .QN(n5504) );
  sdffs1 \DFF_770/Q_reg  ( .DIN(WX5660), .SDIN(n7356), .SSEL(test_se), .CLK(CK), .Q(n7357), .QN(n5505) );
  sdffs1 \DFF_769/Q_reg  ( .DIN(WX5658), .SDIN(n7355), .SSEL(test_se), .CLK(CK), .Q(n7356), .QN(n5506) );
  sdffs1 \DFF_768/Q_reg  ( .DIN(WX5656), .SDIN(CRC_OUT_6_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7355), .QN(n5475) );
  sdffs1 \DFF_767/Q_reg  ( .DIN(WX5205), .SDIN(CRC_OUT_6_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_31), .QN(n5650) );
  sdffs1 \DFF_766/Q_reg  ( .DIN(WX5203), .SDIN(CRC_OUT_6_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_30), .QN(n5645) );
  sdffs1 \DFF_765/Q_reg  ( .DIN(WX5201), .SDIN(CRC_OUT_6_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_29), .QN(n5640) );
  sdffs1 \DFF_764/Q_reg  ( .DIN(WX5199), .SDIN(CRC_OUT_6_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_28), .QN(n5635) );
  sdffs1 \DFF_763/Q_reg  ( .DIN(WX5197), .SDIN(CRC_OUT_6_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_27), .QN(n5630) );
  sdffs1 \DFF_762/Q_reg  ( .DIN(WX5195), .SDIN(CRC_OUT_6_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_26), .QN(n5625) );
  sdffs1 \DFF_761/Q_reg  ( .DIN(WX5193), .SDIN(CRC_OUT_6_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_25), .QN(n5620) );
  sdffs1 \DFF_760/Q_reg  ( .DIN(WX5191), .SDIN(CRC_OUT_6_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_24), .QN(n5615) );
  sdffs1 \DFF_759/Q_reg  ( .DIN(WX5189), .SDIN(CRC_OUT_6_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_23), .QN(n5610) );
  sdffs1 \DFF_758/Q_reg  ( .DIN(WX5187), .SDIN(CRC_OUT_6_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_22), .QN(n5605) );
  sdffs1 \DFF_757/Q_reg  ( .DIN(WX5185), .SDIN(CRC_OUT_6_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_21), .QN(n5600) );
  sdffs1 \DFF_756/Q_reg  ( .DIN(WX5183), .SDIN(CRC_OUT_6_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_20), .QN(n5595) );
  sdffs1 \DFF_755/Q_reg  ( .DIN(WX5181), .SDIN(CRC_OUT_6_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_19), .QN(n5590) );
  sdffs1 \DFF_754/Q_reg  ( .DIN(WX5179), .SDIN(CRC_OUT_6_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_18), .QN(n5585) );
  sdffs1 \DFF_753/Q_reg  ( .DIN(WX5177), .SDIN(CRC_OUT_6_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_17), .QN(n5580) );
  sdffs1 \DFF_752/Q_reg  ( .DIN(WX5175), .SDIN(CRC_OUT_6_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_16), .QN(n5575) );
  sdffs1 \DFF_751/Q_reg  ( .DIN(WX5173), .SDIN(CRC_OUT_6_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_15), .QN(n5570) );
  sdffs1 \DFF_750/Q_reg  ( .DIN(WX5171), .SDIN(CRC_OUT_6_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_14), .QN(n5566) );
  sdffs1 \DFF_749/Q_reg  ( .DIN(WX5169), .SDIN(CRC_OUT_6_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_13), .QN(n5562) );
  sdffs1 \DFF_748/Q_reg  ( .DIN(WX5167), .SDIN(CRC_OUT_6_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_12), .QN(n5558) );
  sdffs1 \DFF_747/Q_reg  ( .DIN(WX5165), .SDIN(CRC_OUT_6_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_11), .QN(n5554) );
  sdffs1 \DFF_746/Q_reg  ( .DIN(WX5163), .SDIN(CRC_OUT_6_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_10), .QN(n5550) );
  sdffs1 \DFF_745/Q_reg  ( .DIN(WX5161), .SDIN(CRC_OUT_6_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_9), .QN(n5546) );
  sdffs1 \DFF_744/Q_reg  ( .DIN(WX5159), .SDIN(CRC_OUT_6_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_8), .QN(n5542) );
  sdffs1 \DFF_743/Q_reg  ( .DIN(WX5157), .SDIN(CRC_OUT_6_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_7), .QN(n5538) );
  sdffs1 \DFF_742/Q_reg  ( .DIN(WX5155), .SDIN(CRC_OUT_6_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_6), .QN(n5534) );
  sdffs1 \DFF_741/Q_reg  ( .DIN(WX5153), .SDIN(CRC_OUT_6_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_5), .QN(n5530) );
  sdffs1 \DFF_740/Q_reg  ( .DIN(WX5151), .SDIN(CRC_OUT_6_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_4), .QN(n5526) );
  sdffs1 \DFF_739/Q_reg  ( .DIN(WX5149), .SDIN(CRC_OUT_6_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_3), .QN(n5522) );
  sdffs1 \DFF_738/Q_reg  ( .DIN(WX5147), .SDIN(CRC_OUT_6_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_2), .QN(n5518) );
  sdffs1 \DFF_737/Q_reg  ( .DIN(WX5145), .SDIN(CRC_OUT_6_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_6_1), .QN(n5514) );
  sdffs1 \DFF_736/Q_reg  ( .DIN(WX5143), .SDIN(n7354), .SSEL(test_se), .CLK(CK), .Q(CRC_OUT_6_0), .QN(n5510) );
  sdffs1 \DFF_735/Q_reg  ( .DIN(WX4777), .SDIN(n7353), .SSEL(test_se), .CLK(CK), .Q(n7354), .QN(n3269) );
  sdffs1 \DFF_734/Q_reg  ( .DIN(WX4775), .SDIN(n7352), .SSEL(test_se), .CLK(CK), .Q(n7353), .QN(n3270) );
  sdffs1 \DFF_733/Q_reg  ( .DIN(WX4773), .SDIN(n7351), .SSEL(test_se), .CLK(CK), .Q(n7352), .QN(n3271) );
  sdffs1 \DFF_732/Q_reg  ( .DIN(WX4771), .SDIN(n7350), .SSEL(test_se), .CLK(CK), .Q(n7351), .QN(n3272) );
  sdffs1 \DFF_731/Q_reg  ( .DIN(WX4769), .SDIN(n7349), .SSEL(test_se), .CLK(CK), .Q(n7350), .QN(n3273) );
  sdffs1 \DFF_730/Q_reg  ( .DIN(WX4767), .SDIN(n7348), .SSEL(test_se), .CLK(CK), .Q(n7349), .QN(n3274) );
  sdffs1 \DFF_729/Q_reg  ( .DIN(WX4765), .SDIN(n7347), .SSEL(test_se), .CLK(CK), .Q(n7348), .QN(n3275) );
  sdffs1 \DFF_728/Q_reg  ( .DIN(WX4763), .SDIN(n7346), .SSEL(test_se), .CLK(CK), .Q(n7347), .QN(n3276) );
  sdffs1 \DFF_727/Q_reg  ( .DIN(WX4761), .SDIN(n7345), .SSEL(test_se), .CLK(CK), .Q(n7346), .QN(n3277) );
  sdffs1 \DFF_726/Q_reg  ( .DIN(WX4759), .SDIN(n7344), .SSEL(test_se), .CLK(CK), .Q(n7345), .QN(n3278) );
  sdffs1 \DFF_725/Q_reg  ( .DIN(WX4757), .SDIN(n7343), .SSEL(test_se), .CLK(CK), .Q(n7344), .QN(n3279) );
  sdffs1 \DFF_724/Q_reg  ( .DIN(WX4755), .SDIN(n7342), .SSEL(test_se), .CLK(CK), .Q(n7343), .QN(n3280) );
  sdffs1 \DFF_723/Q_reg  ( .DIN(WX4753), .SDIN(n7341), .SSEL(test_se), .CLK(CK), .Q(n7342), .QN(n3281) );
  sdffs1 \DFF_722/Q_reg  ( .DIN(WX4751), .SDIN(n7340), .SSEL(test_se), .CLK(CK), .Q(n7341), .QN(n3282) );
  sdffs1 \DFF_721/Q_reg  ( .DIN(WX4749), .SDIN(n7339), .SSEL(test_se), .CLK(CK), .Q(n7340), .QN(n3283) );
  sdffs1 \DFF_720/Q_reg  ( .DIN(WX4747), .SDIN(n7338), .SSEL(test_se), .CLK(CK), .Q(n7339), .QN(n3284) );
  sdffs1 \DFF_719/Q_reg  ( .DIN(WX4745), .SDIN(n7337), .SSEL(test_se), .CLK(CK), .Q(n7338), .QN(n5750) );
  sdffs1 \DFF_718/Q_reg  ( .DIN(WX4743), .SDIN(n7336), .SSEL(test_se), .CLK(CK), .Q(n7337), .QN(n5755) );
  sdffs1 \DFF_717/Q_reg  ( .DIN(WX4741), .SDIN(n7335), .SSEL(test_se), .CLK(CK), .Q(n7336), .QN(n5760) );
  sdffs1 \DFF_716/Q_reg  ( .DIN(WX4739), .SDIN(n7334), .SSEL(test_se), .CLK(CK), .Q(n7335), .QN(n5765) );
  sdffs1 \DFF_715/Q_reg  ( .DIN(WX4737), .SDIN(n7333), .SSEL(test_se), .CLK(CK), .Q(n7334), .QN(n5770) );
  sdffs1 \DFF_714/Q_reg  ( .DIN(WX4735), .SDIN(n7332), .SSEL(test_se), .CLK(CK), .Q(n7333), .QN(n5775) );
  sdffs1 \DFF_713/Q_reg  ( .DIN(WX4733), .SDIN(n7331), .SSEL(test_se), .CLK(CK), .Q(n7332), .QN(n5780) );
  sdffs1 \DFF_712/Q_reg  ( .DIN(WX4731), .SDIN(n7330), .SSEL(test_se), .CLK(CK), .Q(n7331), .QN(n5785) );
  sdffs1 \DFF_711/Q_reg  ( .DIN(WX4729), .SDIN(n7329), .SSEL(test_se), .CLK(CK), .Q(n7330), .QN(n5790) );
  sdffs1 \DFF_710/Q_reg  ( .DIN(WX4727), .SDIN(n7328), .SSEL(test_se), .CLK(CK), .Q(n7329), .QN(n5795) );
  sdffs1 \DFF_709/Q_reg  ( .DIN(WX4725), .SDIN(n7327), .SSEL(test_se), .CLK(CK), .Q(n7328), .QN(n5800) );
  sdffs1 \DFF_708/Q_reg  ( .DIN(WX4723), .SDIN(n7326), .SSEL(test_se), .CLK(CK), .Q(n7327), .QN(n5805) );
  sdffs1 \DFF_707/Q_reg  ( .DIN(WX4721), .SDIN(n7325), .SSEL(test_se), .CLK(CK), .Q(n7326), .QN(n5810) );
  sdffs1 \DFF_706/Q_reg  ( .DIN(WX4719), .SDIN(n7324), .SSEL(test_se), .CLK(CK), .Q(n7325), .QN(n5815) );
  sdffs1 \DFF_705/Q_reg  ( .DIN(WX4717), .SDIN(n7323), .SSEL(test_se), .CLK(CK), .Q(n7324), .QN(n5820) );
  sdffs1 \DFF_704/Q_reg  ( .DIN(WX4715), .SDIN(n7322), .SSEL(test_se), .CLK(CK), .Q(n7323), .QN(n5825) );
  sdffs1 \DFF_703/Q_reg  ( .DIN(WX4713), .SDIN(n7321), .SSEL(test_se), .CLK(CK), .Q(n7322), .QN(n5685) );
  sdffs1 \DFF_702/Q_reg  ( .DIN(WX4711), .SDIN(n7320), .SSEL(test_se), .CLK(CK), .Q(n7321), .QN(n5689) );
  sdffs1 \DFF_701/Q_reg  ( .DIN(WX4709), .SDIN(n7319), .SSEL(test_se), .CLK(CK), .Q(n7320), .QN(n5693) );
  sdffs1 \DFF_700/Q_reg  ( .DIN(WX4707), .SDIN(n7318), .SSEL(test_se), .CLK(CK), .Q(n7319), .QN(n5697) );
  sdffs1 \DFF_699/Q_reg  ( .DIN(WX4705), .SDIN(n7317), .SSEL(test_se), .CLK(CK), .Q(n7318), .QN(n5701) );
  sdffs1 \DFF_698/Q_reg  ( .DIN(WX4703), .SDIN(n7316), .SSEL(test_se), .CLK(CK), .Q(n7317), .QN(n5705) );
  sdffs1 \DFF_697/Q_reg  ( .DIN(WX4701), .SDIN(n7315), .SSEL(test_se), .CLK(CK), .Q(n7316), .QN(n5709) );
  sdffs1 \DFF_696/Q_reg  ( .DIN(WX4699), .SDIN(n7314), .SSEL(test_se), .CLK(CK), .Q(n7315), .QN(n5713) );
  sdffs1 \DFF_695/Q_reg  ( .DIN(WX4697), .SDIN(n7313), .SSEL(test_se), .CLK(CK), .Q(n7314), .QN(n5717) );
  sdffs1 \DFF_694/Q_reg  ( .DIN(WX4695), .SDIN(n7312), .SSEL(test_se), .CLK(CK), .Q(n7313), .QN(n5721) );
  sdffs1 \DFF_693/Q_reg  ( .DIN(WX4693), .SDIN(n7311), .SSEL(test_se), .CLK(CK), .Q(n7312), .QN(n5725) );
  sdffs1 \DFF_692/Q_reg  ( .DIN(WX4691), .SDIN(n7310), .SSEL(test_se), .CLK(CK), .Q(n7311), .QN(n5729) );
  sdffs1 \DFF_691/Q_reg  ( .DIN(WX4689), .SDIN(n7309), .SSEL(test_se), .CLK(CK), .Q(n7310), .QN(n5733) );
  sdffs1 \DFF_690/Q_reg  ( .DIN(WX4687), .SDIN(n7308), .SSEL(test_se), .CLK(CK), .Q(n7309), .QN(n5737) );
  sdffs1 \DFF_689/Q_reg  ( .DIN(WX4685), .SDIN(n7307), .SSEL(test_se), .CLK(CK), .Q(n7308), .QN(n5741) );
  sdffs1 \DFF_688/Q_reg  ( .DIN(WX4683), .SDIN(n7306), .SSEL(test_se), .CLK(CK), .Q(n7307), .QN(n5745) );
  sdffs1 \DFF_687/Q_reg  ( .DIN(WX4681), .SDIN(n7305), .SSEL(test_se), .CLK(CK), .Q(n7306), .QN(n5749) );
  sdffs1 \DFF_686/Q_reg  ( .DIN(WX4679), .SDIN(n7304), .SSEL(test_se), .CLK(CK), .Q(n7305), .QN(n5754) );
  sdffs1 \DFF_685/Q_reg  ( .DIN(WX4677), .SDIN(n7303), .SSEL(test_se), .CLK(CK), .Q(n7304), .QN(n5759) );
  sdffs1 \DFF_684/Q_reg  ( .DIN(WX4675), .SDIN(n7302), .SSEL(test_se), .CLK(CK), .Q(n7303), .QN(n5764) );
  sdffs1 \DFF_683/Q_reg  ( .DIN(WX4673), .SDIN(n7301), .SSEL(test_se), .CLK(CK), .Q(n7302), .QN(n5769) );
  sdffs1 \DFF_682/Q_reg  ( .DIN(WX4671), .SDIN(n7300), .SSEL(test_se), .CLK(CK), .Q(n7301), .QN(n5774) );
  sdffs1 \DFF_681/Q_reg  ( .DIN(WX4669), .SDIN(n7299), .SSEL(test_se), .CLK(CK), .Q(n7300), .QN(n5779) );
  sdffs1 \DFF_680/Q_reg  ( .DIN(WX4667), .SDIN(n7298), .SSEL(test_se), .CLK(CK), .Q(n7299), .QN(n5784) );
  sdffs1 \DFF_679/Q_reg  ( .DIN(WX4665), .SDIN(n7297), .SSEL(test_se), .CLK(CK), .Q(n7298), .QN(n5789) );
  sdffs1 \DFF_678/Q_reg  ( .DIN(WX4663), .SDIN(n7296), .SSEL(test_se), .CLK(CK), .Q(n7297), .QN(n5794) );
  sdffs1 \DFF_677/Q_reg  ( .DIN(WX4661), .SDIN(n7295), .SSEL(test_se), .CLK(CK), .Q(n7296), .QN(n5799) );
  sdffs1 \DFF_676/Q_reg  ( .DIN(WX4659), .SDIN(n7294), .SSEL(test_se), .CLK(CK), .Q(n7295), .QN(n5804) );
  sdffs1 \DFF_675/Q_reg  ( .DIN(WX4657), .SDIN(n7293), .SSEL(test_se), .CLK(CK), .Q(n7294), .QN(n5809) );
  sdffs1 \DFF_674/Q_reg  ( .DIN(WX4655), .SDIN(n7292), .SSEL(test_se), .CLK(CK), .Q(n7293), .QN(n5814) );
  sdffs1 \DFF_673/Q_reg  ( .DIN(WX4653), .SDIN(n7291), .SSEL(test_se), .CLK(CK), .Q(n7292), .QN(n5819) );
  sdffs1 \DFF_672/Q_reg  ( .DIN(WX4651), .SDIN(n7290), .SSEL(test_se), .CLK(CK), .Q(n7291), .QN(n5824) );
  sdffs1 \DFF_671/Q_reg  ( .DIN(WX4649), .SDIN(n7289), .SSEL(test_se), .CLK(CK), .Q(n7290), .QN(n5684) );
  sdffs1 \DFF_670/Q_reg  ( .DIN(WX4647), .SDIN(n7288), .SSEL(test_se), .CLK(CK), .Q(n7289), .QN(n5688) );
  sdffs1 \DFF_669/Q_reg  ( .DIN(WX4645), .SDIN(n7287), .SSEL(test_se), .CLK(CK), .Q(n7288), .QN(n5692) );
  sdffs1 \DFF_668/Q_reg  ( .DIN(WX4643), .SDIN(n7286), .SSEL(test_se), .CLK(CK), .Q(n7287), .QN(n5696) );
  sdffs1 \DFF_667/Q_reg  ( .DIN(WX4641), .SDIN(n7285), .SSEL(test_se), .CLK(CK), .Q(n7286), .QN(n5700) );
  sdffs1 \DFF_666/Q_reg  ( .DIN(WX4639), .SDIN(n7284), .SSEL(test_se), .CLK(CK), .Q(n7285), .QN(n5704) );
  sdffs1 \DFF_665/Q_reg  ( .DIN(WX4637), .SDIN(n7283), .SSEL(test_se), .CLK(CK), .Q(n7284), .QN(n5708) );
  sdffs1 \DFF_664/Q_reg  ( .DIN(WX4635), .SDIN(n7282), .SSEL(test_se), .CLK(CK), .Q(n7283), .QN(n5712) );
  sdffs1 \DFF_663/Q_reg  ( .DIN(WX4633), .SDIN(n7281), .SSEL(test_se), .CLK(CK), .Q(n7282), .QN(n5716) );
  sdffs1 \DFF_662/Q_reg  ( .DIN(WX4631), .SDIN(n7280), .SSEL(test_se), .CLK(CK), .Q(n7281), .QN(n5720) );
  sdffs1 \DFF_661/Q_reg  ( .DIN(WX4629), .SDIN(n7279), .SSEL(test_se), .CLK(CK), .Q(n7280), .QN(n5724) );
  sdffs1 \DFF_660/Q_reg  ( .DIN(WX4627), .SDIN(n7278), .SSEL(test_se), .CLK(CK), .Q(n7279), .QN(n5728) );
  sdffs1 \DFF_659/Q_reg  ( .DIN(WX4625), .SDIN(n7277), .SSEL(test_se), .CLK(CK), .Q(n7278), .QN(n5732) );
  sdffs1 \DFF_658/Q_reg  ( .DIN(WX4623), .SDIN(n7276), .SSEL(test_se), .CLK(CK), .Q(n7277), .QN(n5736) );
  sdffs1 \DFF_657/Q_reg  ( .DIN(WX4621), .SDIN(n7275), .SSEL(test_se), .CLK(CK), .Q(n7276), .QN(n5740) );
  sdffs1 \DFF_656/Q_reg  ( .DIN(WX4619), .SDIN(n5748), .SSEL(test_se), .CLK(CK), .Q(n7275), .QN(n5744) );
  sdffs1 \DFF_655/Q_reg  ( .DIN(WX4617), .SDIN(n5753), .SSEL(test_se), .CLK(CK), .Q(n5748) );
  sdffs1 \DFF_654/Q_reg  ( .DIN(WX4615), .SDIN(n5758), .SSEL(test_se), .CLK(CK), .Q(n5753) );
  sdffs1 \DFF_653/Q_reg  ( .DIN(WX4613), .SDIN(n5763), .SSEL(test_se), .CLK(CK), .Q(n5758) );
  sdffs1 \DFF_652/Q_reg  ( .DIN(WX4611), .SDIN(n5768), .SSEL(test_se), .CLK(CK), .Q(n5763) );
  sdffs1 \DFF_651/Q_reg  ( .DIN(WX4609), .SDIN(n5773), .SSEL(test_se), .CLK(CK), .Q(n5768) );
  sdffs1 \DFF_650/Q_reg  ( .DIN(WX4607), .SDIN(n5778), .SSEL(test_se), .CLK(CK), .Q(n5773) );
  sdffs1 \DFF_649/Q_reg  ( .DIN(WX4605), .SDIN(n5783), .SSEL(test_se), .CLK(CK), .Q(n5778) );
  sdffs1 \DFF_648/Q_reg  ( .DIN(WX4603), .SDIN(n5788), .SSEL(test_se), .CLK(CK), .Q(n5783) );
  sdffs1 \DFF_647/Q_reg  ( .DIN(WX4601), .SDIN(n5793), .SSEL(test_se), .CLK(CK), .Q(n5788) );
  sdffs1 \DFF_646/Q_reg  ( .DIN(WX4599), .SDIN(n5798), .SSEL(test_se), .CLK(CK), .Q(n5793) );
  sdffs1 \DFF_645/Q_reg  ( .DIN(WX4597), .SDIN(n5803), .SSEL(test_se), .CLK(CK), .Q(n5798) );
  sdffs1 \DFF_644/Q_reg  ( .DIN(WX4595), .SDIN(n5808), .SSEL(test_se), .CLK(CK), .Q(n5803) );
  sdffs1 \DFF_643/Q_reg  ( .DIN(WX4593), .SDIN(n5813), .SSEL(test_se), .CLK(CK), .Q(n5808) );
  sdffs1 \DFF_642/Q_reg  ( .DIN(WX4591), .SDIN(n5818), .SSEL(test_se), .CLK(CK), .Q(n5813) );
  sdffs1 \DFF_641/Q_reg  ( .DIN(WX4589), .SDIN(n5823), .SSEL(test_se), .CLK(CK), .Q(n5818) );
  sdffs1 \DFF_640/Q_reg  ( .DIN(WX4587), .SDIN(n5683), .SSEL(test_se), .CLK(CK), .Q(n5823) );
  sdffs1 \DFF_639/Q_reg  ( .DIN(WX4585), .SDIN(n5687), .SSEL(test_se), .CLK(CK), .Q(n5683) );
  sdffs1 \DFF_638/Q_reg  ( .DIN(WX4583), .SDIN(n5691), .SSEL(test_se), .CLK(CK), .Q(n5687) );
  sdffs1 \DFF_637/Q_reg  ( .DIN(WX4581), .SDIN(n5695), .SSEL(test_se), .CLK(CK), .Q(n5691) );
  sdffs1 \DFF_636/Q_reg  ( .DIN(WX4579), .SDIN(n5699), .SSEL(test_se), .CLK(CK), .Q(n5695) );
  sdffs1 \DFF_635/Q_reg  ( .DIN(WX4577), .SDIN(n5703), .SSEL(test_se), .CLK(CK), .Q(n5699) );
  sdffs1 \DFF_634/Q_reg  ( .DIN(WX4575), .SDIN(n5707), .SSEL(test_se), .CLK(CK), .Q(n5703) );
  sdffs1 \DFF_633/Q_reg  ( .DIN(WX4573), .SDIN(n5711), .SSEL(test_se), .CLK(CK), .Q(n5707) );
  sdffs1 \DFF_632/Q_reg  ( .DIN(WX4571), .SDIN(n5715), .SSEL(test_se), .CLK(CK), .Q(n5711) );
  sdffs1 \DFF_631/Q_reg  ( .DIN(WX4569), .SDIN(n5719), .SSEL(test_se), .CLK(CK), .Q(n5715) );
  sdffs1 \DFF_630/Q_reg  ( .DIN(WX4567), .SDIN(n5723), .SSEL(test_se), .CLK(CK), .Q(n5719) );
  sdffs1 \DFF_629/Q_reg  ( .DIN(WX4565), .SDIN(n5727), .SSEL(test_se), .CLK(CK), .Q(n5723) );
  sdffs1 \DFF_628/Q_reg  ( .DIN(WX4563), .SDIN(n5731), .SSEL(test_se), .CLK(CK), .Q(n5727) );
  sdffs1 \DFF_627/Q_reg  ( .DIN(WX4561), .SDIN(n5735), .SSEL(test_se), .CLK(CK), .Q(n5731) );
  sdffs1 \DFF_626/Q_reg  ( .DIN(WX4559), .SDIN(n5739), .SSEL(test_se), .CLK(CK), .Q(n5735) );
  sdffs1 \DFF_625/Q_reg  ( .DIN(WX4557), .SDIN(n5743), .SSEL(test_se), .CLK(CK), .Q(n5739) );
  sdffs1 \DFF_624/Q_reg  ( .DIN(WX4555), .SDIN(n7274), .SSEL(test_se), .CLK(CK), .Q(n5743) );
  sdffs1 \DFF_623/Q_reg  ( .DIN(WX4553), .SDIN(n7273), .SSEL(test_se), .CLK(CK), .Q(n7274), .QN(n5747) );
  sdffs1 \DFF_622/Q_reg  ( .DIN(WX4551), .SDIN(n7272), .SSEL(test_se), .CLK(CK), .Q(n7273), .QN(n5752) );
  sdffs1 \DFF_621/Q_reg  ( .DIN(WX4549), .SDIN(n7271), .SSEL(test_se), .CLK(CK), .Q(n7272), .QN(n5757) );
  sdffs1 \DFF_620/Q_reg  ( .DIN(WX4547), .SDIN(n7270), .SSEL(test_se), .CLK(CK), .Q(n7271), .QN(n5762) );
  sdffs1 \DFF_619/Q_reg  ( .DIN(WX4545), .SDIN(n7269), .SSEL(test_se), .CLK(CK), .Q(n7270), .QN(n5767) );
  sdffs1 \DFF_618/Q_reg  ( .DIN(WX4543), .SDIN(n7268), .SSEL(test_se), .CLK(CK), .Q(n7269), .QN(n5772) );
  sdffs1 \DFF_617/Q_reg  ( .DIN(WX4541), .SDIN(n7267), .SSEL(test_se), .CLK(CK), .Q(n7268), .QN(n5777) );
  sdffs1 \DFF_616/Q_reg  ( .DIN(WX4539), .SDIN(n7266), .SSEL(test_se), .CLK(CK), .Q(n7267), .QN(n5782) );
  sdffs1 \DFF_615/Q_reg  ( .DIN(WX4537), .SDIN(n7265), .SSEL(test_se), .CLK(CK), .Q(n7266), .QN(n5787) );
  sdffs1 \DFF_614/Q_reg  ( .DIN(WX4535), .SDIN(n7264), .SSEL(test_se), .CLK(CK), .Q(n7265), .QN(n5792) );
  sdffs1 \DFF_613/Q_reg  ( .DIN(WX4533), .SDIN(n7263), .SSEL(test_se), .CLK(CK), .Q(n7264), .QN(n5797) );
  sdffs1 \DFF_612/Q_reg  ( .DIN(WX4531), .SDIN(n7262), .SSEL(test_se), .CLK(CK), .Q(n7263), .QN(n5802) );
  sdffs1 \DFF_611/Q_reg  ( .DIN(WX4529), .SDIN(n7261), .SSEL(test_se), .CLK(CK), .Q(n7262), .QN(n5807) );
  sdffs1 \DFF_610/Q_reg  ( .DIN(WX4527), .SDIN(n7260), .SSEL(test_se), .CLK(CK), .Q(n7261), .QN(n5812) );
  sdffs1 \DFF_609/Q_reg  ( .DIN(WX4525), .SDIN(n7259), .SSEL(test_se), .CLK(CK), .Q(n7260), .QN(n5817) );
  sdffs1 \DFF_608/Q_reg  ( .DIN(WX4523), .SDIN(n7258), .SSEL(test_se), .CLK(CK), .Q(n7259), .QN(n5822) );
  sdffs1 \DFF_607/Q_reg  ( .DIN(WX4425), .SDIN(n7257), .SSEL(test_se), .CLK(CK), .Q(n7258), .QN(n5652) );
  sdffs1 \DFF_606/Q_reg  ( .DIN(WX4423), .SDIN(n7256), .SSEL(test_se), .CLK(CK), .Q(n7257), .QN(n5653) );
  sdffs1 \DFF_605/Q_reg  ( .DIN(WX4421), .SDIN(n7255), .SSEL(test_se), .CLK(CK), .Q(n7256), .QN(n5654) );
  sdffs1 \DFF_604/Q_reg  ( .DIN(WX4419), .SDIN(n7254), .SSEL(test_se), .CLK(CK), .Q(n7255), .QN(n5655) );
  sdffs1 \DFF_603/Q_reg  ( .DIN(WX4417), .SDIN(n7253), .SSEL(test_se), .CLK(CK), .Q(n7254), .QN(n5656) );
  sdffs1 \DFF_602/Q_reg  ( .DIN(WX4415), .SDIN(n7252), .SSEL(test_se), .CLK(CK), .Q(n7253), .QN(n5657) );
  sdffs1 \DFF_601/Q_reg  ( .DIN(WX4413), .SDIN(n7251), .SSEL(test_se), .CLK(CK), .Q(n7252), .QN(n5658) );
  sdffs1 \DFF_600/Q_reg  ( .DIN(WX4411), .SDIN(n7250), .SSEL(test_se), .CLK(CK), .Q(n7251), .QN(n5659) );
  sdffs1 \DFF_599/Q_reg  ( .DIN(WX4409), .SDIN(n7249), .SSEL(test_se), .CLK(CK), .Q(n7250), .QN(n5660) );
  sdffs1 \DFF_598/Q_reg  ( .DIN(WX4407), .SDIN(n7248), .SSEL(test_se), .CLK(CK), .Q(n7249), .QN(n5661) );
  sdffs1 \DFF_597/Q_reg  ( .DIN(WX4405), .SDIN(n7247), .SSEL(test_se), .CLK(CK), .Q(n7248), .QN(n5662) );
  sdffs1 \DFF_596/Q_reg  ( .DIN(WX4403), .SDIN(n7246), .SSEL(test_se), .CLK(CK), .Q(n7247), .QN(n5663) );
  sdffs1 \DFF_595/Q_reg  ( .DIN(WX4401), .SDIN(n7245), .SSEL(test_se), .CLK(CK), .Q(n7246), .QN(n5664) );
  sdffs1 \DFF_594/Q_reg  ( .DIN(WX4399), .SDIN(n7244), .SSEL(test_se), .CLK(CK), .Q(n7245), .QN(n5665) );
  sdffs1 \DFF_593/Q_reg  ( .DIN(WX4397), .SDIN(n7243), .SSEL(test_se), .CLK(CK), .Q(n7244), .QN(n5666) );
  sdffs1 \DFF_592/Q_reg  ( .DIN(WX4395), .SDIN(n7242), .SSEL(test_se), .CLK(CK), .Q(n7243), .QN(n5667) );
  sdffs1 \DFF_591/Q_reg  ( .DIN(WX4393), .SDIN(n7241), .SSEL(test_se), .CLK(CK), .Q(n7242), .QN(n5668) );
  sdffs1 \DFF_590/Q_reg  ( .DIN(WX4391), .SDIN(n7240), .SSEL(test_se), .CLK(CK), .Q(n7241), .QN(n5669) );
  sdffs1 \DFF_589/Q_reg  ( .DIN(WX4389), .SDIN(n7239), .SSEL(test_se), .CLK(CK), .Q(n7240), .QN(n5670) );
  sdffs1 \DFF_588/Q_reg  ( .DIN(WX4387), .SDIN(n7238), .SSEL(test_se), .CLK(CK), .Q(n7239), .QN(n5671) );
  sdffs1 \DFF_587/Q_reg  ( .DIN(WX4385), .SDIN(n7237), .SSEL(test_se), .CLK(CK), .Q(n7238), .QN(n5672) );
  sdffs1 \DFF_586/Q_reg  ( .DIN(WX4383), .SDIN(n7236), .SSEL(test_se), .CLK(CK), .Q(n7237), .QN(n5673) );
  sdffs1 \DFF_585/Q_reg  ( .DIN(WX4381), .SDIN(n7235), .SSEL(test_se), .CLK(CK), .Q(n7236), .QN(n5674) );
  sdffs1 \DFF_584/Q_reg  ( .DIN(WX4379), .SDIN(n7234), .SSEL(test_se), .CLK(CK), .Q(n7235), .QN(n5675) );
  sdffs1 \DFF_583/Q_reg  ( .DIN(WX4377), .SDIN(n7233), .SSEL(test_se), .CLK(CK), .Q(n7234), .QN(n5676) );
  sdffs1 \DFF_582/Q_reg  ( .DIN(WX4375), .SDIN(n7232), .SSEL(test_se), .CLK(CK), .Q(n7233), .QN(n5677) );
  sdffs1 \DFF_581/Q_reg  ( .DIN(WX4373), .SDIN(n7231), .SSEL(test_se), .CLK(CK), .Q(n7232), .QN(n5678) );
  sdffs1 \DFF_580/Q_reg  ( .DIN(WX4371), .SDIN(n7230), .SSEL(test_se), .CLK(CK), .Q(n7231), .QN(n5679) );
  sdffs1 \DFF_579/Q_reg  ( .DIN(WX4369), .SDIN(n7229), .SSEL(test_se), .CLK(CK), .Q(n7230), .QN(n5680) );
  sdffs1 \DFF_578/Q_reg  ( .DIN(WX4367), .SDIN(n7228), .SSEL(test_se), .CLK(CK), .Q(n7229), .QN(n5681) );
  sdffs1 \DFF_577/Q_reg  ( .DIN(WX4365), .SDIN(n7227), .SSEL(test_se), .CLK(CK), .Q(n7228), .QN(n5682) );
  sdffs1 \DFF_576/Q_reg  ( .DIN(WX4363), .SDIN(CRC_OUT_7_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7227), .QN(n5651) );
  sdffs1 \DFF_575/Q_reg  ( .DIN(WX3912), .SDIN(CRC_OUT_7_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_31), .QN(n5826) );
  sdffs1 \DFF_574/Q_reg  ( .DIN(WX3910), .SDIN(CRC_OUT_7_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_30), .QN(n5821) );
  sdffs1 \DFF_573/Q_reg  ( .DIN(WX3908), .SDIN(CRC_OUT_7_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_29), .QN(n5816) );
  sdffs1 \DFF_572/Q_reg  ( .DIN(WX3906), .SDIN(CRC_OUT_7_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_28), .QN(n5811) );
  sdffs1 \DFF_571/Q_reg  ( .DIN(WX3904), .SDIN(CRC_OUT_7_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_27), .QN(n5806) );
  sdffs1 \DFF_570/Q_reg  ( .DIN(WX3902), .SDIN(CRC_OUT_7_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_26), .QN(n5801) );
  sdffs1 \DFF_569/Q_reg  ( .DIN(WX3900), .SDIN(CRC_OUT_7_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_25), .QN(n5796) );
  sdffs1 \DFF_568/Q_reg  ( .DIN(WX3898), .SDIN(CRC_OUT_7_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_24), .QN(n5791) );
  sdffs1 \DFF_567/Q_reg  ( .DIN(WX3896), .SDIN(CRC_OUT_7_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_23), .QN(n5786) );
  sdffs1 \DFF_566/Q_reg  ( .DIN(WX3894), .SDIN(CRC_OUT_7_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_22), .QN(n5781) );
  sdffs1 \DFF_565/Q_reg  ( .DIN(WX3892), .SDIN(CRC_OUT_7_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_21), .QN(n5776) );
  sdffs1 \DFF_564/Q_reg  ( .DIN(WX3890), .SDIN(CRC_OUT_7_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_20), .QN(n5771) );
  sdffs1 \DFF_563/Q_reg  ( .DIN(WX3888), .SDIN(CRC_OUT_7_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_19), .QN(n5766) );
  sdffs1 \DFF_562/Q_reg  ( .DIN(WX3886), .SDIN(CRC_OUT_7_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_18), .QN(n5761) );
  sdffs1 \DFF_561/Q_reg  ( .DIN(WX3884), .SDIN(CRC_OUT_7_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_17), .QN(n5756) );
  sdffs1 \DFF_560/Q_reg  ( .DIN(WX3882), .SDIN(CRC_OUT_7_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_16), .QN(n5751) );
  sdffs1 \DFF_559/Q_reg  ( .DIN(WX3880), .SDIN(CRC_OUT_7_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_15), .QN(n5746) );
  sdffs1 \DFF_558/Q_reg  ( .DIN(WX3878), .SDIN(CRC_OUT_7_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_14), .QN(n5742) );
  sdffs1 \DFF_557/Q_reg  ( .DIN(WX3876), .SDIN(CRC_OUT_7_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_13), .QN(n5738) );
  sdffs1 \DFF_556/Q_reg  ( .DIN(WX3874), .SDIN(CRC_OUT_7_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_12), .QN(n5734) );
  sdffs1 \DFF_555/Q_reg  ( .DIN(WX3872), .SDIN(CRC_OUT_7_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_11), .QN(n5730) );
  sdffs1 \DFF_554/Q_reg  ( .DIN(WX3870), .SDIN(CRC_OUT_7_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_10), .QN(n5726) );
  sdffs1 \DFF_553/Q_reg  ( .DIN(WX3868), .SDIN(CRC_OUT_7_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_9), .QN(n5722) );
  sdffs1 \DFF_552/Q_reg  ( .DIN(WX3866), .SDIN(CRC_OUT_7_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_8), .QN(n5718) );
  sdffs1 \DFF_551/Q_reg  ( .DIN(WX3864), .SDIN(CRC_OUT_7_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_7), .QN(n5714) );
  sdffs1 \DFF_550/Q_reg  ( .DIN(WX3862), .SDIN(CRC_OUT_7_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_6), .QN(n5710) );
  sdffs1 \DFF_549/Q_reg  ( .DIN(WX3860), .SDIN(CRC_OUT_7_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_5), .QN(n5706) );
  sdffs1 \DFF_548/Q_reg  ( .DIN(WX3858), .SDIN(CRC_OUT_7_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_4), .QN(n5702) );
  sdffs1 \DFF_547/Q_reg  ( .DIN(WX3856), .SDIN(CRC_OUT_7_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_3), .QN(n5698) );
  sdffs1 \DFF_546/Q_reg  ( .DIN(WX3854), .SDIN(CRC_OUT_7_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_2), .QN(n5694) );
  sdffs1 \DFF_545/Q_reg  ( .DIN(WX3852), .SDIN(CRC_OUT_7_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_7_1), .QN(n5690) );
  sdffs1 \DFF_544/Q_reg  ( .DIN(WX3850), .SDIN(n7226), .SSEL(test_se), .CLK(CK), .Q(CRC_OUT_7_0), .QN(n5686) );
  sdffs1 \DFF_543/Q_reg  ( .DIN(WX3484), .SDIN(n7225), .SSEL(test_se), .CLK(CK), .Q(n7226), .QN(n3285) );
  sdffs1 \DFF_542/Q_reg  ( .DIN(WX3482), .SDIN(n7224), .SSEL(test_se), .CLK(CK), .Q(n7225), .QN(n3287) );
  sdffs1 \DFF_541/Q_reg  ( .DIN(WX3480), .SDIN(n7223), .SSEL(test_se), .CLK(CK), .Q(n7224), .QN(n3289) );
  sdffs1 \DFF_540/Q_reg  ( .DIN(WX3478), .SDIN(n7222), .SSEL(test_se), .CLK(CK), .Q(n7223), .QN(n3291) );
  sdffs1 \DFF_539/Q_reg  ( .DIN(WX3476), .SDIN(n7221), .SSEL(test_se), .CLK(CK), .Q(n7222), .QN(n3293) );
  sdffs1 \DFF_538/Q_reg  ( .DIN(WX3474), .SDIN(n7220), .SSEL(test_se), .CLK(CK), .Q(n7221), .QN(n3295) );
  sdffs1 \DFF_537/Q_reg  ( .DIN(WX3472), .SDIN(n7219), .SSEL(test_se), .CLK(CK), .Q(n7220), .QN(n3297) );
  sdffs1 \DFF_536/Q_reg  ( .DIN(WX3470), .SDIN(n7218), .SSEL(test_se), .CLK(CK), .Q(n7219), .QN(n3299) );
  sdffs1 \DFF_535/Q_reg  ( .DIN(WX3468), .SDIN(n7217), .SSEL(test_se), .CLK(CK), .Q(n7218), .QN(n3301) );
  sdffs1 \DFF_534/Q_reg  ( .DIN(WX3466), .SDIN(n7216), .SSEL(test_se), .CLK(CK), .Q(n7217), .QN(n3303) );
  sdffs1 \DFF_533/Q_reg  ( .DIN(WX3464), .SDIN(n7215), .SSEL(test_se), .CLK(CK), .Q(n7216), .QN(n3305) );
  sdffs1 \DFF_532/Q_reg  ( .DIN(WX3462), .SDIN(n7214), .SSEL(test_se), .CLK(CK), .Q(n7215), .QN(n3307) );
  sdffs1 \DFF_531/Q_reg  ( .DIN(WX3460), .SDIN(n7213), .SSEL(test_se), .CLK(CK), .Q(n7214), .QN(n3309) );
  sdffs1 \DFF_530/Q_reg  ( .DIN(WX3458), .SDIN(n7212), .SSEL(test_se), .CLK(CK), .Q(n7213), .QN(n3311) );
  sdffs1 \DFF_529/Q_reg  ( .DIN(WX3456), .SDIN(n7211), .SSEL(test_se), .CLK(CK), .Q(n7212), .QN(n3313) );
  sdffs1 \DFF_528/Q_reg  ( .DIN(WX3454), .SDIN(n7210), .SSEL(test_se), .CLK(CK), .Q(n7211), .QN(n3315) );
  sdffs1 \DFF_527/Q_reg  ( .DIN(WX3452), .SDIN(n7209), .SSEL(test_se), .CLK(CK), .Q(n7210), .QN(n5974) );
  sdffs1 \DFF_526/Q_reg  ( .DIN(WX3450), .SDIN(n7208), .SSEL(test_se), .CLK(CK), .Q(n7209), .QN(n5983) );
  sdffs1 \DFF_525/Q_reg  ( .DIN(WX3448), .SDIN(n7207), .SSEL(test_se), .CLK(CK), .Q(n7208), .QN(n5992) );
  sdffs1 \DFF_524/Q_reg  ( .DIN(WX3446), .SDIN(n7206), .SSEL(test_se), .CLK(CK), .Q(n7207), .QN(n6001) );
  sdffs1 \DFF_523/Q_reg  ( .DIN(WX3444), .SDIN(n7205), .SSEL(test_se), .CLK(CK), .Q(n7206), .QN(n6010) );
  sdffs1 \DFF_522/Q_reg  ( .DIN(WX3442), .SDIN(n7204), .SSEL(test_se), .CLK(CK), .Q(n7205), .QN(n6019) );
  sdffs1 \DFF_521/Q_reg  ( .DIN(WX3440), .SDIN(n7203), .SSEL(test_se), .CLK(CK), .Q(n7204), .QN(n6028) );
  sdffs1 \DFF_520/Q_reg  ( .DIN(WX3438), .SDIN(n7202), .SSEL(test_se), .CLK(CK), .Q(n7203), .QN(n6037) );
  sdffs1 \DFF_519/Q_reg  ( .DIN(WX3436), .SDIN(n7201), .SSEL(test_se), .CLK(CK), .Q(n7202), .QN(n6046) );
  sdffs1 \DFF_518/Q_reg  ( .DIN(WX3434), .SDIN(n7200), .SSEL(test_se), .CLK(CK), .Q(n7201), .QN(n6055) );
  sdffs1 \DFF_517/Q_reg  ( .DIN(WX3432), .SDIN(n7199), .SSEL(test_se), .CLK(CK), .Q(n7200), .QN(n6064) );
  sdffs1 \DFF_516/Q_reg  ( .DIN(WX3430), .SDIN(n7198), .SSEL(test_se), .CLK(CK), .Q(n7199), .QN(n6073) );
  sdffs1 \DFF_515/Q_reg  ( .DIN(WX3428), .SDIN(n7197), .SSEL(test_se), .CLK(CK), .Q(n7198), .QN(n6082) );
  sdffs1 \DFF_514/Q_reg  ( .DIN(WX3426), .SDIN(n7196), .SSEL(test_se), .CLK(CK), .Q(n7197), .QN(n6091) );
  sdffs1 \DFF_513/Q_reg  ( .DIN(WX3424), .SDIN(n7195), .SSEL(test_se), .CLK(CK), .Q(n7196), .QN(n6100) );
  sdffs1 \DFF_512/Q_reg  ( .DIN(WX3422), .SDIN(n7194), .SSEL(test_se), .CLK(CK), .Q(n7195), .QN(n6109) );
  sdffs1 \DFF_511/Q_reg  ( .DIN(WX3420), .SDIN(n7193), .SSEL(test_se), .CLK(CK), .Q(n7194), .QN(n5861) );
  sdffs1 \DFF_510/Q_reg  ( .DIN(WX3418), .SDIN(n7192), .SSEL(test_se), .CLK(CK), .Q(n7193), .QN(n5868) );
  sdffs1 \DFF_509/Q_reg  ( .DIN(WX3416), .SDIN(n7191), .SSEL(test_se), .CLK(CK), .Q(n7192), .QN(n5875) );
  sdffs1 \DFF_508/Q_reg  ( .DIN(WX3414), .SDIN(n7190), .SSEL(test_se), .CLK(CK), .Q(n7191), .QN(n5882) );
  sdffs1 \DFF_507/Q_reg  ( .DIN(WX3412), .SDIN(n7189), .SSEL(test_se), .CLK(CK), .Q(n7190), .QN(n5889) );
  sdffs1 \DFF_506/Q_reg  ( .DIN(WX3410), .SDIN(n7188), .SSEL(test_se), .CLK(CK), .Q(n7189), .QN(n5896) );
  sdffs1 \DFF_505/Q_reg  ( .DIN(WX3408), .SDIN(n7187), .SSEL(test_se), .CLK(CK), .Q(n7188), .QN(n5903) );
  sdffs1 \DFF_504/Q_reg  ( .DIN(WX3406), .SDIN(n7186), .SSEL(test_se), .CLK(CK), .Q(n7187), .QN(n5910) );
  sdffs1 \DFF_503/Q_reg  ( .DIN(WX3404), .SDIN(n7185), .SSEL(test_se), .CLK(CK), .Q(n7186), .QN(n5917) );
  sdffs1 \DFF_502/Q_reg  ( .DIN(WX3402), .SDIN(n7184), .SSEL(test_se), .CLK(CK), .Q(n7185), .QN(n5924) );
  sdffs1 \DFF_501/Q_reg  ( .DIN(WX3400), .SDIN(n7183), .SSEL(test_se), .CLK(CK), .Q(n7184), .QN(n5931) );
  sdffs1 \DFF_500/Q_reg  ( .DIN(WX3398), .SDIN(n7182), .SSEL(test_se), .CLK(CK), .Q(n7183), .QN(n5938) );
  sdffs1 \DFF_499/Q_reg  ( .DIN(WX3396), .SDIN(n7181), .SSEL(test_se), .CLK(CK), .Q(n7182), .QN(n5945) );
  sdffs1 \DFF_498/Q_reg  ( .DIN(WX3394), .SDIN(n7180), .SSEL(test_se), .CLK(CK), .Q(n7181), .QN(n5952) );
  sdffs1 \DFF_497/Q_reg  ( .DIN(WX3392), .SDIN(n7179), .SSEL(test_se), .CLK(CK), .Q(n7180), .QN(n5959) );
  sdffs1 \DFF_496/Q_reg  ( .DIN(WX3390), .SDIN(n7178), .SSEL(test_se), .CLK(CK), .Q(n7179), .QN(n5966) );
  sdffs1 \DFF_495/Q_reg  ( .DIN(WX3388), .SDIN(n7177), .SSEL(test_se), .CLK(CK), .Q(n7178), .QN(n5973) );
  sdffs1 \DFF_494/Q_reg  ( .DIN(WX3386), .SDIN(n7176), .SSEL(test_se), .CLK(CK), .Q(n7177), .QN(n5982) );
  sdffs1 \DFF_493/Q_reg  ( .DIN(WX3384), .SDIN(n7175), .SSEL(test_se), .CLK(CK), .Q(n7176), .QN(n5991) );
  sdffs1 \DFF_492/Q_reg  ( .DIN(WX3382), .SDIN(n7174), .SSEL(test_se), .CLK(CK), .Q(n7175), .QN(n6000) );
  sdffs1 \DFF_491/Q_reg  ( .DIN(WX3380), .SDIN(n7173), .SSEL(test_se), .CLK(CK), .Q(n7174), .QN(n6009) );
  sdffs1 \DFF_490/Q_reg  ( .DIN(WX3378), .SDIN(n7172), .SSEL(test_se), .CLK(CK), .Q(n7173), .QN(n6018) );
  sdffs1 \DFF_489/Q_reg  ( .DIN(WX3376), .SDIN(n7171), .SSEL(test_se), .CLK(CK), .Q(n7172), .QN(n6027) );
  sdffs1 \DFF_488/Q_reg  ( .DIN(WX3374), .SDIN(n7170), .SSEL(test_se), .CLK(CK), .Q(n7171), .QN(n6036) );
  sdffs1 \DFF_487/Q_reg  ( .DIN(WX3372), .SDIN(n7169), .SSEL(test_se), .CLK(CK), .Q(n7170), .QN(n6045) );
  sdffs1 \DFF_486/Q_reg  ( .DIN(WX3370), .SDIN(n7168), .SSEL(test_se), .CLK(CK), .Q(n7169), .QN(n6054) );
  sdffs1 \DFF_485/Q_reg  ( .DIN(WX3368), .SDIN(n7167), .SSEL(test_se), .CLK(CK), .Q(n7168), .QN(n6063) );
  sdffs1 \DFF_484/Q_reg  ( .DIN(WX3366), .SDIN(n7166), .SSEL(test_se), .CLK(CK), .Q(n7167), .QN(n6072) );
  sdffs1 \DFF_483/Q_reg  ( .DIN(WX3364), .SDIN(n7165), .SSEL(test_se), .CLK(CK), .Q(n7166), .QN(n6081) );
  sdffs1 \DFF_482/Q_reg  ( .DIN(WX3362), .SDIN(n7164), .SSEL(test_se), .CLK(CK), .Q(n7165), .QN(n6090) );
  sdffs1 \DFF_481/Q_reg  ( .DIN(WX3360), .SDIN(n7163), .SSEL(test_se), .CLK(CK), .Q(n7164), .QN(n6099) );
  sdffs1 \DFF_480/Q_reg  ( .DIN(WX3358), .SDIN(n7162), .SSEL(test_se), .CLK(CK), .Q(n7163), .QN(n6108) );
  sdffs1 \DFF_479/Q_reg  ( .DIN(WX3356), .SDIN(n7161), .SSEL(test_se), .CLK(CK), .Q(n7162), .QN(n5860) );
  sdffs1 \DFF_478/Q_reg  ( .DIN(WX3354), .SDIN(n7160), .SSEL(test_se), .CLK(CK), .Q(n7161), .QN(n5867) );
  sdffs1 \DFF_477/Q_reg  ( .DIN(WX3352), .SDIN(n7159), .SSEL(test_se), .CLK(CK), .Q(n7160), .QN(n5874) );
  sdffs1 \DFF_476/Q_reg  ( .DIN(WX3350), .SDIN(n7158), .SSEL(test_se), .CLK(CK), .Q(n7159), .QN(n5881) );
  sdffs1 \DFF_475/Q_reg  ( .DIN(WX3348), .SDIN(n7157), .SSEL(test_se), .CLK(CK), .Q(n7158), .QN(n5888) );
  sdffs1 \DFF_474/Q_reg  ( .DIN(WX3346), .SDIN(n7156), .SSEL(test_se), .CLK(CK), .Q(n7157), .QN(n5895) );
  sdffs1 \DFF_473/Q_reg  ( .DIN(WX3344), .SDIN(n7155), .SSEL(test_se), .CLK(CK), .Q(n7156), .QN(n5902) );
  sdffs1 \DFF_472/Q_reg  ( .DIN(WX3342), .SDIN(n7154), .SSEL(test_se), .CLK(CK), .Q(n7155), .QN(n5909) );
  sdffs1 \DFF_471/Q_reg  ( .DIN(WX3340), .SDIN(n7153), .SSEL(test_se), .CLK(CK), .Q(n7154), .QN(n5916) );
  sdffs1 \DFF_470/Q_reg  ( .DIN(WX3338), .SDIN(n7152), .SSEL(test_se), .CLK(CK), .Q(n7153), .QN(n5923) );
  sdffs1 \DFF_469/Q_reg  ( .DIN(WX3336), .SDIN(n7151), .SSEL(test_se), .CLK(CK), .Q(n7152), .QN(n5930) );
  sdffs1 \DFF_468/Q_reg  ( .DIN(WX3334), .SDIN(n7150), .SSEL(test_se), .CLK(CK), .Q(n7151), .QN(n5937) );
  sdffs1 \DFF_467/Q_reg  ( .DIN(WX3332), .SDIN(n7149), .SSEL(test_se), .CLK(CK), .Q(n7150), .QN(n5944) );
  sdffs1 \DFF_466/Q_reg  ( .DIN(WX3330), .SDIN(n7148), .SSEL(test_se), .CLK(CK), .Q(n7149), .QN(n5951) );
  sdffs1 \DFF_465/Q_reg  ( .DIN(WX3328), .SDIN(n7147), .SSEL(test_se), .CLK(CK), .Q(n7148), .QN(n5958) );
  sdffs1 \DFF_464/Q_reg  ( .DIN(WX3326), .SDIN(n5972), .SSEL(test_se), .CLK(CK), .Q(n7147), .QN(n5965) );
  sdffs1 \DFF_463/Q_reg  ( .DIN(WX3324), .SDIN(n5981), .SSEL(test_se), .CLK(CK), .Q(n5972) );
  sdffs1 \DFF_462/Q_reg  ( .DIN(WX3322), .SDIN(n5990), .SSEL(test_se), .CLK(CK), .Q(n5981) );
  sdffs1 \DFF_461/Q_reg  ( .DIN(WX3320), .SDIN(n5999), .SSEL(test_se), .CLK(CK), .Q(n5990) );
  sdffs1 \DFF_460/Q_reg  ( .DIN(WX3318), .SDIN(n6008), .SSEL(test_se), .CLK(CK), .Q(n5999) );
  sdffs1 \DFF_459/Q_reg  ( .DIN(WX3316), .SDIN(n6017), .SSEL(test_se), .CLK(CK), .Q(n6008) );
  sdffs1 \DFF_458/Q_reg  ( .DIN(WX3314), .SDIN(n6026), .SSEL(test_se), .CLK(CK), .Q(n6017) );
  sdffs1 \DFF_457/Q_reg  ( .DIN(WX3312), .SDIN(n6035), .SSEL(test_se), .CLK(CK), .Q(n6026) );
  sdffs1 \DFF_456/Q_reg  ( .DIN(WX3310), .SDIN(n6044), .SSEL(test_se), .CLK(CK), .Q(n6035) );
  sdffs1 \DFF_455/Q_reg  ( .DIN(WX3308), .SDIN(n6053), .SSEL(test_se), .CLK(CK), .Q(n6044) );
  sdffs1 \DFF_454/Q_reg  ( .DIN(WX3306), .SDIN(n6062), .SSEL(test_se), .CLK(CK), .Q(n6053) );
  sdffs1 \DFF_453/Q_reg  ( .DIN(WX3304), .SDIN(n6071), .SSEL(test_se), .CLK(CK), .Q(n6062) );
  sdffs1 \DFF_452/Q_reg  ( .DIN(WX3302), .SDIN(n6080), .SSEL(test_se), .CLK(CK), .Q(n6071) );
  sdffs1 \DFF_451/Q_reg  ( .DIN(WX3300), .SDIN(n6089), .SSEL(test_se), .CLK(CK), .Q(n6080) );
  sdffs1 \DFF_450/Q_reg  ( .DIN(WX3298), .SDIN(n6098), .SSEL(test_se), .CLK(CK), .Q(n6089) );
  sdffs1 \DFF_449/Q_reg  ( .DIN(WX3296), .SDIN(n6107), .SSEL(test_se), .CLK(CK), .Q(n6098) );
  sdffs1 \DFF_448/Q_reg  ( .DIN(WX3294), .SDIN(n5859), .SSEL(test_se), .CLK(CK), .Q(n6107) );
  sdffs1 \DFF_447/Q_reg  ( .DIN(WX3292), .SDIN(n5866), .SSEL(test_se), .CLK(CK), .Q(n5859) );
  sdffs1 \DFF_446/Q_reg  ( .DIN(WX3290), .SDIN(n5873), .SSEL(test_se), .CLK(CK), .Q(n5866) );
  sdffs1 \DFF_445/Q_reg  ( .DIN(WX3288), .SDIN(n5880), .SSEL(test_se), .CLK(CK), .Q(n5873) );
  sdffs1 \DFF_444/Q_reg  ( .DIN(WX3286), .SDIN(n5887), .SSEL(test_se), .CLK(CK), .Q(n5880) );
  sdffs1 \DFF_443/Q_reg  ( .DIN(WX3284), .SDIN(n5894), .SSEL(test_se), .CLK(CK), .Q(n5887) );
  sdffs1 \DFF_442/Q_reg  ( .DIN(WX3282), .SDIN(n5901), .SSEL(test_se), .CLK(CK), .Q(n5894) );
  sdffs1 \DFF_441/Q_reg  ( .DIN(WX3280), .SDIN(n5908), .SSEL(test_se), .CLK(CK), .Q(n5901) );
  sdffs1 \DFF_440/Q_reg  ( .DIN(WX3278), .SDIN(n5915), .SSEL(test_se), .CLK(CK), .Q(n5908) );
  sdffs1 \DFF_439/Q_reg  ( .DIN(WX3276), .SDIN(n5922), .SSEL(test_se), .CLK(CK), .Q(n5915) );
  sdffs1 \DFF_438/Q_reg  ( .DIN(WX3274), .SDIN(n5929), .SSEL(test_se), .CLK(CK), .Q(n5922) );
  sdffs1 \DFF_437/Q_reg  ( .DIN(WX3272), .SDIN(n5936), .SSEL(test_se), .CLK(CK), .Q(n5929) );
  sdffs1 \DFF_436/Q_reg  ( .DIN(WX3270), .SDIN(n5943), .SSEL(test_se), .CLK(CK), .Q(n5936) );
  sdffs1 \DFF_435/Q_reg  ( .DIN(WX3268), .SDIN(n5950), .SSEL(test_se), .CLK(CK), .Q(n5943) );
  sdffs1 \DFF_434/Q_reg  ( .DIN(WX3266), .SDIN(n5957), .SSEL(test_se), .CLK(CK), .Q(n5950) );
  sdffs1 \DFF_433/Q_reg  ( .DIN(WX3264), .SDIN(n5964), .SSEL(test_se), .CLK(CK), .Q(n5957) );
  sdffs1 \DFF_432/Q_reg  ( .DIN(WX3262), .SDIN(n7146), .SSEL(test_se), .CLK(CK), .Q(n5964) );
  sdffs1 \DFF_431/Q_reg  ( .DIN(WX3260), .SDIN(n7145), .SSEL(test_se), .CLK(CK), .Q(n7146), .QN(n5971) );
  sdffs1 \DFF_430/Q_reg  ( .DIN(WX3258), .SDIN(n7144), .SSEL(test_se), .CLK(CK), .Q(n7145), .QN(n5980) );
  sdffs1 \DFF_429/Q_reg  ( .DIN(WX3256), .SDIN(n7143), .SSEL(test_se), .CLK(CK), .Q(n7144), .QN(n5989) );
  sdffs1 \DFF_428/Q_reg  ( .DIN(WX3254), .SDIN(n7142), .SSEL(test_se), .CLK(CK), .Q(n7143), .QN(n5998) );
  sdffs1 \DFF_427/Q_reg  ( .DIN(WX3252), .SDIN(n7141), .SSEL(test_se), .CLK(CK), .Q(n7142), .QN(n6007) );
  sdffs1 \DFF_426/Q_reg  ( .DIN(WX3250), .SDIN(n7140), .SSEL(test_se), .CLK(CK), .Q(n7141), .QN(n6016) );
  sdffs1 \DFF_425/Q_reg  ( .DIN(WX3248), .SDIN(n7139), .SSEL(test_se), .CLK(CK), .Q(n7140), .QN(n6025) );
  sdffs1 \DFF_424/Q_reg  ( .DIN(WX3246), .SDIN(n7138), .SSEL(test_se), .CLK(CK), .Q(n7139), .QN(n6034) );
  sdffs1 \DFF_423/Q_reg  ( .DIN(WX3244), .SDIN(n7137), .SSEL(test_se), .CLK(CK), .Q(n7138), .QN(n6043) );
  sdffs1 \DFF_422/Q_reg  ( .DIN(WX3242), .SDIN(n7136), .SSEL(test_se), .CLK(CK), .Q(n7137), .QN(n6052) );
  sdffs1 \DFF_421/Q_reg  ( .DIN(WX3240), .SDIN(n7135), .SSEL(test_se), .CLK(CK), .Q(n7136), .QN(n6061) );
  sdffs1 \DFF_420/Q_reg  ( .DIN(WX3238), .SDIN(n7134), .SSEL(test_se), .CLK(CK), .Q(n7135), .QN(n6070) );
  sdffs1 \DFF_419/Q_reg  ( .DIN(WX3236), .SDIN(n7133), .SSEL(test_se), .CLK(CK), .Q(n7134), .QN(n6079) );
  sdffs1 \DFF_418/Q_reg  ( .DIN(WX3234), .SDIN(n7132), .SSEL(test_se), .CLK(CK), .Q(n7133), .QN(n6088) );
  sdffs1 \DFF_417/Q_reg  ( .DIN(WX3232), .SDIN(n7131), .SSEL(test_se), .CLK(CK), .Q(n7132), .QN(n6097) );
  sdffs1 \DFF_416/Q_reg  ( .DIN(WX3230), .SDIN(n7130), .SSEL(test_se), .CLK(CK), .Q(n7131), .QN(n6106) );
  sdffs1 \DFF_415/Q_reg  ( .DIN(WX3132), .SDIN(n7129), .SSEL(test_se), .CLK(CK), .Q(n7130), .QN(n5828) );
  sdffs1 \DFF_414/Q_reg  ( .DIN(WX3130), .SDIN(n7128), .SSEL(test_se), .CLK(CK), .Q(n7129), .QN(n5829) );
  sdffs1 \DFF_413/Q_reg  ( .DIN(WX3128), .SDIN(n7127), .SSEL(test_se), .CLK(CK), .Q(n7128), .QN(n5830) );
  sdffs1 \DFF_412/Q_reg  ( .DIN(WX3126), .SDIN(n7126), .SSEL(test_se), .CLK(CK), .Q(n7127), .QN(n5831) );
  sdffs1 \DFF_411/Q_reg  ( .DIN(WX3124), .SDIN(n7125), .SSEL(test_se), .CLK(CK), .Q(n7126), .QN(n5832) );
  sdffs1 \DFF_410/Q_reg  ( .DIN(WX3122), .SDIN(n7124), .SSEL(test_se), .CLK(CK), .Q(n7125), .QN(n5833) );
  sdffs1 \DFF_409/Q_reg  ( .DIN(WX3120), .SDIN(n7123), .SSEL(test_se), .CLK(CK), .Q(n7124), .QN(n5834) );
  sdffs1 \DFF_408/Q_reg  ( .DIN(WX3118), .SDIN(n7122), .SSEL(test_se), .CLK(CK), .Q(n7123), .QN(n5835) );
  sdffs1 \DFF_407/Q_reg  ( .DIN(WX3116), .SDIN(n7121), .SSEL(test_se), .CLK(CK), .Q(n7122), .QN(n5836) );
  sdffs1 \DFF_406/Q_reg  ( .DIN(WX3114), .SDIN(n7120), .SSEL(test_se), .CLK(CK), .Q(n7121), .QN(n5837) );
  sdffs1 \DFF_405/Q_reg  ( .DIN(WX3112), .SDIN(n7119), .SSEL(test_se), .CLK(CK), .Q(n7120), .QN(n5838) );
  sdffs1 \DFF_404/Q_reg  ( .DIN(WX3110), .SDIN(n7118), .SSEL(test_se), .CLK(CK), .Q(n7119), .QN(n5839) );
  sdffs1 \DFF_403/Q_reg  ( .DIN(WX3108), .SDIN(n7117), .SSEL(test_se), .CLK(CK), .Q(n7118), .QN(n5840) );
  sdffs1 \DFF_402/Q_reg  ( .DIN(WX3106), .SDIN(n7116), .SSEL(test_se), .CLK(CK), .Q(n7117), .QN(n5841) );
  sdffs1 \DFF_401/Q_reg  ( .DIN(WX3104), .SDIN(n7115), .SSEL(test_se), .CLK(CK), .Q(n7116), .QN(n5842) );
  sdffs1 \DFF_400/Q_reg  ( .DIN(WX3102), .SDIN(n7114), .SSEL(test_se), .CLK(CK), .Q(n7115), .QN(n5843) );
  sdffs1 \DFF_399/Q_reg  ( .DIN(WX3100), .SDIN(n7113), .SSEL(test_se), .CLK(CK), .Q(n7114), .QN(n5844) );
  sdffs1 \DFF_398/Q_reg  ( .DIN(WX3098), .SDIN(n7112), .SSEL(test_se), .CLK(CK), .Q(n7113), .QN(n5845) );
  sdffs1 \DFF_397/Q_reg  ( .DIN(WX3096), .SDIN(n7111), .SSEL(test_se), .CLK(CK), .Q(n7112), .QN(n5846) );
  sdffs1 \DFF_396/Q_reg  ( .DIN(WX3094), .SDIN(n7110), .SSEL(test_se), .CLK(CK), .Q(n7111), .QN(n5847) );
  sdffs1 \DFF_395/Q_reg  ( .DIN(WX3092), .SDIN(n7109), .SSEL(test_se), .CLK(CK), .Q(n7110), .QN(n5848) );
  sdffs1 \DFF_394/Q_reg  ( .DIN(WX3090), .SDIN(n7108), .SSEL(test_se), .CLK(CK), .Q(n7109), .QN(n5849) );
  sdffs1 \DFF_393/Q_reg  ( .DIN(WX3088), .SDIN(n7107), .SSEL(test_se), .CLK(CK), .Q(n7108), .QN(n5850) );
  sdffs1 \DFF_392/Q_reg  ( .DIN(WX3086), .SDIN(n7106), .SSEL(test_se), .CLK(CK), .Q(n7107), .QN(n5851) );
  sdffs1 \DFF_391/Q_reg  ( .DIN(WX3084), .SDIN(n7105), .SSEL(test_se), .CLK(CK), .Q(n7106), .QN(n5852) );
  sdffs1 \DFF_390/Q_reg  ( .DIN(WX3082), .SDIN(n7104), .SSEL(test_se), .CLK(CK), .Q(n7105), .QN(n5853) );
  sdffs1 \DFF_389/Q_reg  ( .DIN(WX3080), .SDIN(n7103), .SSEL(test_se), .CLK(CK), .Q(n7104), .QN(n5854) );
  sdffs1 \DFF_388/Q_reg  ( .DIN(WX3078), .SDIN(n7102), .SSEL(test_se), .CLK(CK), .Q(n7103), .QN(n5855) );
  sdffs1 \DFF_387/Q_reg  ( .DIN(WX3076), .SDIN(n7101), .SSEL(test_se), .CLK(CK), .Q(n7102), .QN(n5856) );
  sdffs1 \DFF_386/Q_reg  ( .DIN(WX3074), .SDIN(n7100), .SSEL(test_se), .CLK(CK), .Q(n7101), .QN(n5857) );
  sdffs1 \DFF_385/Q_reg  ( .DIN(WX3072), .SDIN(n7099), .SSEL(test_se), .CLK(CK), .Q(n7100), .QN(n5858) );
  sdffs1 \DFF_384/Q_reg  ( .DIN(WX3070), .SDIN(CRC_OUT_8_31), .SSEL(test_se), 
        .CLK(CK), .Q(n7099), .QN(n5827) );
  sdffs1 \DFF_383/Q_reg  ( .DIN(WX2619), .SDIN(CRC_OUT_8_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_31), .QN(n6114) );
  sdffs1 \DFF_382/Q_reg  ( .DIN(WX2617), .SDIN(CRC_OUT_8_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_30), .QN(n6105) );
  sdffs1 \DFF_381/Q_reg  ( .DIN(WX2615), .SDIN(CRC_OUT_8_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_29), .QN(n6096) );
  sdffs1 \DFF_380/Q_reg  ( .DIN(WX2613), .SDIN(CRC_OUT_8_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_28), .QN(n6087) );
  sdffs1 \DFF_379/Q_reg  ( .DIN(WX2611), .SDIN(CRC_OUT_8_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_27), .QN(n6078) );
  sdffs1 \DFF_378/Q_reg  ( .DIN(WX2609), .SDIN(CRC_OUT_8_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_26), .QN(n6069) );
  sdffs1 \DFF_377/Q_reg  ( .DIN(WX2607), .SDIN(CRC_OUT_8_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_25), .QN(n6060) );
  sdffs1 \DFF_376/Q_reg  ( .DIN(WX2605), .SDIN(CRC_OUT_8_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_24), .QN(n6051) );
  sdffs1 \DFF_375/Q_reg  ( .DIN(WX2603), .SDIN(CRC_OUT_8_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_23), .QN(n6042) );
  sdffs1 \DFF_374/Q_reg  ( .DIN(WX2601), .SDIN(CRC_OUT_8_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_22), .QN(n6033) );
  sdffs1 \DFF_373/Q_reg  ( .DIN(WX2599), .SDIN(CRC_OUT_8_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_21), .QN(n6024) );
  sdffs1 \DFF_372/Q_reg  ( .DIN(WX2597), .SDIN(CRC_OUT_8_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_20), .QN(n6015) );
  sdffs1 \DFF_371/Q_reg  ( .DIN(WX2595), .SDIN(CRC_OUT_8_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_19), .QN(n6006) );
  sdffs1 \DFF_370/Q_reg  ( .DIN(WX2593), .SDIN(CRC_OUT_8_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_18), .QN(n5997) );
  sdffs1 \DFF_369/Q_reg  ( .DIN(WX2591), .SDIN(CRC_OUT_8_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_17), .QN(n5988) );
  sdffs1 \DFF_368/Q_reg  ( .DIN(WX2589), .SDIN(CRC_OUT_8_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_16), .QN(n5979) );
  sdffs1 \DFF_367/Q_reg  ( .DIN(WX2587), .SDIN(CRC_OUT_8_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_15), .QN(n5970) );
  sdffs1 \DFF_366/Q_reg  ( .DIN(WX2585), .SDIN(CRC_OUT_8_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_14), .QN(n5963) );
  sdffs1 \DFF_365/Q_reg  ( .DIN(WX2583), .SDIN(CRC_OUT_8_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_13), .QN(n5956) );
  sdffs1 \DFF_364/Q_reg  ( .DIN(WX2581), .SDIN(CRC_OUT_8_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_12), .QN(n5949) );
  sdffs1 \DFF_363/Q_reg  ( .DIN(WX2579), .SDIN(CRC_OUT_8_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_11), .QN(n5942) );
  sdffs1 \DFF_362/Q_reg  ( .DIN(WX2577), .SDIN(CRC_OUT_8_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_10), .QN(n5935) );
  sdffs1 \DFF_361/Q_reg  ( .DIN(WX2575), .SDIN(CRC_OUT_8_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_9), .QN(n5928) );
  sdffs1 \DFF_360/Q_reg  ( .DIN(WX2573), .SDIN(CRC_OUT_8_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_8), .QN(n5921) );
  sdffs1 \DFF_359/Q_reg  ( .DIN(WX2571), .SDIN(CRC_OUT_8_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_7), .QN(n5914) );
  sdffs1 \DFF_358/Q_reg  ( .DIN(WX2569), .SDIN(CRC_OUT_8_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_6), .QN(n5907) );
  sdffs1 \DFF_357/Q_reg  ( .DIN(WX2567), .SDIN(CRC_OUT_8_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_5), .QN(n5900) );
  sdffs1 \DFF_356/Q_reg  ( .DIN(WX2565), .SDIN(CRC_OUT_8_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_4), .QN(n5893) );
  sdffs1 \DFF_355/Q_reg  ( .DIN(WX2563), .SDIN(CRC_OUT_8_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_3), .QN(n5886) );
  sdffs1 \DFF_354/Q_reg  ( .DIN(WX2561), .SDIN(CRC_OUT_8_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_2), .QN(n5879) );
  sdffs1 \DFF_353/Q_reg  ( .DIN(WX2559), .SDIN(CRC_OUT_8_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_8_1), .QN(n5872) );
  sdffs1 \DFF_352/Q_reg  ( .DIN(WX2557), .SDIN(n7098), .SSEL(test_se), .CLK(CK), .Q(CRC_OUT_8_0), .QN(n5865) );
  sdffs1 \DFF_351/Q_reg  ( .DIN(WX2191), .SDIN(n7097), .SSEL(test_se), .CLK(CK), .Q(n7098), .QN(n3286) );
  sdffs1 \DFF_350/Q_reg  ( .DIN(WX2189), .SDIN(n7096), .SSEL(test_se), .CLK(CK), .Q(n7097), .QN(n3288) );
  sdffs1 \DFF_349/Q_reg  ( .DIN(WX2187), .SDIN(n7095), .SSEL(test_se), .CLK(CK), .Q(n7096), .QN(n3290) );
  sdffs1 \DFF_348/Q_reg  ( .DIN(WX2185), .SDIN(n7094), .SSEL(test_se), .CLK(CK), .Q(n7095), .QN(n3292) );
  sdffs1 \DFF_347/Q_reg  ( .DIN(WX2183), .SDIN(n7093), .SSEL(test_se), .CLK(CK), .Q(n7094), .QN(n3294) );
  sdffs1 \DFF_346/Q_reg  ( .DIN(WX2181), .SDIN(n7092), .SSEL(test_se), .CLK(CK), .Q(n7093), .QN(n3296) );
  sdffs1 \DFF_345/Q_reg  ( .DIN(WX2179), .SDIN(n7091), .SSEL(test_se), .CLK(CK), .Q(n7092), .QN(n3298) );
  sdffs1 \DFF_344/Q_reg  ( .DIN(WX2177), .SDIN(n7090), .SSEL(test_se), .CLK(CK), .Q(n7091), .QN(n3300) );
  sdffs1 \DFF_343/Q_reg  ( .DIN(WX2175), .SDIN(n7089), .SSEL(test_se), .CLK(CK), .Q(n7090), .QN(n3302) );
  sdffs1 \DFF_342/Q_reg  ( .DIN(WX2173), .SDIN(n7088), .SSEL(test_se), .CLK(CK), .Q(n7089), .QN(n3304) );
  sdffs1 \DFF_341/Q_reg  ( .DIN(WX2171), .SDIN(n7087), .SSEL(test_se), .CLK(CK), .Q(n7088), .QN(n3306) );
  sdffs1 \DFF_340/Q_reg  ( .DIN(WX2169), .SDIN(n7086), .SSEL(test_se), .CLK(CK), .Q(n7087), .QN(n3308) );
  sdffs1 \DFF_339/Q_reg  ( .DIN(WX2167), .SDIN(n7085), .SSEL(test_se), .CLK(CK), .Q(n7086), .QN(n3310) );
  sdffs1 \DFF_338/Q_reg  ( .DIN(WX2165), .SDIN(n7084), .SSEL(test_se), .CLK(CK), .Q(n7085), .QN(n3312) );
  sdffs1 \DFF_337/Q_reg  ( .DIN(WX2163), .SDIN(n7083), .SSEL(test_se), .CLK(CK), .Q(n7084), .QN(n3314) );
  sdffs1 \DFF_336/Q_reg  ( .DIN(WX2161), .SDIN(n7082), .SSEL(test_se), .CLK(CK), .Q(n7083), .QN(n3316) );
  sdffs1 \DFF_335/Q_reg  ( .DIN(WX2159), .SDIN(n7081), .SSEL(test_se), .CLK(CK), .Q(n7082), .QN(n5978) );
  sdffs1 \DFF_334/Q_reg  ( .DIN(WX2157), .SDIN(n7080), .SSEL(test_se), .CLK(CK), .Q(n7081), .QN(n5987) );
  sdffs1 \DFF_333/Q_reg  ( .DIN(WX2155), .SDIN(n7079), .SSEL(test_se), .CLK(CK), .Q(n7080), .QN(n5996) );
  sdffs1 \DFF_332/Q_reg  ( .DIN(WX2153), .SDIN(n7078), .SSEL(test_se), .CLK(CK), .Q(n7079), .QN(n6005) );
  sdffs1 \DFF_331/Q_reg  ( .DIN(WX2151), .SDIN(n7077), .SSEL(test_se), .CLK(CK), .Q(n7078), .QN(n6014) );
  sdffs1 \DFF_330/Q_reg  ( .DIN(WX2149), .SDIN(n7076), .SSEL(test_se), .CLK(CK), .Q(n7077), .QN(n6023) );
  sdffs1 \DFF_329/Q_reg  ( .DIN(WX2147), .SDIN(n7075), .SSEL(test_se), .CLK(CK), .Q(n7076), .QN(n6032) );
  sdffs1 \DFF_328/Q_reg  ( .DIN(WX2145), .SDIN(n7074), .SSEL(test_se), .CLK(CK), .Q(n7075), .QN(n6041) );
  sdffs1 \DFF_327/Q_reg  ( .DIN(WX2143), .SDIN(n7073), .SSEL(test_se), .CLK(CK), .Q(n7074), .QN(n6050) );
  sdffs1 \DFF_326/Q_reg  ( .DIN(WX2141), .SDIN(n7072), .SSEL(test_se), .CLK(CK), .Q(n7073), .QN(n6059) );
  sdffs1 \DFF_325/Q_reg  ( .DIN(WX2139), .SDIN(n7071), .SSEL(test_se), .CLK(CK), .Q(n7072), .QN(n6068) );
  sdffs1 \DFF_324/Q_reg  ( .DIN(WX2137), .SDIN(n7070), .SSEL(test_se), .CLK(CK), .Q(n7071), .QN(n6077) );
  sdffs1 \DFF_323/Q_reg  ( .DIN(WX2135), .SDIN(n7069), .SSEL(test_se), .CLK(CK), .Q(n7070), .QN(n6086) );
  sdffs1 \DFF_322/Q_reg  ( .DIN(WX2133), .SDIN(n7068), .SSEL(test_se), .CLK(CK), .Q(n7069), .QN(n6095) );
  sdffs1 \DFF_321/Q_reg  ( .DIN(WX2131), .SDIN(n7067), .SSEL(test_se), .CLK(CK), .Q(n7068), .QN(n6104) );
  sdffs1 \DFF_320/Q_reg  ( .DIN(WX2129), .SDIN(n7066), .SSEL(test_se), .CLK(CK), .Q(n7067), .QN(n6113) );
  sdffs1 \DFF_319/Q_reg  ( .DIN(WX2127), .SDIN(n7065), .SSEL(test_se), .CLK(CK), .Q(n7066), .QN(n5864) );
  sdffs1 \DFF_318/Q_reg  ( .DIN(WX2125), .SDIN(n7064), .SSEL(test_se), .CLK(CK), .Q(n7065), .QN(n5871) );
  sdffs1 \DFF_317/Q_reg  ( .DIN(WX2123), .SDIN(n7063), .SSEL(test_se), .CLK(CK), .Q(n7064), .QN(n5878) );
  sdffs1 \DFF_316/Q_reg  ( .DIN(WX2121), .SDIN(n7062), .SSEL(test_se), .CLK(CK), .Q(n7063), .QN(n5885) );
  sdffs1 \DFF_315/Q_reg  ( .DIN(WX2119), .SDIN(n7061), .SSEL(test_se), .CLK(CK), .Q(n7062), .QN(n5892) );
  sdffs1 \DFF_314/Q_reg  ( .DIN(WX2117), .SDIN(n7060), .SSEL(test_se), .CLK(CK), .Q(n7061), .QN(n5899) );
  sdffs1 \DFF_313/Q_reg  ( .DIN(WX2115), .SDIN(n7059), .SSEL(test_se), .CLK(CK), .Q(n7060), .QN(n5906) );
  sdffs1 \DFF_312/Q_reg  ( .DIN(WX2113), .SDIN(n7058), .SSEL(test_se), .CLK(CK), .Q(n7059), .QN(n5913) );
  sdffs1 \DFF_311/Q_reg  ( .DIN(WX2111), .SDIN(n7057), .SSEL(test_se), .CLK(CK), .Q(n7058), .QN(n5920) );
  sdffs1 \DFF_310/Q_reg  ( .DIN(WX2109), .SDIN(n7056), .SSEL(test_se), .CLK(CK), .Q(n7057), .QN(n5927) );
  sdffs1 \DFF_309/Q_reg  ( .DIN(WX2107), .SDIN(n7055), .SSEL(test_se), .CLK(CK), .Q(n7056), .QN(n5934) );
  sdffs1 \DFF_308/Q_reg  ( .DIN(WX2105), .SDIN(n7054), .SSEL(test_se), .CLK(CK), .Q(n7055), .QN(n5941) );
  sdffs1 \DFF_307/Q_reg  ( .DIN(WX2103), .SDIN(n7053), .SSEL(test_se), .CLK(CK), .Q(n7054), .QN(n5948) );
  sdffs1 \DFF_306/Q_reg  ( .DIN(WX2101), .SDIN(n7052), .SSEL(test_se), .CLK(CK), .Q(n7053), .QN(n5955) );
  sdffs1 \DFF_305/Q_reg  ( .DIN(WX2099), .SDIN(n7051), .SSEL(test_se), .CLK(CK), .Q(n7052), .QN(n5962) );
  sdffs1 \DFF_304/Q_reg  ( .DIN(WX2097), .SDIN(n7050), .SSEL(test_se), .CLK(CK), .Q(n7051), .QN(n5969) );
  sdffs1 \DFF_303/Q_reg  ( .DIN(WX2095), .SDIN(n7049), .SSEL(test_se), .CLK(CK), .Q(n7050), .QN(n5977) );
  sdffs1 \DFF_302/Q_reg  ( .DIN(WX2093), .SDIN(n7048), .SSEL(test_se), .CLK(CK), .Q(n7049), .QN(n5986) );
  sdffs1 \DFF_301/Q_reg  ( .DIN(WX2091), .SDIN(n7047), .SSEL(test_se), .CLK(CK), .Q(n7048), .QN(n5995) );
  sdffs1 \DFF_300/Q_reg  ( .DIN(WX2089), .SDIN(n7046), .SSEL(test_se), .CLK(CK), .Q(n7047), .QN(n6004) );
  sdffs1 \DFF_299/Q_reg  ( .DIN(WX2087), .SDIN(n7045), .SSEL(test_se), .CLK(CK), .Q(n7046), .QN(n6013) );
  sdffs1 \DFF_298/Q_reg  ( .DIN(WX2085), .SDIN(n7044), .SSEL(test_se), .CLK(CK), .Q(n7045), .QN(n6022) );
  sdffs1 \DFF_297/Q_reg  ( .DIN(WX2083), .SDIN(n7043), .SSEL(test_se), .CLK(CK), .Q(n7044), .QN(n6031) );
  sdffs1 \DFF_296/Q_reg  ( .DIN(WX2081), .SDIN(n7042), .SSEL(test_se), .CLK(CK), .Q(n7043), .QN(n6040) );
  sdffs1 \DFF_295/Q_reg  ( .DIN(WX2079), .SDIN(n7041), .SSEL(test_se), .CLK(CK), .Q(n7042), .QN(n6049) );
  sdffs1 \DFF_294/Q_reg  ( .DIN(WX2077), .SDIN(n7040), .SSEL(test_se), .CLK(CK), .Q(n7041), .QN(n6058) );
  sdffs1 \DFF_293/Q_reg  ( .DIN(WX2075), .SDIN(n7039), .SSEL(test_se), .CLK(CK), .Q(n7040), .QN(n6067) );
  sdffs1 \DFF_292/Q_reg  ( .DIN(WX2073), .SDIN(n7038), .SSEL(test_se), .CLK(CK), .Q(n7039), .QN(n6076) );
  sdffs1 \DFF_291/Q_reg  ( .DIN(WX2071), .SDIN(n7037), .SSEL(test_se), .CLK(CK), .Q(n7038), .QN(n6085) );
  sdffs1 \DFF_290/Q_reg  ( .DIN(WX2069), .SDIN(n7036), .SSEL(test_se), .CLK(CK), .Q(n7037), .QN(n6094) );
  sdffs1 \DFF_289/Q_reg  ( .DIN(WX2067), .SDIN(n7035), .SSEL(test_se), .CLK(CK), .Q(n7036), .QN(n6103) );
  sdffs1 \DFF_288/Q_reg  ( .DIN(WX2065), .SDIN(n5863), .SSEL(test_se), .CLK(CK), .Q(n7035), .QN(n6112) );
  sdffs1 \DFF_287/Q_reg  ( .DIN(WX2063), .SDIN(n5870), .SSEL(test_se), .CLK(CK), .Q(n5863) );
  sdffs1 \DFF_286/Q_reg  ( .DIN(WX2061), .SDIN(n5877), .SSEL(test_se), .CLK(CK), .Q(n5870) );
  sdffs1 \DFF_285/Q_reg  ( .DIN(WX2059), .SDIN(n5884), .SSEL(test_se), .CLK(CK), .Q(n5877) );
  sdffs1 \DFF_284/Q_reg  ( .DIN(WX2057), .SDIN(n5891), .SSEL(test_se), .CLK(CK), .Q(n5884) );
  sdffs1 \DFF_283/Q_reg  ( .DIN(WX2055), .SDIN(n5898), .SSEL(test_se), .CLK(CK), .Q(n5891) );
  sdffs1 \DFF_282/Q_reg  ( .DIN(WX2053), .SDIN(n5905), .SSEL(test_se), .CLK(CK), .Q(n5898) );
  sdffs1 \DFF_281/Q_reg  ( .DIN(WX2051), .SDIN(n5912), .SSEL(test_se), .CLK(CK), .Q(n5905) );
  sdffs1 \DFF_280/Q_reg  ( .DIN(WX2049), .SDIN(n5919), .SSEL(test_se), .CLK(CK), .Q(n5912) );
  sdffs1 \DFF_279/Q_reg  ( .DIN(WX2047), .SDIN(n5926), .SSEL(test_se), .CLK(CK), .Q(n5919) );
  sdffs1 \DFF_278/Q_reg  ( .DIN(WX2045), .SDIN(n5933), .SSEL(test_se), .CLK(CK), .Q(n5926) );
  sdffs1 \DFF_277/Q_reg  ( .DIN(WX2043), .SDIN(n5940), .SSEL(test_se), .CLK(CK), .Q(n5933) );
  sdffs1 \DFF_276/Q_reg  ( .DIN(WX2041), .SDIN(n5947), .SSEL(test_se), .CLK(CK), .Q(n5940) );
  sdffs1 \DFF_275/Q_reg  ( .DIN(WX2039), .SDIN(n5954), .SSEL(test_se), .CLK(CK), .Q(n5947) );
  sdffs1 \DFF_274/Q_reg  ( .DIN(WX2037), .SDIN(n5961), .SSEL(test_se), .CLK(CK), .Q(n5954) );
  sdffs1 \DFF_273/Q_reg  ( .DIN(WX2035), .SDIN(n5968), .SSEL(test_se), .CLK(CK), .Q(n5961) );
  sdffs1 \DFF_272/Q_reg  ( .DIN(WX2033), .SDIN(n5976), .SSEL(test_se), .CLK(CK), .Q(n5968) );
  sdffs1 \DFF_271/Q_reg  ( .DIN(WX2031), .SDIN(n5985), .SSEL(test_se), .CLK(CK), .Q(n5976) );
  sdffs1 \DFF_270/Q_reg  ( .DIN(WX2029), .SDIN(n5994), .SSEL(test_se), .CLK(CK), .Q(n5985) );
  sdffs1 \DFF_269/Q_reg  ( .DIN(WX2027), .SDIN(n6003), .SSEL(test_se), .CLK(CK), .Q(n5994) );
  sdffs1 \DFF_268/Q_reg  ( .DIN(WX2025), .SDIN(n6012), .SSEL(test_se), .CLK(CK), .Q(n6003) );
  sdffs1 \DFF_267/Q_reg  ( .DIN(WX2023), .SDIN(n6021), .SSEL(test_se), .CLK(CK), .Q(n6012) );
  sdffs1 \DFF_266/Q_reg  ( .DIN(WX2021), .SDIN(n6030), .SSEL(test_se), .CLK(CK), .Q(n6021) );
  sdffs1 \DFF_265/Q_reg  ( .DIN(WX2019), .SDIN(n6039), .SSEL(test_se), .CLK(CK), .Q(n6030) );
  sdffs1 \DFF_264/Q_reg  ( .DIN(WX2017), .SDIN(n6048), .SSEL(test_se), .CLK(CK), .Q(n6039) );
  sdffs1 \DFF_263/Q_reg  ( .DIN(WX2015), .SDIN(n6057), .SSEL(test_se), .CLK(CK), .Q(n6048) );
  sdffs1 \DFF_262/Q_reg  ( .DIN(WX2013), .SDIN(n6066), .SSEL(test_se), .CLK(CK), .Q(n6057) );
  sdffs1 \DFF_261/Q_reg  ( .DIN(WX2011), .SDIN(n6075), .SSEL(test_se), .CLK(CK), .Q(n6066) );
  sdffs1 \DFF_260/Q_reg  ( .DIN(WX2009), .SDIN(n6084), .SSEL(test_se), .CLK(CK), .Q(n6075) );
  sdffs1 \DFF_259/Q_reg  ( .DIN(WX2007), .SDIN(n6093), .SSEL(test_se), .CLK(CK), .Q(n6084) );
  sdffs1 \DFF_258/Q_reg  ( .DIN(WX2005), .SDIN(n6102), .SSEL(test_se), .CLK(CK), .Q(n6093) );
  sdffs1 \DFF_257/Q_reg  ( .DIN(WX2003), .SDIN(n6111), .SSEL(test_se), .CLK(CK), .Q(n6102) );
  sdffs1 \DFF_256/Q_reg  ( .DIN(WX2001), .SDIN(n7034), .SSEL(test_se), .CLK(CK), .Q(n6111) );
  sdffs1 \DFF_255/Q_reg  ( .DIN(WX1999), .SDIN(n7033), .SSEL(test_se), .CLK(CK), .Q(n7034), .QN(n5862) );
  sdffs1 \DFF_254/Q_reg  ( .DIN(WX1997), .SDIN(n7032), .SSEL(test_se), .CLK(CK), .Q(n7033), .QN(n5869) );
  sdffs1 \DFF_253/Q_reg  ( .DIN(WX1995), .SDIN(n7031), .SSEL(test_se), .CLK(CK), .Q(n7032), .QN(n5876) );
  sdffs1 \DFF_252/Q_reg  ( .DIN(WX1993), .SDIN(n7030), .SSEL(test_se), .CLK(CK), .Q(n7031), .QN(n5883) );
  sdffs1 \DFF_251/Q_reg  ( .DIN(WX1991), .SDIN(n7029), .SSEL(test_se), .CLK(CK), .Q(n7030), .QN(n5890) );
  sdffs1 \DFF_250/Q_reg  ( .DIN(WX1989), .SDIN(n7028), .SSEL(test_se), .CLK(CK), .Q(n7029), .QN(n5897) );
  sdffs1 \DFF_249/Q_reg  ( .DIN(WX1987), .SDIN(n7027), .SSEL(test_se), .CLK(CK), .Q(n7028), .QN(n5904) );
  sdffs1 \DFF_248/Q_reg  ( .DIN(WX1985), .SDIN(n7026), .SSEL(test_se), .CLK(CK), .Q(n7027), .QN(n5911) );
  sdffs1 \DFF_247/Q_reg  ( .DIN(WX1983), .SDIN(n7025), .SSEL(test_se), .CLK(CK), .Q(n7026), .QN(n5918) );
  sdffs1 \DFF_246/Q_reg  ( .DIN(WX1981), .SDIN(n7024), .SSEL(test_se), .CLK(CK), .Q(n7025), .QN(n5925) );
  sdffs1 \DFF_245/Q_reg  ( .DIN(WX1979), .SDIN(n7023), .SSEL(test_se), .CLK(CK), .Q(n7024), .QN(n5932) );
  sdffs1 \DFF_244/Q_reg  ( .DIN(WX1977), .SDIN(n7022), .SSEL(test_se), .CLK(CK), .Q(n7023), .QN(n5939) );
  sdffs1 \DFF_243/Q_reg  ( .DIN(WX1975), .SDIN(n7021), .SSEL(test_se), .CLK(CK), .Q(n7022), .QN(n5946) );
  sdffs1 \DFF_242/Q_reg  ( .DIN(WX1973), .SDIN(n7020), .SSEL(test_se), .CLK(CK), .Q(n7021), .QN(n5953) );
  sdffs1 \DFF_241/Q_reg  ( .DIN(WX1971), .SDIN(n7019), .SSEL(test_se), .CLK(CK), .Q(n7020), .QN(n5960) );
  sdffs1 \DFF_240/Q_reg  ( .DIN(WX1969), .SDIN(n7018), .SSEL(test_se), .CLK(CK), .Q(n7019), .QN(n5967) );
  sdffs1 \DFF_239/Q_reg  ( .DIN(WX1967), .SDIN(n7017), .SSEL(test_se), .CLK(CK), .Q(n7018), .QN(n5975) );
  sdffs1 \DFF_238/Q_reg  ( .DIN(WX1965), .SDIN(n7016), .SSEL(test_se), .CLK(CK), .Q(n7017), .QN(n5984) );
  sdffs1 \DFF_237/Q_reg  ( .DIN(WX1963), .SDIN(n7015), .SSEL(test_se), .CLK(CK), .Q(n7016), .QN(n5993) );
  sdffs1 \DFF_236/Q_reg  ( .DIN(WX1961), .SDIN(n7014), .SSEL(test_se), .CLK(CK), .Q(n7015), .QN(n6002) );
  sdffs1 \DFF_235/Q_reg  ( .DIN(WX1959), .SDIN(n7013), .SSEL(test_se), .CLK(CK), .Q(n7014), .QN(n6011) );
  sdffs1 \DFF_234/Q_reg  ( .DIN(WX1957), .SDIN(n7012), .SSEL(test_se), .CLK(CK), .Q(n7013), .QN(n6020) );
  sdffs1 \DFF_233/Q_reg  ( .DIN(WX1955), .SDIN(n7011), .SSEL(test_se), .CLK(CK), .Q(n7012), .QN(n6029) );
  sdffs1 \DFF_232/Q_reg  ( .DIN(WX1953), .SDIN(n7010), .SSEL(test_se), .CLK(CK), .Q(n7011), .QN(n6038) );
  sdffs1 \DFF_231/Q_reg  ( .DIN(WX1951), .SDIN(n7009), .SSEL(test_se), .CLK(CK), .Q(n7010), .QN(n6047) );
  sdffs1 \DFF_230/Q_reg  ( .DIN(WX1949), .SDIN(n7008), .SSEL(test_se), .CLK(CK), .Q(n7009), .QN(n6056) );
  sdffs1 \DFF_229/Q_reg  ( .DIN(WX1947), .SDIN(n7007), .SSEL(test_se), .CLK(CK), .Q(n7008), .QN(n6065) );
  sdffs1 \DFF_228/Q_reg  ( .DIN(WX1945), .SDIN(n7006), .SSEL(test_se), .CLK(CK), .Q(n7007), .QN(n6074) );
  sdffs1 \DFF_227/Q_reg  ( .DIN(WX1943), .SDIN(n7005), .SSEL(test_se), .CLK(CK), .Q(n7006), .QN(n6083) );
  sdffs1 \DFF_226/Q_reg  ( .DIN(WX1941), .SDIN(n7004), .SSEL(test_se), .CLK(CK), .Q(n7005), .QN(n6092) );
  sdffs1 \DFF_225/Q_reg  ( .DIN(WX1939), .SDIN(n7003), .SSEL(test_se), .CLK(CK), .Q(n7004), .QN(n6101) );
  sdffs1 \DFF_224/Q_reg  ( .DIN(WX1937), .SDIN(n7002), .SSEL(test_se), .CLK(CK), .Q(n7003), .QN(n6110) );
  sdffs1 \DFF_223/Q_reg  ( .DIN(WX1839), .SDIN(n7001), .SSEL(test_se), .CLK(CK), .Q(n7002), .QN(n6116) );
  sdffs1 \DFF_222/Q_reg  ( .DIN(WX1837), .SDIN(n7000), .SSEL(test_se), .CLK(CK), .Q(n7001), .QN(n6117) );
  sdffs1 \DFF_221/Q_reg  ( .DIN(WX1835), .SDIN(n6999), .SSEL(test_se), .CLK(CK), .Q(n7000), .QN(n6118) );
  sdffs1 \DFF_220/Q_reg  ( .DIN(WX1833), .SDIN(n6998), .SSEL(test_se), .CLK(CK), .Q(n6999), .QN(n6119) );
  sdffs1 \DFF_219/Q_reg  ( .DIN(WX1831), .SDIN(n6997), .SSEL(test_se), .CLK(CK), .Q(n6998), .QN(n6120) );
  sdffs1 \DFF_218/Q_reg  ( .DIN(WX1829), .SDIN(n6996), .SSEL(test_se), .CLK(CK), .Q(n6997), .QN(n6121) );
  sdffs1 \DFF_217/Q_reg  ( .DIN(WX1827), .SDIN(n6995), .SSEL(test_se), .CLK(CK), .Q(n6996), .QN(n6122) );
  sdffs1 \DFF_216/Q_reg  ( .DIN(WX1825), .SDIN(n6994), .SSEL(test_se), .CLK(CK), .Q(n6995), .QN(n6123) );
  sdffs1 \DFF_215/Q_reg  ( .DIN(WX1823), .SDIN(n6993), .SSEL(test_se), .CLK(CK), .Q(n6994), .QN(n6124) );
  sdffs1 \DFF_214/Q_reg  ( .DIN(WX1821), .SDIN(n6992), .SSEL(test_se), .CLK(CK), .Q(n6993), .QN(n6125) );
  sdffs1 \DFF_213/Q_reg  ( .DIN(WX1819), .SDIN(n6991), .SSEL(test_se), .CLK(CK), .Q(n6992), .QN(n6126) );
  sdffs1 \DFF_212/Q_reg  ( .DIN(WX1817), .SDIN(n6990), .SSEL(test_se), .CLK(CK), .Q(n6991), .QN(n6127) );
  sdffs1 \DFF_211/Q_reg  ( .DIN(WX1815), .SDIN(n6989), .SSEL(test_se), .CLK(CK), .Q(n6990), .QN(n6128) );
  sdffs1 \DFF_210/Q_reg  ( .DIN(WX1813), .SDIN(n6988), .SSEL(test_se), .CLK(CK), .Q(n6989), .QN(n6129) );
  sdffs1 \DFF_209/Q_reg  ( .DIN(WX1811), .SDIN(n6987), .SSEL(test_se), .CLK(CK), .Q(n6988), .QN(n6130) );
  sdffs1 \DFF_208/Q_reg  ( .DIN(WX1809), .SDIN(n6986), .SSEL(test_se), .CLK(CK), .Q(n6987), .QN(n6131) );
  sdffs1 \DFF_207/Q_reg  ( .DIN(WX1807), .SDIN(n6985), .SSEL(test_se), .CLK(CK), .Q(n6986), .QN(n6132) );
  sdffs1 \DFF_206/Q_reg  ( .DIN(WX1805), .SDIN(n6984), .SSEL(test_se), .CLK(CK), .Q(n6985), .QN(n6133) );
  sdffs1 \DFF_205/Q_reg  ( .DIN(WX1803), .SDIN(n6983), .SSEL(test_se), .CLK(CK), .Q(n6984), .QN(n6134) );
  sdffs1 \DFF_204/Q_reg  ( .DIN(WX1801), .SDIN(n6982), .SSEL(test_se), .CLK(CK), .Q(n6983), .QN(n6135) );
  sdffs1 \DFF_203/Q_reg  ( .DIN(WX1799), .SDIN(n6981), .SSEL(test_se), .CLK(CK), .Q(n6982), .QN(n6136) );
  sdffs1 \DFF_202/Q_reg  ( .DIN(WX1797), .SDIN(n6980), .SSEL(test_se), .CLK(CK), .Q(n6981), .QN(n6137) );
  sdffs1 \DFF_201/Q_reg  ( .DIN(WX1795), .SDIN(n6979), .SSEL(test_se), .CLK(CK), .Q(n6980), .QN(n6138) );
  sdffs1 \DFF_200/Q_reg  ( .DIN(WX1793), .SDIN(n6978), .SSEL(test_se), .CLK(CK), .Q(n6979), .QN(n6139) );
  sdffs1 \DFF_199/Q_reg  ( .DIN(WX1791), .SDIN(n6977), .SSEL(test_se), .CLK(CK), .Q(n6978), .QN(n6140) );
  sdffs1 \DFF_198/Q_reg  ( .DIN(WX1789), .SDIN(n6976), .SSEL(test_se), .CLK(CK), .Q(n6977), .QN(n6141) );
  sdffs1 \DFF_197/Q_reg  ( .DIN(WX1787), .SDIN(n6975), .SSEL(test_se), .CLK(CK), .Q(n6976), .QN(n6142) );
  sdffs1 \DFF_196/Q_reg  ( .DIN(WX1785), .SDIN(n6974), .SSEL(test_se), .CLK(CK), .Q(n6975), .QN(n6143) );
  sdffs1 \DFF_195/Q_reg  ( .DIN(WX1783), .SDIN(n6973), .SSEL(test_se), .CLK(CK), .Q(n6974), .QN(n6144) );
  sdffs1 \DFF_194/Q_reg  ( .DIN(WX1781), .SDIN(n6972), .SSEL(test_se), .CLK(CK), .Q(n6973), .QN(n6145) );
  sdffs1 \DFF_193/Q_reg  ( .DIN(WX1779), .SDIN(n6971), .SSEL(test_se), .CLK(CK), .Q(n6972), .QN(n6146) );
  sdffs1 \DFF_192/Q_reg  ( .DIN(WX1777), .SDIN(CRC_OUT_9_31), .SSEL(test_se), 
        .CLK(CK), .Q(n6971), .QN(n6115) );
  sdffs1 \DFF_191/Q_reg  ( .DIN(WX1326), .SDIN(CRC_OUT_9_30), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_31), .QN(n6178) );
  sdffs1 \DFF_190/Q_reg  ( .DIN(WX1324), .SDIN(CRC_OUT_9_29), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_30), .QN(n6147) );
  sdffs1 \DFF_189/Q_reg  ( .DIN(WX1322), .SDIN(CRC_OUT_9_28), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_29), .QN(n6148) );
  sdffs1 \DFF_188/Q_reg  ( .DIN(WX1320), .SDIN(CRC_OUT_9_27), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_28), .QN(n6149) );
  sdffs1 \DFF_187/Q_reg  ( .DIN(WX1318), .SDIN(CRC_OUT_9_26), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_27), .QN(n6150) );
  sdffs1 \DFF_186/Q_reg  ( .DIN(WX1316), .SDIN(CRC_OUT_9_25), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_26), .QN(n6151) );
  sdffs1 \DFF_185/Q_reg  ( .DIN(WX1314), .SDIN(CRC_OUT_9_24), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_25), .QN(n6152) );
  sdffs1 \DFF_184/Q_reg  ( .DIN(WX1312), .SDIN(CRC_OUT_9_23), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_24), .QN(n6153) );
  sdffs1 \DFF_183/Q_reg  ( .DIN(WX1310), .SDIN(CRC_OUT_9_22), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_23), .QN(n6154) );
  sdffs1 \DFF_182/Q_reg  ( .DIN(WX1308), .SDIN(CRC_OUT_9_21), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_22), .QN(n6155) );
  sdffs1 \DFF_181/Q_reg  ( .DIN(WX1306), .SDIN(CRC_OUT_9_20), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_21), .QN(n6156) );
  sdffs1 \DFF_180/Q_reg  ( .DIN(WX1304), .SDIN(CRC_OUT_9_19), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_20), .QN(n6157) );
  sdffs1 \DFF_179/Q_reg  ( .DIN(WX1302), .SDIN(CRC_OUT_9_18), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_19), .QN(n6158) );
  sdffs1 \DFF_178/Q_reg  ( .DIN(WX1300), .SDIN(CRC_OUT_9_17), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_18), .QN(n6159) );
  sdffs1 \DFF_177/Q_reg  ( .DIN(WX1298), .SDIN(CRC_OUT_9_16), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_17), .QN(n6160) );
  sdffs1 \DFF_176/Q_reg  ( .DIN(WX1296), .SDIN(CRC_OUT_9_15), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_16), .QN(n6161) );
  sdffs1 \DFF_175/Q_reg  ( .DIN(WX1294), .SDIN(CRC_OUT_9_14), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_15), .QN(n6162) );
  sdffs1 \DFF_174/Q_reg  ( .DIN(WX1292), .SDIN(CRC_OUT_9_13), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_14), .QN(n6163) );
  sdffs1 \DFF_173/Q_reg  ( .DIN(WX1290), .SDIN(CRC_OUT_9_12), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_13), .QN(n6164) );
  sdffs1 \DFF_172/Q_reg  ( .DIN(WX1288), .SDIN(CRC_OUT_9_11), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_12), .QN(n6165) );
  sdffs1 \DFF_171/Q_reg  ( .DIN(WX1286), .SDIN(CRC_OUT_9_10), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_11), .QN(n6166) );
  sdffs1 \DFF_170/Q_reg  ( .DIN(WX1284), .SDIN(CRC_OUT_9_9), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_10), .QN(n6167) );
  sdffs1 \DFF_169/Q_reg  ( .DIN(WX1282), .SDIN(CRC_OUT_9_8), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_9), .QN(n6168) );
  sdffs1 \DFF_168/Q_reg  ( .DIN(WX1280), .SDIN(CRC_OUT_9_7), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_8), .QN(n6169) );
  sdffs1 \DFF_167/Q_reg  ( .DIN(WX1278), .SDIN(CRC_OUT_9_6), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_7), .QN(n6170) );
  sdffs1 \DFF_166/Q_reg  ( .DIN(WX1276), .SDIN(CRC_OUT_9_5), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_6), .QN(n6171) );
  sdffs1 \DFF_165/Q_reg  ( .DIN(WX1274), .SDIN(CRC_OUT_9_4), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_5), .QN(n6172) );
  sdffs1 \DFF_164/Q_reg  ( .DIN(WX1272), .SDIN(CRC_OUT_9_3), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_4), .QN(n6173) );
  sdffs1 \DFF_163/Q_reg  ( .DIN(WX1270), .SDIN(CRC_OUT_9_2), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_3), .QN(n6174) );
  sdffs1 \DFF_162/Q_reg  ( .DIN(WX1268), .SDIN(CRC_OUT_9_1), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_2), .QN(n6175) );
  sdffs1 \DFF_161/Q_reg  ( .DIN(WX1266), .SDIN(CRC_OUT_9_0), .SSEL(test_se), 
        .CLK(CK), .Q(CRC_OUT_9_1), .QN(n6176) );
  sdffs1 \DFF_160/Q_reg  ( .DIN(WX1264), .SDIN(n6970), .SSEL(test_se), .CLK(CK), .Q(CRC_OUT_9_0), .QN(n6177) );
  sdffs1 \DFF_159/Q_reg  ( .DIN(WX898), .SDIN(n6969), .SSEL(test_se), .CLK(CK), 
        .Q(n6970), .QN(n6462) );
  sdffs1 \DFF_158/Q_reg  ( .DIN(WX896), .SDIN(n6968), .SSEL(test_se), .CLK(CK), 
        .Q(n6969), .QN(n6530) );
  sdffs1 \DFF_157/Q_reg  ( .DIN(WX894), .SDIN(n6967), .SSEL(test_se), .CLK(CK), 
        .Q(n6968), .QN(n6437) );
  sdffs1 \DFF_156/Q_reg  ( .DIN(WX892), .SDIN(n6966), .SSEL(test_se), .CLK(CK), 
        .Q(n6967), .QN(n6468) );
  sdffs1 \DFF_155/Q_reg  ( .DIN(WX890), .SDIN(n6965), .SSEL(test_se), .CLK(CK), 
        .Q(n6966), .QN(n6471) );
  sdffs1 \DFF_154/Q_reg  ( .DIN(WX888), .SDIN(n6964), .SSEL(test_se), .CLK(CK), 
        .Q(n6965), .QN(n6459) );
  sdffs1 \DFF_153/Q_reg  ( .DIN(WX886), .SDIN(n6963), .SSEL(test_se), .CLK(CK), 
        .Q(n6964), .QN(n6441) );
  sdffs1 \DFF_152/Q_reg  ( .DIN(WX884), .SDIN(n6962), .SSEL(test_se), .CLK(CK), 
        .Q(n6963), .QN(n6465) );
  sdffs1 \DFF_151/Q_reg  ( .DIN(WX882), .SDIN(n6961), .SSEL(test_se), .CLK(CK), 
        .Q(n6962), .QN(n6453) );
  sdffs1 \DFF_150/Q_reg  ( .DIN(WX880), .SDIN(n6960), .SSEL(test_se), .CLK(CK), 
        .Q(n6961), .QN(n6506) );
  sdffs1 \DFF_149/Q_reg  ( .DIN(WX878), .SDIN(n6959), .SSEL(test_se), .CLK(CK), 
        .Q(n6960), .QN(n6450) );
  sdffs1 \DFF_148/Q_reg  ( .DIN(WX876), .SDIN(n6958), .SSEL(test_se), .CLK(CK), 
        .Q(n6959), .QN(n6444) );
  sdffs1 \DFF_147/Q_reg  ( .DIN(WX874), .SDIN(n6957), .SSEL(test_se), .CLK(CK), 
        .Q(n6958), .QN(n6456) );
  sdffs1 \DFF_146/Q_reg  ( .DIN(WX872), .SDIN(n6956), .SSEL(test_se), .CLK(CK), 
        .Q(n6957), .QN(n6447) );
  sdffs1 \DFF_145/Q_reg  ( .DIN(WX870), .SDIN(n6955), .SSEL(test_se), .CLK(CK), 
        .Q(n6956), .QN(n6525) );
  sdffs1 \DFF_144/Q_reg  ( .DIN(WX868), .SDIN(n6954), .SSEL(test_se), .CLK(CK), 
        .Q(n6955), .QN(n6438) );
  sdffs1 \DFF_143/Q_reg  ( .DIN(WX866), .SDIN(n6953), .SSEL(test_se), .CLK(CK), 
        .Q(n6954), .QN(n6510) );
  sdffs1 \DFF_142/Q_reg  ( .DIN(WX864), .SDIN(n6952), .SSEL(test_se), .CLK(CK), 
        .Q(n6953), .QN(n6495) );
  sdffs1 \DFF_141/Q_reg  ( .DIN(WX862), .SDIN(n6951), .SSEL(test_se), .CLK(CK), 
        .Q(n6952), .QN(n6491) );
  sdffs1 \DFF_140/Q_reg  ( .DIN(WX860), .SDIN(n6950), .SSEL(test_se), .CLK(CK), 
        .Q(n6951), .QN(n6477) );
  sdffs1 \DFF_139/Q_reg  ( .DIN(WX858), .SDIN(n6949), .SSEL(test_se), .CLK(CK), 
        .Q(n6950), .QN(n6522) );
  sdffs1 \DFF_138/Q_reg  ( .DIN(WX856), .SDIN(n6948), .SSEL(test_se), .CLK(CK), 
        .Q(n6949), .QN(n6517) );
  sdffs1 \DFF_137/Q_reg  ( .DIN(WX854), .SDIN(n6947), .SSEL(test_se), .CLK(CK), 
        .Q(n6948), .QN(n6516) );
  sdffs1 \DFF_136/Q_reg  ( .DIN(WX852), .SDIN(n6946), .SSEL(test_se), .CLK(CK), 
        .Q(n6947), .QN(n6511) );
  sdffs1 \DFF_135/Q_reg  ( .DIN(WX850), .SDIN(n6945), .SSEL(test_se), .CLK(CK), 
        .Q(n6946), .QN(n6501) );
  sdffs1 \DFF_134/Q_reg  ( .DIN(WX848), .SDIN(n6944), .SSEL(test_se), .CLK(CK), 
        .Q(n6945), .QN(n6500) );
  sdffs1 \DFF_133/Q_reg  ( .DIN(WX846), .SDIN(n6943), .SSEL(test_se), .CLK(CK), 
        .Q(n6944), .QN(n6492) );
  sdffs1 \DFF_132/Q_reg  ( .DIN(WX844), .SDIN(n6942), .SSEL(test_se), .CLK(CK), 
        .Q(n6943), .QN(n6486) );
  sdffs1 \DFF_131/Q_reg  ( .DIN(WX842), .SDIN(n6941), .SSEL(test_se), .CLK(CK), 
        .Q(n6942), .QN(n6483) );
  sdffs1 \DFF_130/Q_reg  ( .DIN(WX840), .SDIN(n6940), .SSEL(test_se), .CLK(CK), 
        .Q(n6941), .QN(n6482) );
  sdffs1 \DFF_129/Q_reg  ( .DIN(WX838), .SDIN(n6939), .SSEL(test_se), .CLK(CK), 
        .Q(n6940), .QN(n6474) );
  sdffs1 \DFF_128/Q_reg  ( .DIN(WX836), .SDIN(n6938), .SSEL(test_se), .CLK(CK), 
        .Q(n6939), .QN(n6534) );
  sdffs1 \DFF_127/Q_reg  ( .DIN(WX834), .SDIN(n6937), .SSEL(test_se), .CLK(CK), 
        .Q(n6938), .QN(n6463) );
  sdffs1 \DFF_126/Q_reg  ( .DIN(WX832), .SDIN(n6936), .SSEL(test_se), .CLK(CK), 
        .Q(n6937), .QN(n6527) );
  sdffs1 \DFF_125/Q_reg  ( .DIN(WX830), .SDIN(n6935), .SSEL(test_se), .CLK(CK), 
        .Q(n6936), .QN(n6436) );
  sdffs1 \DFF_124/Q_reg  ( .DIN(WX828), .SDIN(n6934), .SSEL(test_se), .CLK(CK), 
        .Q(n6935), .QN(n6469) );
  sdffs1 \DFF_123/Q_reg  ( .DIN(WX826), .SDIN(n6933), .SSEL(test_se), .CLK(CK), 
        .Q(n6934), .QN(n6472) );
  sdffs1 \DFF_122/Q_reg  ( .DIN(WX824), .SDIN(n6932), .SSEL(test_se), .CLK(CK), 
        .Q(n6933), .QN(n6460) );
  sdffs1 \DFF_121/Q_reg  ( .DIN(WX822), .SDIN(n6931), .SSEL(test_se), .CLK(CK), 
        .Q(n6932), .QN(n6442) );
  sdffs1 \DFF_120/Q_reg  ( .DIN(WX820), .SDIN(n6930), .SSEL(test_se), .CLK(CK), 
        .Q(n6931), .QN(n6466) );
  sdffs1 \DFF_119/Q_reg  ( .DIN(WX818), .SDIN(n6929), .SSEL(test_se), .CLK(CK), 
        .Q(n6930), .QN(n6454) );
  sdffs1 \DFF_118/Q_reg  ( .DIN(WX816), .SDIN(n6928), .SSEL(test_se), .CLK(CK), 
        .Q(n6929), .QN(n6504) );
  sdffs1 \DFF_117/Q_reg  ( .DIN(WX814), .SDIN(n6927), .SSEL(test_se), .CLK(CK), 
        .Q(n6928), .QN(n6451) );
  sdffs1 \DFF_116/Q_reg  ( .DIN(WX812), .SDIN(n6926), .SSEL(test_se), .CLK(CK), 
        .Q(n6927), .QN(n6445) );
  sdffs1 \DFF_115/Q_reg  ( .DIN(WX810), .SDIN(n6925), .SSEL(test_se), .CLK(CK), 
        .Q(n6926), .QN(n6457) );
  sdffs1 \DFF_114/Q_reg  ( .DIN(WX808), .SDIN(n6924), .SSEL(test_se), .CLK(CK), 
        .Q(n6925), .QN(n6448) );
  sdffs1 \DFF_113/Q_reg  ( .DIN(WX806), .SDIN(n6923), .SSEL(test_se), .CLK(CK), 
        .Q(n6924), .QN(n6523) );
  sdffs1 \DFF_112/Q_reg  ( .DIN(WX804), .SDIN(n6922), .SSEL(test_se), .CLK(CK), 
        .Q(n6923), .QN(n6439) );
  sdffs1 \DFF_111/Q_reg  ( .DIN(WX802), .SDIN(n6921), .SSEL(test_se), .CLK(CK), 
        .Q(n6922), .QN(n6539) );
  sdffs1 \DFF_110/Q_reg  ( .DIN(WX800), .SDIN(n6920), .SSEL(test_se), .CLK(CK), 
        .Q(n6921), .QN(n6496) );
  sdffs1 \DFF_109/Q_reg  ( .DIN(WX798), .SDIN(n6919), .SSEL(test_se), .CLK(CK), 
        .Q(n6920), .QN(n6544) );
  sdffs1 \DFF_108/Q_reg  ( .DIN(WX796), .SDIN(n6918), .SSEL(test_se), .CLK(CK), 
        .Q(n6919), .QN(n6478) );
  sdffs1 \DFF_107/Q_reg  ( .DIN(WX794), .SDIN(n6917), .SSEL(test_se), .CLK(CK), 
        .Q(n6918), .QN(n6535) );
  sdffs1 \DFF_106/Q_reg  ( .DIN(WX792), .SDIN(n6916), .SSEL(test_se), .CLK(CK), 
        .Q(n6917), .QN(n6518) );
  sdffs1 \DFF_105/Q_reg  ( .DIN(WX790), .SDIN(n6915), .SSEL(test_se), .CLK(CK), 
        .Q(n6916), .QN(n6537) );
  sdffs1 \DFF_104/Q_reg  ( .DIN(WX788), .SDIN(n6914), .SSEL(test_se), .CLK(CK), 
        .Q(n6915), .QN(n6512) );
  sdffs1 \DFF_103/Q_reg  ( .DIN(WX786), .SDIN(n6913), .SSEL(test_se), .CLK(CK), 
        .Q(n6914), .QN(n6502) );
  sdffs1 \DFF_102/Q_reg  ( .DIN(WX784), .SDIN(n6912), .SSEL(test_se), .CLK(CK), 
        .Q(n6913), .QN(n6541) );
  sdffs1 \DFF_101/Q_reg  ( .DIN(WX782), .SDIN(n6911), .SSEL(test_se), .CLK(CK), 
        .Q(n6912), .QN(n6493) );
  sdffs1 \DFF_100/Q_reg  ( .DIN(WX780), .SDIN(n6910), .SSEL(test_se), .CLK(CK), 
        .Q(n6911), .QN(n6487) );
  sdffs1 \DFF_99/Q_reg  ( .DIN(WX778), .SDIN(n6909), .SSEL(test_se), .CLK(CK), 
        .Q(n6910), .QN(n6484) );
  sdffs1 \DFF_98/Q_reg  ( .DIN(WX776), .SDIN(n6908), .SSEL(test_se), .CLK(CK), 
        .Q(n6909), .QN(n6547) );
  sdffs1 \DFF_97/Q_reg  ( .DIN(WX774), .SDIN(n6907), .SSEL(test_se), .CLK(CK), 
        .Q(n6908), .QN(n6475) );
  sdffs1 \DFF_96/Q_reg  ( .DIN(WX772), .SDIN(n6906), .SSEL(test_se), .CLK(CK), 
        .Q(n6907), .QN(n6531) );
  sdffs1 \DFF_95/Q_reg  ( .DIN(WX770), .SDIN(n6905), .SSEL(test_se), .CLK(CK), 
        .Q(n6906), .QN(n6464) );
  sdffs1 \DFF_94/Q_reg  ( .DIN(WX768), .SDIN(n6904), .SSEL(test_se), .CLK(CK), 
        .Q(n6905), .QN(n6528) );
  sdffs1 \DFF_93/Q_reg  ( .DIN(WX766), .SDIN(n6903), .SSEL(test_se), .CLK(CK), 
        .Q(n6904), .QN(n6562) );
  sdffs1 \DFF_92/Q_reg  ( .DIN(WX764), .SDIN(n6902), .SSEL(test_se), .CLK(CK), 
        .Q(n6903), .QN(n6470) );
  sdffs1 \DFF_91/Q_reg  ( .DIN(WX762), .SDIN(n6901), .SSEL(test_se), .CLK(CK), 
        .Q(n6902), .QN(n6473) );
  sdffs1 \DFF_90/Q_reg  ( .DIN(WX760), .SDIN(n6900), .SSEL(test_se), .CLK(CK), 
        .Q(n6901), .QN(n6461) );
  sdffs1 \DFF_89/Q_reg  ( .DIN(WX758), .SDIN(n6899), .SSEL(test_se), .CLK(CK), 
        .Q(n6900), .QN(n6443) );
  sdffs1 \DFF_88/Q_reg  ( .DIN(WX756), .SDIN(n6898), .SSEL(test_se), .CLK(CK), 
        .Q(n6899), .QN(n6467) );
  sdffs1 \DFF_87/Q_reg  ( .DIN(WX754), .SDIN(n6897), .SSEL(test_se), .CLK(CK), 
        .Q(n6898), .QN(n6455) );
  sdffs1 \DFF_86/Q_reg  ( .DIN(WX752), .SDIN(n6896), .SSEL(test_se), .CLK(CK), 
        .Q(n6897), .QN(n6505) );
  sdffs1 \DFF_85/Q_reg  ( .DIN(WX750), .SDIN(n6895), .SSEL(test_se), .CLK(CK), 
        .Q(n6896), .QN(n6452) );
  sdffs1 \DFF_84/Q_reg  ( .DIN(WX748), .SDIN(n6894), .SSEL(test_se), .CLK(CK), 
        .Q(n6895), .QN(n6446) );
  sdffs1 \DFF_83/Q_reg  ( .DIN(WX746), .SDIN(n6893), .SSEL(test_se), .CLK(CK), 
        .Q(n6894), .QN(n6458) );
  sdffs1 \DFF_82/Q_reg  ( .DIN(WX744), .SDIN(n6892), .SSEL(test_se), .CLK(CK), 
        .Q(n6893), .QN(n6449) );
  sdffs1 \DFF_81/Q_reg  ( .DIN(WX742), .SDIN(n6891), .SSEL(test_se), .CLK(CK), 
        .Q(n6892), .QN(n6524) );
  sdffs1 \DFF_80/Q_reg  ( .DIN(WX740), .SDIN(n6890), .SSEL(test_se), .CLK(CK), 
        .Q(n6891), .QN(n6440) );
  sdffs1 \DFF_79/Q_reg  ( .DIN(WX738), .SDIN(n6889), .SSEL(test_se), .CLK(CK), 
        .Q(n6890), .QN(n6508) );
  sdffs1 \DFF_78/Q_reg  ( .DIN(WX736), .SDIN(n6888), .SSEL(test_se), .CLK(CK), 
        .Q(n6889), .QN(n6497) );
  sdffs1 \DFF_77/Q_reg  ( .DIN(WX734), .SDIN(n6887), .SSEL(test_se), .CLK(CK), 
        .Q(n6888), .QN(n6489) );
  sdffs1 \DFF_76/Q_reg  ( .DIN(WX732), .SDIN(n6886), .SSEL(test_se), .CLK(CK), 
        .Q(n6887), .QN(n6479) );
  sdffs1 \DFF_75/Q_reg  ( .DIN(WX730), .SDIN(n6885), .SSEL(test_se), .CLK(CK), 
        .Q(n6886), .QN(n6520) );
  sdffs1 \DFF_74/Q_reg  ( .DIN(WX728), .SDIN(n6884), .SSEL(test_se), .CLK(CK), 
        .Q(n6885), .QN(n6519) );
  sdffs1 \DFF_73/Q_reg  ( .DIN(WX726), .SDIN(n6883), .SSEL(test_se), .CLK(CK), 
        .Q(n6884), .QN(n6514) );
  sdffs1 \DFF_72/Q_reg  ( .DIN(WX724), .SDIN(n6882), .SSEL(test_se), .CLK(CK), 
        .Q(n6883), .QN(n6513) );
  sdffs1 \DFF_71/Q_reg  ( .DIN(WX722), .SDIN(n6881), .SSEL(test_se), .CLK(CK), 
        .Q(n6882), .QN(n6503) );
  sdffs1 \DFF_70/Q_reg  ( .DIN(WX720), .SDIN(n6880), .SSEL(test_se), .CLK(CK), 
        .Q(n6881), .QN(n6498) );
  sdffs1 \DFF_69/Q_reg  ( .DIN(WX718), .SDIN(n6879), .SSEL(test_se), .CLK(CK), 
        .Q(n6880), .QN(n6494) );
  sdffs1 \DFF_68/Q_reg  ( .DIN(WX716), .SDIN(n6878), .SSEL(test_se), .CLK(CK), 
        .Q(n6879), .QN(n6488) );
  sdffs1 \DFF_67/Q_reg  ( .DIN(WX714), .SDIN(n6877), .SSEL(test_se), .CLK(CK), 
        .Q(n6878), .QN(n6485) );
  sdffs1 \DFF_66/Q_reg  ( .DIN(WX712), .SDIN(n6876), .SSEL(test_se), .CLK(CK), 
        .Q(n6877), .QN(n6480) );
  sdffs1 \DFF_65/Q_reg  ( .DIN(WX710), .SDIN(n6875), .SSEL(test_se), .CLK(CK), 
        .Q(n6876), .QN(n6476) );
  sdffs1 \DFF_64/Q_reg  ( .DIN(WX708), .SDIN(n6874), .SSEL(test_se), .CLK(CK), 
        .Q(n6875), .QN(n6532) );
  sdffs1 \DFF_63/Q_reg  ( .DIN(WX706), .SDIN(n6873), .SSEL(test_se), .CLK(CK), 
        .Q(n6874), .QN(n6553) );
  sdffs1 \DFF_62/Q_reg  ( .DIN(WX704), .SDIN(n6872), .SSEL(test_se), .CLK(CK), 
        .Q(n6873), .QN(n6529) );
  sdffs1 \DFF_61/Q_reg  ( .DIN(WX702), .SDIN(n6871), .SSEL(test_se), .CLK(CK), 
        .Q(n6872), .QN(n6435) );
  sdffs1 \DFF_60/Q_reg  ( .DIN(WX700), .SDIN(n6870), .SSEL(test_se), .CLK(CK), 
        .Q(n6871), .QN(n6551) );
  sdffs1 \DFF_59/Q_reg  ( .DIN(WX698), .SDIN(n6869), .SSEL(test_se), .CLK(CK), 
        .Q(n6870), .QN(n6550) );
  sdffs1 \DFF_58/Q_reg  ( .DIN(WX696), .SDIN(n6868), .SSEL(test_se), .CLK(CK), 
        .Q(n6869), .QN(n6554) );
  sdffs1 \DFF_57/Q_reg  ( .DIN(WX694), .SDIN(n6867), .SSEL(test_se), .CLK(CK), 
        .Q(n6868), .QN(n6560) );
  sdffs1 \DFF_56/Q_reg  ( .DIN(WX692), .SDIN(n6866), .SSEL(test_se), .CLK(CK), 
        .Q(n6867), .QN(n6552) );
  sdffs1 \DFF_55/Q_reg  ( .DIN(WX690), .SDIN(n6865), .SSEL(test_se), .CLK(CK), 
        .Q(n6866), .QN(n6556) );
  sdffs1 \DFF_54/Q_reg  ( .DIN(WX688), .SDIN(n6864), .SSEL(test_se), .CLK(CK), 
        .Q(n6865), .QN(n6507) );
  sdffs1 \DFF_53/Q_reg  ( .DIN(WX686), .SDIN(n6863), .SSEL(test_se), .CLK(CK), 
        .Q(n6864), .QN(n6557) );
  sdffs1 \DFF_52/Q_reg  ( .DIN(WX684), .SDIN(n6862), .SSEL(test_se), .CLK(CK), 
        .Q(n6863), .QN(n6559) );
  sdffs1 \DFF_51/Q_reg  ( .DIN(WX682), .SDIN(n6861), .SSEL(test_se), .CLK(CK), 
        .Q(n6862), .QN(n6555) );
  sdffs1 \DFF_50/Q_reg  ( .DIN(WX680), .SDIN(n6860), .SSEL(test_se), .CLK(CK), 
        .Q(n6861), .QN(n6558) );
  sdffs1 \DFF_49/Q_reg  ( .DIN(WX678), .SDIN(n6859), .SSEL(test_se), .CLK(CK), 
        .Q(n6860), .QN(n6526) );
  sdffs1 \DFF_48/Q_reg  ( .DIN(WX676), .SDIN(n6858), .SSEL(test_se), .CLK(CK), 
        .Q(n6859), .QN(n6561) );
  sdffs1 \DFF_47/Q_reg  ( .DIN(WX674), .SDIN(n6857), .SSEL(test_se), .CLK(CK), 
        .Q(n6858), .QN(n6509) );
  sdffs1 \DFF_46/Q_reg  ( .DIN(WX672), .SDIN(n6856), .SSEL(test_se), .CLK(CK), 
        .Q(n6857), .QN(n6542) );
  sdffs1 \DFF_45/Q_reg  ( .DIN(WX670), .SDIN(n6855), .SSEL(test_se), .CLK(CK), 
        .Q(n6856), .QN(n6490) );
  sdffs1 \DFF_44/Q_reg  ( .DIN(WX668), .SDIN(n6854), .SSEL(test_se), .CLK(CK), 
        .Q(n6855), .QN(n6548) );
  sdffs1 \DFF_43/Q_reg  ( .DIN(WX666), .SDIN(n6853), .SSEL(test_se), .CLK(CK), 
        .Q(n6854), .QN(n6521) );
  sdffs1 \DFF_42/Q_reg  ( .DIN(WX664), .SDIN(n6852), .SSEL(test_se), .CLK(CK), 
        .Q(n6853), .QN(n6536) );
  sdffs1 \DFF_41/Q_reg  ( .DIN(WX662), .SDIN(n6851), .SSEL(test_se), .CLK(CK), 
        .Q(n6852), .QN(n6515) );
  sdffs1 \DFF_40/Q_reg  ( .DIN(WX660), .SDIN(n6850), .SSEL(test_se), .CLK(CK), 
        .Q(n6851), .QN(n6538) );
  sdffs1 \DFF_39/Q_reg  ( .DIN(WX658), .SDIN(n6849), .SSEL(test_se), .CLK(CK), 
        .Q(n6850), .QN(n6540) );
  sdffs1 \DFF_38/Q_reg  ( .DIN(WX656), .SDIN(n6848), .SSEL(test_se), .CLK(CK), 
        .Q(n6849), .QN(n6499) );
  sdffs1 \DFF_37/Q_reg  ( .DIN(WX654), .SDIN(n6847), .SSEL(test_se), .CLK(CK), 
        .Q(n6848), .QN(n6543) );
  sdffs1 \DFF_36/Q_reg  ( .DIN(WX652), .SDIN(n6846), .SSEL(test_se), .CLK(CK), 
        .Q(n6847), .QN(n6545) );
  sdffs1 \DFF_35/Q_reg  ( .DIN(WX650), .SDIN(n6845), .SSEL(test_se), .CLK(CK), 
        .Q(n6846), .QN(n6546) );
  sdffs1 \DFF_34/Q_reg  ( .DIN(WX648), .SDIN(n6844), .SSEL(test_se), .CLK(CK), 
        .Q(n6845), .QN(n6481) );
  sdffs1 \DFF_33/Q_reg  ( .DIN(WX646), .SDIN(n6843), .SSEL(test_se), .CLK(CK), 
        .Q(n6844), .QN(n6549) );
  sdffs1 \DFF_32/Q_reg  ( .DIN(WX644), .SDIN(n6842), .SSEL(test_se), .CLK(CK), 
        .Q(n6843), .QN(n6533) );
  sdffs1 \DFF_31/Q_reg  ( .DIN(WX546), .SDIN(n6841), .SSEL(test_se), .CLK(CK), 
        .Q(n6842), .QN(n6179) );
  sdffs1 \DFF_30/Q_reg  ( .DIN(WX544), .SDIN(n6840), .SSEL(test_se), .CLK(CK), 
        .Q(n6841), .QN(n6180) );
  sdffs1 \DFF_29/Q_reg  ( .DIN(WX542), .SDIN(n6839), .SSEL(test_se), .CLK(CK), 
        .Q(n6840), .QN(n6181) );
  sdffs1 \DFF_28/Q_reg  ( .DIN(WX540), .SDIN(n6838), .SSEL(test_se), .CLK(CK), 
        .Q(n6839), .QN(n6182) );
  sdffs1 \DFF_27/Q_reg  ( .DIN(WX538), .SDIN(n6837), .SSEL(test_se), .CLK(CK), 
        .Q(n6838), .QN(n6183) );
  sdffs1 \DFF_26/Q_reg  ( .DIN(WX536), .SDIN(n6836), .SSEL(test_se), .CLK(CK), 
        .Q(n6837), .QN(n6184) );
  sdffs1 \DFF_25/Q_reg  ( .DIN(WX534), .SDIN(n6835), .SSEL(test_se), .CLK(CK), 
        .Q(n6836), .QN(n6185) );
  sdffs1 \DFF_24/Q_reg  ( .DIN(WX532), .SDIN(n6834), .SSEL(test_se), .CLK(CK), 
        .Q(n6835), .QN(n6186) );
  sdffs1 \DFF_23/Q_reg  ( .DIN(WX530), .SDIN(n6833), .SSEL(test_se), .CLK(CK), 
        .Q(n6834), .QN(n6187) );
  sdffs1 \DFF_22/Q_reg  ( .DIN(WX528), .SDIN(n6832), .SSEL(test_se), .CLK(CK), 
        .Q(n6833), .QN(n6188) );
  sdffs1 \DFF_21/Q_reg  ( .DIN(WX526), .SDIN(n6831), .SSEL(test_se), .CLK(CK), 
        .Q(n6832), .QN(n6189) );
  sdffs1 \DFF_20/Q_reg  ( .DIN(WX524), .SDIN(n6830), .SSEL(test_se), .CLK(CK), 
        .Q(n6831), .QN(n6190) );
  sdffs1 \DFF_19/Q_reg  ( .DIN(WX522), .SDIN(n6829), .SSEL(test_se), .CLK(CK), 
        .Q(n6830), .QN(n6191) );
  sdffs1 \DFF_18/Q_reg  ( .DIN(WX520), .SDIN(n6828), .SSEL(test_se), .CLK(CK), 
        .Q(n6829), .QN(n6192) );
  sdffs1 \DFF_17/Q_reg  ( .DIN(WX518), .SDIN(n6827), .SSEL(test_se), .CLK(CK), 
        .Q(n6828), .QN(n6193) );
  sdffs1 \DFF_16/Q_reg  ( .DIN(WX516), .SDIN(n6826), .SSEL(test_se), .CLK(CK), 
        .Q(n6827), .QN(n6194) );
  sdffs1 \DFF_15/Q_reg  ( .DIN(WX514), .SDIN(n6825), .SSEL(test_se), .CLK(CK), 
        .Q(n6826), .QN(n6195) );
  sdffs1 \DFF_14/Q_reg  ( .DIN(WX512), .SDIN(n6824), .SSEL(test_se), .CLK(CK), 
        .Q(n6825), .QN(n6196) );
  sdffs1 \DFF_13/Q_reg  ( .DIN(WX510), .SDIN(n6823), .SSEL(test_se), .CLK(CK), 
        .Q(n6824), .QN(n6286) );
  sdffs1 \DFF_12/Q_reg  ( .DIN(WX508), .SDIN(n6822), .SSEL(test_se), .CLK(CK), 
        .Q(n6823), .QN(n6342) );
  sdffs1 \DFF_11/Q_reg  ( .DIN(WX506), .SDIN(n6821), .SSEL(test_se), .CLK(CK), 
        .Q(n6822), .QN(n6354) );
  sdffs1 \DFF_10/Q_reg  ( .DIN(WX504), .SDIN(n6820), .SSEL(test_se), .CLK(CK), 
        .Q(n6821), .QN(n6376) );
  sdffs1 \DFF_9/Q_reg  ( .DIN(WX502), .SDIN(n6819), .SSEL(test_se), .CLK(CK), 
        .Q(n6820), .QN(n6377) );
  sdffs1 \DFF_8/Q_reg  ( .DIN(WX500), .SDIN(n6818), .SSEL(test_se), .CLK(CK), 
        .Q(n6819), .QN(n6378) );
  sdffs1 \DFF_7/Q_reg  ( .DIN(WX498), .SDIN(n6817), .SSEL(test_se), .CLK(CK), 
        .Q(n6818), .QN(n6379) );
  sdffs1 \DFF_6/Q_reg  ( .DIN(WX496), .SDIN(n6816), .SSEL(test_se), .CLK(CK), 
        .Q(n6817), .QN(n6380) );
  sdffs1 \DFF_5/Q_reg  ( .DIN(WX494), .SDIN(n6815), .SSEL(test_se), .CLK(CK), 
        .Q(n6816), .QN(n6381) );
  sdffs1 \DFF_4/Q_reg  ( .DIN(WX492), .SDIN(n6814), .SSEL(test_se), .CLK(CK), 
        .Q(n6815), .QN(n6382) );
  sdffs1 \DFF_3/Q_reg  ( .DIN(WX490), .SDIN(n6813), .SSEL(test_se), .CLK(CK), 
        .Q(n6814), .QN(n6431) );
  sdffs1 \DFF_2/Q_reg  ( .DIN(WX488), .SDIN(n6812), .SSEL(test_se), .CLK(CK), 
        .Q(n6813), .QN(n6432) );
  sdffs1 \DFF_1/Q_reg  ( .DIN(WX486), .SDIN(n6811), .SSEL(test_se), .CLK(CK), 
        .Q(n6812), .QN(n6433) );
  sdffs1 \DFF_0/Q_reg  ( .DIN(WX484), .SDIN(test_si), .SSEL(test_se), .CLK(CK), 
        .Q(n6811), .QN(n6434) );
  nor5s1 trig32_0U1 ( .DIN1(trig32_0n1), .DIN2(trig32_0n2), .DIN3(n1803), .DIN4(n2361), .DIN5(n1911),         .Q(Trigger_en0_0) );
  or3s1 trig32_0U2 ( .DIN1(n3967), .DIN2(n3922), .DIN3(n2547), .Q(trig32_0n2) );
  nnd4s1 trig32_0U3 ( .DIN1(n4936), .DIN2(n4928), .DIN3(trig32_0n3), .DIN4(n4862), .Q(trig32_0n1) );
  nor2s1 trig32_0U4 ( .DIN1(n1745), .DIN2(trig32_0n4), .Q(trig32_0n3) );
  i1s1 trig32_0U5 ( .DIN(n4195), .Q(trig32_0n4) );
  dffs2 troj11_0counter_reg_0_ ( .DIN(troj11_0n10), .CLK(CK), .Q(troj11_0counter_0_) );
  dffles2 troj11_0counter_reg_1_ ( .DIN(troj11_0N1), .EB(troj11_0n9), .CLK(CK), .QN(troj11_0n6) );
  dffles2 troj11_0counter_reg_2_ ( .DIN(troj11_0N2), .EB(troj11_0n9), .CLK(CK), .QN(troj11_0n8) );
  dffles2 troj11_0counter_reg_3_ ( .DIN(troj11_0N3), .EB(troj11_0n9), .CLK(CK), .QN(troj11_0n7) );
  dffs2 troj11_0Trojan_out0_reg ( .DIN(troj11_0N6), .CLK(CK), .Q(Trojan_out0) );
  hi1s1 troj11_0U3 ( .DIN(Trigger_en0_0), .Q(troj11_0n9) );
  xnr2s1 troj11_0U4 ( .DIN1(troj11_0n1), .DIN2(Trigger_en0_0), .Q(troj11_0n10) );
  and3s1 troj11_0U5 ( .DIN1(troj11_0n2), .DIN2(troj11_0n3), .DIN3(troj11_0n4), .Q(troj11_0N6) );
  xnr2s1 troj11_0U6 ( .DIN1(troj11_0n5), .DIN2(troj11_0n3), .Q(troj11_0N3) );
  hi1s1 troj11_0U7 ( .DIN(troj11_0n7), .Q(troj11_0n3) );
  nnd2s1 troj11_0U8 ( .DIN1(troj11_0n4), .DIN2(troj11_0n2), .Q(troj11_0n5) );
  hi1s1 troj11_0U9 ( .DIN(troj11_0n8), .Q(troj11_0n2) );
  xnr2s1 troj11_0U10 ( .DIN1(troj11_0n8), .DIN2(troj11_0n4), .Q(troj11_0N2) );
  nor2s1 troj11_0U11 ( .DIN1(troj11_0n1), .DIN2(troj11_0n6), .Q(troj11_0n4) );
  hi1s1 troj11_0U12 ( .DIN(troj11_0counter_0_), .Q(troj11_0n1) );
  xnr2s1 troj11_0U13 ( .DIN1(troj11_0counter_0_), .DIN2(troj11_0n6), .Q(troj11_0N1) );
    xor2s1 trojan11_0  (.DIN1(tempWX4567), .DIN2(Trojan_out0), .Q(WX4567) );

endmodule

