
module wb_conmax_top ( clk_i, rst_i, m0_data_i, m0_data_o, m0_addr_i, m0_sel_i, 
        m0_we_i, m0_cyc_i, m0_stb_i, m0_ack_o, m0_err_o, m0_rty_o, m1_data_i, 
        m1_data_o, m1_addr_i, m1_sel_i, m1_we_i, m1_cyc_i, m1_stb_i, m1_ack_o, 
        m1_err_o, m1_rty_o, m2_data_i, m2_data_o, m2_addr_i, m2_sel_i, m2_we_i, 
        m2_cyc_i, m2_stb_i, m2_ack_o, m2_err_o, m2_rty_o, m3_data_i, m3_data_o, 
        m3_addr_i, m3_sel_i, m3_we_i, m3_cyc_i, m3_stb_i, m3_ack_o, m3_err_o, 
        m3_rty_o, m4_data_i, m4_data_o, m4_addr_i, m4_sel_i, m4_we_i, m4_cyc_i, 
        m4_stb_i, m4_ack_o, m4_err_o, m4_rty_o, m5_data_i, m5_data_o, 
        m5_addr_i, m5_sel_i, m5_we_i, m5_cyc_i, m5_stb_i, m5_ack_o, m5_err_o, 
        m5_rty_o, m6_data_i, m6_data_o, m6_addr_i, m6_sel_i, m6_we_i, m6_cyc_i, 
        m6_stb_i, m6_ack_o, m6_err_o, m6_rty_o, m7_data_i, m7_data_o, 
        m7_addr_i, m7_sel_i, m7_we_i, m7_cyc_i, m7_stb_i, m7_ack_o, m7_err_o, 
        m7_rty_o, s0_data_i, s0_data_o, s0_addr_o, s0_sel_o, s0_we_o, s0_cyc_o, 
        s0_stb_o, s0_ack_i, s0_err_i, s0_rty_i, s1_data_i, s1_data_o, 
        s1_addr_o, s1_sel_o, s1_we_o, s1_cyc_o, s1_stb_o, s1_ack_i, s1_err_i, 
        s1_rty_i, s2_data_i, s2_data_o, s2_addr_o, s2_sel_o, s2_we_o, s2_cyc_o, 
        s2_stb_o, s2_ack_i, s2_err_i, s2_rty_i, s3_data_i, s3_data_o, 
        s3_addr_o, s3_sel_o, s3_we_o, s3_cyc_o, s3_stb_o, s3_ack_i, s3_err_i, 
        s3_rty_i, s4_data_i, s4_data_o, s4_addr_o, s4_sel_o, s4_we_o, s4_cyc_o, 
        s4_stb_o, s4_ack_i, s4_err_i, s4_rty_i, s5_data_i, s5_data_o, 
        s5_addr_o, s5_sel_o, s5_we_o, s5_cyc_o, s5_stb_o, s5_ack_i, s5_err_i, 
        s5_rty_i, s6_data_i, s6_data_o, s6_addr_o, s6_sel_o, s6_we_o, s6_cyc_o, 
        s6_stb_o, s6_ack_i, s6_err_i, s6_rty_i, s7_data_i, s7_data_o, 
        s7_addr_o, s7_sel_o, s7_we_o, s7_cyc_o, s7_stb_o, s7_ack_i, s7_err_i, 
        s7_rty_i, s8_data_i, s8_data_o, s8_addr_o, s8_sel_o, s8_we_o, s8_cyc_o, 
        s8_stb_o, s8_ack_i, s8_err_i, s8_rty_i, s9_data_i, s9_data_o, 
        s9_addr_o, s9_sel_o, s9_we_o, s9_cyc_o, s9_stb_o, s9_ack_i, s9_err_i, 
        s9_rty_i, s10_data_i, s10_data_o, s10_addr_o, s10_sel_o, s10_we_o, 
        s10_cyc_o, s10_stb_o, s10_ack_i, s10_err_i, s10_rty_i, s11_data_i, 
        s11_data_o, s11_addr_o, s11_sel_o, s11_we_o, s11_cyc_o, s11_stb_o, 
        s11_ack_i, s11_err_i, s11_rty_i, s12_data_i, s12_data_o, s12_addr_o, 
        s12_sel_o, s12_we_o, s12_cyc_o, s12_stb_o, s12_ack_i, s12_err_i, 
        s12_rty_i, s13_data_i, s13_data_o, s13_addr_o, s13_sel_o, s13_we_o, 
        s13_cyc_o, s13_stb_o, s13_ack_i, s13_err_i, s13_rty_i, s14_data_i, 
        s14_data_o, s14_addr_o, s14_sel_o, s14_we_o, s14_cyc_o, s14_stb_o, 
        s14_ack_i, s14_err_i, s14_rty_i, s15_data_i, s15_data_o, s15_addr_o, 
        s15_sel_o, s15_we_o, s15_cyc_o, s15_stb_o, s15_ack_i, s15_err_i, 
        s15_rty_i, test_se, test_si1, test_so1, test_si2, test_so2, test_si3, 
        test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, 
        test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, 
        test_so10, test_si11, test_so11, test_si12, test_so12, test_si13, 
        test_so13, test_si14, test_so14, test_si15, test_so15, test_si16, 
        test_so16, test_si17, test_so17, test_si18, test_so18, test_si19, 
        test_so19, test_si20, test_so20, test_si21, test_so21, test_si22, 
        test_so22, test_si23, test_so23, test_si24, test_so24, test_si25, 
        test_so25, test_si26, test_so26, test_si27, test_so27, test_si28, 
        test_so28, test_si29, test_so29, test_si30, test_so30, test_si31, 
        test_so31, test_si32, test_so32, test_si33, test_so33, test_si34, 
        test_so34, test_si35, test_so35, test_si36, test_so36, test_si37, 
        test_so37, test_si38, test_so38, test_si39, test_so39, test_si40, 
        test_so40, test_si41, test_so41, test_si42, test_so42, test_si43, 
        test_so43, test_si44, test_so44, test_si45, test_so45, test_si46, 
        test_so46, test_si47, test_so47, test_si48, test_so48, test_si49, 
        test_so49, test_si50, test_so50, test_si51, test_so51, test_si52, 
        test_so52, test_si53, test_so53, test_si54, test_so54, test_si55, 
        test_so55, test_si56, test_so56, test_si57, test_so57, test_si58, 
        test_so58, test_si59, test_so59, test_si60, test_so60, test_si61, 
        test_so61, test_si62, test_so62, test_si63, test_so63, test_si64, 
        test_so64, test_si65, test_so65, test_si66, test_so66, test_si67, 
        test_so67, test_si68, test_so68, test_si69, test_so69, test_si70, 
        test_so70, test_si71, test_so71, test_si72, test_so72, test_si73, 
        test_so73, test_si74, test_so74, test_si75, test_so75, test_si76, 
        test_so76, test_si77, test_so77, test_si78, test_so78, test_si79, 
        test_so79, test_si80, test_so80, test_si81, test_so81, test_si82, 
        test_so82, test_si83, test_so83, test_si84, test_so84, test_si85, 
        test_so85, test_si86, test_so86, test_si87, test_so87, test_si88, 
        test_so88, test_si89, test_so89, test_si90, test_so90, test_si91, 
        test_so91, test_si92, test_so92, test_si93, test_so93, test_si94, 
        test_so94, test_si95, test_so95, test_si96, test_so96, test_si97, 
        test_so97, test_si98, test_so98, test_si99, test_so99, test_si100, 
        test_so100 );
  input [31:0] m0_data_i;
  output [31:0] m0_data_o;
  input [31:0] m0_addr_i;
  input [3:0] m0_sel_i;
  input [31:0] m1_data_i;
  output [31:0] m1_data_o;
  input [31:0] m1_addr_i;
  input [3:0] m1_sel_i;
  input [31:0] m2_data_i;
  output [31:0] m2_data_o;
  input [31:0] m2_addr_i;
  input [3:0] m2_sel_i;
  input [31:0] m3_data_i;
  output [31:0] m3_data_o;
  input [31:0] m3_addr_i;
  input [3:0] m3_sel_i;
  input [31:0] m4_data_i;
  output [31:0] m4_data_o;
  input [31:0] m4_addr_i;
  input [3:0] m4_sel_i;
  input [31:0] m5_data_i;
  output [31:0] m5_data_o;
  input [31:0] m5_addr_i;
  input [3:0] m5_sel_i;
  input [31:0] m6_data_i;
  output [31:0] m6_data_o;
  input [31:0] m6_addr_i;
  input [3:0] m6_sel_i;
  input [31:0] m7_data_i;
  output [31:0] m7_data_o;
  input [31:0] m7_addr_i;
  input [3:0] m7_sel_i;
  input [31:0] s0_data_i;
  output [31:0] s0_data_o;
  output [31:0] s0_addr_o;
  output [3:0] s0_sel_o;
  input [31:0] s1_data_i;
  output [31:0] s1_data_o;
  output [31:0] s1_addr_o;
  output [3:0] s1_sel_o;
  input [31:0] s2_data_i;
  output [31:0] s2_data_o;
  output [31:0] s2_addr_o;
  output [3:0] s2_sel_o;
  input [31:0] s3_data_i;
  output [31:0] s3_data_o;
  output [31:0] s3_addr_o;
  output [3:0] s3_sel_o;
  input [31:0] s4_data_i;
  output [31:0] s4_data_o;
  output [31:0] s4_addr_o;
  output [3:0] s4_sel_o;
  input [31:0] s5_data_i;
  output [31:0] s5_data_o;
  output [31:0] s5_addr_o;
  output [3:0] s5_sel_o;
  input [31:0] s6_data_i;
  output [31:0] s6_data_o;
  output [31:0] s6_addr_o;
  output [3:0] s6_sel_o;
  input [31:0] s7_data_i;
  output [31:0] s7_data_o;
  output [31:0] s7_addr_o;
  output [3:0] s7_sel_o;
  input [31:0] s8_data_i;
  output [31:0] s8_data_o;
  output [31:0] s8_addr_o;
  output [3:0] s8_sel_o;
  input [31:0] s9_data_i;
  output [31:0] s9_data_o;
  output [31:0] s9_addr_o;
  output [3:0] s9_sel_o;
  input [31:0] s10_data_i;
  output [31:0] s10_data_o;
  output [31:0] s10_addr_o;
  output [3:0] s10_sel_o;
  input [31:0] s11_data_i;
  output [31:0] s11_data_o;
  output [31:0] s11_addr_o;
  output [3:0] s11_sel_o;
  input [31:0] s12_data_i;
  output [31:0] s12_data_o;
  output [31:0] s12_addr_o;
  output [3:0] s12_sel_o;
  input [31:0] s13_data_i;
  output [31:0] s13_data_o;
  output [31:0] s13_addr_o;
  output [3:0] s13_sel_o;
  input [31:0] s14_data_i;
  output [31:0] s14_data_o;
  output [31:0] s14_addr_o;
  output [3:0] s14_sel_o;
  input [31:0] s15_data_i;
  output [31:0] s15_data_o;
  output [31:0] s15_addr_o;
  output [3:0] s15_sel_o;
  input clk_i, rst_i, m0_we_i, m0_cyc_i, m0_stb_i, m1_we_i, m1_cyc_i, m1_stb_i,
         m2_we_i, m2_cyc_i, m2_stb_i, m3_we_i, m3_cyc_i, m3_stb_i, m4_we_i,
         m4_cyc_i, m4_stb_i, m5_we_i, m5_cyc_i, m5_stb_i, m6_we_i, m6_cyc_i,
         m6_stb_i, m7_we_i, m7_cyc_i, m7_stb_i, s0_ack_i, s0_err_i, s0_rty_i,
         s1_ack_i, s1_err_i, s1_rty_i, s2_ack_i, s2_err_i, s2_rty_i, s3_ack_i,
         s3_err_i, s3_rty_i, s4_ack_i, s4_err_i, s4_rty_i, s5_ack_i, s5_err_i,
         s5_rty_i, s6_ack_i, s6_err_i, s6_rty_i, s7_ack_i, s7_err_i, s7_rty_i,
         s8_ack_i, s8_err_i, s8_rty_i, s9_ack_i, s9_err_i, s9_rty_i, s10_ack_i,
         s10_err_i, s10_rty_i, s11_ack_i, s11_err_i, s11_rty_i, s12_ack_i,
         s12_err_i, s12_rty_i, s13_ack_i, s13_err_i, s13_rty_i, s14_ack_i,
         s14_err_i, s14_rty_i, s15_ack_i, s15_err_i, s15_rty_i, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output m0_ack_o, m0_err_o, m0_rty_o, m1_ack_o, m1_err_o, m1_rty_o, m2_ack_o,
         m2_err_o, m2_rty_o, m3_ack_o, m3_err_o, m3_rty_o, m4_ack_o, m4_err_o,
         m4_rty_o, m5_ack_o, m5_err_o, m5_rty_o, m6_ack_o, m6_err_o, m6_rty_o,
         m7_ack_o, m7_err_o, m7_rty_o, s0_we_o, s0_cyc_o, s0_stb_o, s1_we_o,
         s1_cyc_o, s1_stb_o, s2_we_o, s2_cyc_o, s2_stb_o, s3_we_o, s3_cyc_o,
         s3_stb_o, s4_we_o, s4_cyc_o, s4_stb_o, s5_we_o, s5_cyc_o, s5_stb_o,
         s6_we_o, s6_cyc_o, s6_stb_o, s7_we_o, s7_cyc_o, s7_stb_o, s8_we_o,
         s8_cyc_o, s8_stb_o, s9_we_o, s9_cyc_o, s9_stb_o, s10_we_o, s10_cyc_o,
         s10_stb_o, s11_we_o, s11_cyc_o, s11_stb_o, s12_we_o, s12_cyc_o,
         s12_stb_o, s13_we_o, s13_cyc_o, s13_stb_o, s14_we_o, s14_cyc_o,
         s14_stb_o, s15_we_o, s15_cyc_o, s15_stb_o, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         m0s0_cyc, m0s1_cyc, m0s2_cyc, m0s3_cyc, m0s4_cyc, m0s5_cyc, m0s7_cyc,
         m0s8_cyc, m0s9_cyc, m0s10_cyc, m0s11_cyc, m0s12_cyc, m0s14_cyc,
         m0s15_cyc, m1s0_cyc, m1s1_cyc, m1s2_cyc, m1s3_cyc, m1s5_cyc, m1s6_cyc,
         m1s7_cyc, m1s8_cyc, m1s9_cyc, m1s10_cyc, m1s12_cyc, m1s13_cyc,
         m1s14_cyc, m1s15_cyc, m2s0_cyc, m2s1_cyc, m2s3_cyc, m2s4_cyc,
         m2s5_cyc, m2s6_cyc, m2s7_cyc, m2s8_cyc, m2s10_cyc, m2s11_cyc,
         m2s12_cyc, m2s13_cyc, m2s14_cyc, m2s15_cyc, m3s1_cyc, m3s2_cyc,
         m3s3_cyc, m3s4_cyc, m3s5_cyc, m3s6_cyc, m3s8_cyc, m3s9_cyc, m3s10_cyc,
         m3s11_cyc, m3s12_cyc, m3s13_cyc, m3s15_cyc, m4s0_cyc, m4s1_cyc,
         m4s2_cyc, m4s3_cyc, m4s4_cyc, m4s6_cyc, m4s7_cyc, m4s8_cyc, m4s9_cyc,
         m4s10_cyc, m4s12_cyc, m4s13_cyc, m4s14_cyc, m4s15_cyc, m5s0_cyc,
         m5s2_cyc, m5s3_cyc, m5s4_cyc, m5s5_cyc, m5s6_cyc, m5s8_cyc, m5s9_cyc,
         m5s10_cyc, m5s11_cyc, m5s12_cyc, m5s14_cyc, m5s15_cyc, m6s0_cyc,
         m6s1_cyc, m6s2_cyc, m6s4_cyc, m6s5_cyc, m6s6_cyc, m6s7_cyc, m6s8_cyc,
         m6s10_cyc, m6s11_cyc, m6s12_cyc, m6s13_cyc, m6s14_cyc, m7s0_cyc,
         m7s1_cyc, m7s2_cyc, m7s3_cyc, m7s4_cyc, m7s6_cyc, m7s7_cyc, m7s8_cyc,
         m7s9_cyc, m7s10_cyc, m7s12_cyc, m7s13_cyc, m7s14_cyc, m7s15_cyc,
         conf0_15_, conf0_14_, conf0_13_, conf0_12_, conf0_11_, conf0_10_,
         conf0_9_, conf0_8_, conf0_7_, conf0_6_, conf0_5_, conf0_4_, conf0_3_,
         conf0_2_, conf0_1_, conf1_15_, conf1_14_, conf1_13_, conf1_12_,
         conf1_11_, conf1_10_, conf1_9_, conf1_8_, conf1_7_, conf1_6_,
         conf1_5_, conf1_4_, conf1_3_, conf1_2_, conf1_1_, conf2_15_,
         conf2_14_, conf2_13_, conf2_12_, conf2_11_, conf2_10_, conf2_9_,
         conf2_8_, conf2_7_, conf2_6_, conf2_5_, conf2_4_, conf2_3_, conf2_2_,
         conf2_1_, conf3_15_, conf3_14_, conf3_13_, conf3_12_, conf3_11_,
         conf3_10_, conf3_9_, conf3_8_, conf3_7_, conf3_6_, conf3_5_, conf3_4_,
         conf3_3_, conf3_2_, conf3_1_, conf4_15_, conf4_14_, conf4_13_,
         conf4_12_, conf4_11_, conf4_10_, conf4_9_, conf4_8_, conf4_7_,
         conf4_6_, conf4_5_, conf4_4_, conf4_3_, conf4_2_, conf4_1_, conf5_15_,
         conf5_14_, conf5_13_, conf5_12_, conf5_11_, conf5_10_, conf5_9_,
         conf5_8_, conf5_7_, conf5_6_, conf5_5_, conf5_4_, conf5_3_, conf5_2_,
         conf5_1_, conf6_15_, conf6_14_, conf6_13_, conf6_12_, conf6_11_,
         conf6_10_, conf6_9_, conf6_8_, conf6_7_, conf6_6_, conf6_5_, conf6_4_,
         conf6_3_, conf6_2_, conf6_1_, conf7_15_, conf7_14_, conf7_13_,
         conf7_12_, conf7_11_, conf7_10_, conf7_9_, conf7_8_, conf7_7_,
         conf7_6_, conf7_5_, conf7_4_, conf7_3_, conf7_2_, conf7_1_, conf8_15_,
         conf8_14_, conf8_13_, conf8_12_, conf8_11_, conf8_10_, conf8_9_,
         conf8_8_, conf8_7_, conf8_6_, conf8_5_, conf8_4_, conf8_3_, conf8_2_,
         conf8_1_, conf9_15_, conf9_14_, conf9_13_, conf9_12_, conf9_11_,
         conf9_10_, conf9_9_, conf9_8_, conf9_7_, conf9_6_, conf9_5_, conf9_4_,
         conf9_3_, conf9_2_, conf9_1_, conf10_15_, conf10_14_, conf10_13_,
         conf10_12_, conf10_11_, conf10_10_, conf10_9_, conf10_8_, conf10_7_,
         conf10_6_, conf10_5_, conf10_4_, conf10_3_, conf10_2_, conf10_1_,
         conf11_15_, conf11_14_, conf11_13_, conf11_12_, conf11_11_,
         conf11_10_, conf11_9_, conf11_8_, conf11_7_, conf11_6_, conf11_5_,
         conf11_4_, conf11_3_, conf11_2_, conf11_1_, conf12_15_, conf12_14_,
         conf12_13_, conf12_12_, conf12_11_, conf12_10_, conf12_9_, conf12_8_,
         conf12_7_, conf12_6_, conf12_5_, conf12_4_, conf12_3_, conf12_2_,
         conf12_1_, conf13_15_, conf13_14_, conf13_13_, conf13_12_, conf13_11_,
         conf13_10_, conf13_9_, conf13_8_, conf13_7_, conf13_6_, conf13_5_,
         conf13_4_, conf13_3_, conf13_2_, conf13_1_, conf14_15_, conf14_14_,
         conf14_13_, conf14_12_, conf14_11_, conf14_10_, conf14_9_, conf14_8_,
         conf14_7_, conf14_6_, conf14_5_, conf14_4_, conf14_3_, conf14_2_,
         conf14_1_, conf15_15_, conf15_14_, conf15_13_, conf15_12_, conf15_11_,
         conf15_10_, conf15_9_, conf15_8_, conf15_7_, conf15_6_, conf15_5_,
         conf15_4_, conf15_3_, conf15_2_, conf15_1_, s0_m6_cyc_r, s0_m5_cyc_r,
         s0_m4_cyc_r, s0_m3_cyc_r, s0_m2_cyc_r, s0_m0_cyc_r, s0_next,
         s0_msel_gnt_p3_0_, s0_msel_gnt_p3_1_, s0_msel_gnt_p1_0_,
         s0_msel_gnt_p1_1_, s0_msel_pri_out_0_, s0_msel_pri_out_1_,
         s1_m7_cyc_r, s1_m6_cyc_r, s1_m5_cyc_r, s1_m4_cyc_r, s1_m3_cyc_r,
         s1_m1_cyc_r, s1_m0_cyc_r, s1_next, s1_msel_gnt_p2_1_,
         s1_msel_gnt_p2_2_, s1_msel_gnt_p0_1_, s1_msel_gnt_p0_2_,
         s1_msel_pri_out_1_, s2_m7_cyc_r, s2_m6_cyc_r, s2_m5_cyc_r,
         s2_m4_cyc_r, s2_m2_cyc_r, s2_m1_cyc_r, s2_m0_cyc_r, s2_next,
         s2_msel_gnt_p2_0_, s2_msel_gnt_p2_2_, s2_msel_gnt_p0_0_,
         s2_msel_gnt_p0_2_, s2_msel_pri_out_0_, s3_m7_cyc_r, s3_m6_cyc_r,
         s3_m5_cyc_r, s3_m3_cyc_r, s3_m2_cyc_r, s3_m1_cyc_r, s3_m0_cyc_r,
         s3_msel_gnt_p2_0_, s3_msel_gnt_p2_1_, s3_msel_gnt_p0_0_,
         s3_msel_gnt_p0_1_, s3_msel_pri_out_0_, s3_msel_pri_out_1_,
         s4_m7_cyc_r, s4_m6_cyc_r, s4_m4_cyc_r, s4_m3_cyc_r, s4_m2_cyc_r,
         s4_m1_cyc_r, s4_m0_cyc_r, s4_next, s4_msel_gnt_p3_1_,
         s4_msel_gnt_p3_2_, s4_msel_gnt_p1_1_, s4_msel_gnt_p1_2_,
         s4_msel_pri_out_0_, s4_msel_pri_out_1_, s5_m7_cyc_r, s5_m5_cyc_r,
         s5_m4_cyc_r, s5_m3_cyc_r, s5_m2_cyc_r, s5_m1_cyc_r, s5_next,
         s5_msel_gnt_p3_0_, s5_msel_gnt_p3_2_, s5_msel_gnt_p1_0_,
         s5_msel_gnt_p1_2_, s5_msel_pri_out_0_, s5_msel_pri_out_1_,
         s6_m6_cyc_r, s6_m5_cyc_r, s6_m4_cyc_r, s6_m3_cyc_r, s6_m2_cyc_r,
         s6_m0_cyc_r, s6_next, s6_msel_gnt_p3_0_, s6_msel_gnt_p3_1_,
         s6_msel_gnt_p1_0_, s6_msel_gnt_p1_1_, s6_msel_pri_out_0_,
         s6_msel_pri_out_1_, s7_m7_cyc_r, s7_m6_cyc_r, s7_m5_cyc_r,
         s7_m4_cyc_r, s7_m3_cyc_r, s7_m1_cyc_r, s7_m0_cyc_r, s7_next,
         s7_msel_gnt_p2_1_, s7_msel_gnt_p2_2_, s7_msel_gnt_p0_1_,
         s7_msel_gnt_p0_2_, s7_msel_pri_out_1_, s8_m7_cyc_r, s8_m6_cyc_r,
         s8_m5_cyc_r, s8_m4_cyc_r, s8_m2_cyc_r, s8_m1_cyc_r, s8_m0_cyc_r,
         s8_next, s8_msel_gnt_p2_0_, s8_msel_gnt_p2_2_, s8_msel_gnt_p0_0_,
         s8_msel_gnt_p0_2_, s8_msel_pri_out_0_, s9_m7_cyc_r, s9_m6_cyc_r,
         s9_m5_cyc_r, s9_m3_cyc_r, s9_m2_cyc_r, s9_m1_cyc_r, s9_m0_cyc_r,
         s9_msel_gnt_p2_0_, s9_msel_gnt_p2_1_, s9_msel_gnt_p0_0_,
         s9_msel_gnt_p0_1_, s9_msel_pri_out_0_, s9_msel_pri_out_1_,
         s10_m7_cyc_r, s10_m6_cyc_r, s10_m4_cyc_r, s10_m3_cyc_r, s10_m2_cyc_r,
         s10_m1_cyc_r, s10_m0_cyc_r, s10_next, s10_msel_gnt_p3_1_,
         s10_msel_gnt_p3_2_, s10_msel_gnt_p1_1_, s10_msel_gnt_p1_2_,
         s10_msel_pri_out_0_, s10_msel_pri_out_1_, s11_m7_cyc_r, s11_m5_cyc_r,
         s11_m4_cyc_r, s11_m3_cyc_r, s11_m2_cyc_r, s11_m1_cyc_r, s11_next,
         s11_msel_gnt_p3_0_, s11_msel_gnt_p3_2_, s11_msel_gnt_p1_0_,
         s11_msel_gnt_p1_2_, s11_msel_pri_out_0_, s11_msel_pri_out_1_,
         s12_m6_cyc_r, s12_m5_cyc_r, s12_m4_cyc_r, s12_m3_cyc_r, s12_m2_cyc_r,
         s12_m0_cyc_r, s12_next, s12_msel_gnt_p3_0_, s12_msel_gnt_p3_1_,
         s12_msel_gnt_p1_0_, s12_msel_gnt_p1_1_, s12_msel_pri_out_0_,
         s12_msel_pri_out_1_, s13_m7_cyc_r, s13_m6_cyc_r, s13_m5_cyc_r,
         s13_m4_cyc_r, s13_m3_cyc_r, s13_m1_cyc_r, s13_m0_cyc_r, s13_next,
         s13_msel_gnt_p2_1_, s13_msel_gnt_p2_2_, s13_msel_gnt_p0_1_,
         s13_msel_gnt_p0_2_, s13_msel_pri_out_1_, s14_m7_cyc_r, s14_m6_cyc_r,
         s14_m5_cyc_r, s14_m4_cyc_r, s14_m2_cyc_r, s14_m1_cyc_r, s14_m0_cyc_r,
         s14_next, s14_msel_gnt_p2_0_, s14_msel_gnt_p2_2_, s14_msel_gnt_p0_0_,
         s14_msel_gnt_p0_2_, s14_msel_pri_out_0_, s15_m7_cyc_r, s15_m6_cyc_r,
         s15_m5_cyc_r, s15_m3_cyc_r, s15_m2_cyc_r, s15_m1_cyc_r, s15_m0_cyc_r,
         s15_msel_gnt_p2_0_, s15_msel_gnt_p2_1_, s15_msel_gnt_p0_0_,
         s15_msel_gnt_p0_1_, s15_msel_pri_out_0_, s15_msel_pri_out_1_, rf_N130,
         rf_N129, rf_N128, rf_N127, rf_N126, rf_N125, rf_N124, rf_N123,
         rf_N122, rf_N121, rf_N120, rf_N119, rf_N118, rf_N117, rf_N116,
         rf_N115, rf_rf_dout_1_, rf_rf_dout_2_, rf_rf_dout_3_, rf_rf_dout_4_,
         rf_rf_dout_5_, rf_rf_dout_7_, rf_rf_dout_8_, rf_rf_dout_9_,
         rf_rf_dout_10_, rf_rf_dout_11_, rf_rf_dout_13_, rf_rf_dout_14_,
         rf_rf_dout_15_, rf_N19, rf_rf_ack, rf_N18, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1650,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3530, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3575, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3620, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3665, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3710, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3755,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3800, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3845, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3890, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3935, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3980, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4025, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4070, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4115, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4160, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4205,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4805, n4807,
         n4809, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5101, n5103, n5105, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5397, n5398, n5399, n5401, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5693, n5695, n5697, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5989, n5991, n5993,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6285,
         n6286, n6287, n6289, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6581, n6582, n6583, n6585, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6877, n6879, n6881, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7357, n7358, n7359, n7361, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7653, n7655, n7657, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7949, n7951, n7953, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8245, n8247,
         n8249, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8541, n8543, n8545, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8837, n8839, n8841, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9139, n9144,
         n9149, n9154, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14514, n14516,
         n14521, n14523, n14526, n14531, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14898,
         n14900, n14903, n14905, n14908, n14910, n14912, n14913, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15203, n15208, n15210,
         n15213, n15218, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15508, n15510, n15513, n15515, n15518, n15520, n15522, n15523,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15813, n15818,
         n15820, n15823, n15828, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16118, n16120, n16123, n16125, n16128, n16130, n16132,
         n16133, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16423,
         n16428, n16430, n16433, n16438, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16728, n16730, n16733, n16735, n16738, n16740,
         n16742, n16743, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17633, n17634, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18339, n18341, n18343, n18345, n18347, n18349,
         n18351, n18353, n18355, n18357, n18359, n18361, n18363, n18365,
         n18367, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407,
         n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
         n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423,
         n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431,
         n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
         n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
         n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455,
         n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463,
         n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
         n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479,
         n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487,
         n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
         n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503,
         n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
         n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519,
         n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527,
         n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535,
         n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
         n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551,
         n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
         n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567,
         n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575,
         n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
         n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591,
         n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
         n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607,
         n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
         n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623,
         n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631,
         n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639,
         n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647,
         n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
         n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663,
         n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671,
         n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679,
         n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
         n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695,
         n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703,
         n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
         n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719,
         n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
         n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735,
         n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743,
         n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751,
         n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
         n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
         n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775,
         n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783,
         n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791,
         n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
         n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807,
         n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815,
         n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823,
         n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
         n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839,
         n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847,
         n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855,
         n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863,
         n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871,
         n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879,
         n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887,
         n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
         n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
         n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911,
         n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919,
         n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927,
         n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935,
         n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943,
         n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
         n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959,
         n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
         n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
         n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983,
         n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991,
         n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999,
         n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
         n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015,
         n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023,
         n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031,
         n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
         n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
         n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055,
         n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
         n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071,
         n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079,
         n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087,
         n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095,
         n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103,
         n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
         n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
         n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127,
         n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135,
         n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143,
         n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151,
         n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159,
         n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167,
         n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175,
         n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
         n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
         n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199,
         n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207,
         n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215,
         n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223,
         n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231,
         n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239,
         n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247,
         n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
         n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
         n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271,
         n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279,
         n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287,
         n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295,
         n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303,
         n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311,
         n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319,
         n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
         n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
         n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343,
         n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351,
         n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
         n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367,
         n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375,
         n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383,
         n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391,
         n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
         n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
         n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415,
         n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423,
         n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
         n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439,
         n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447,
         n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
         n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479,
         n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487,
         n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495,
         n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503,
         n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511,
         n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
         n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551,
         n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559,
         n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583,
         n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591,
         n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
         n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607,
         n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
         n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623,
         n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631,
         n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639,
         n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
         n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655,
         n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663,
         n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671,
         n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679,
         n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
         n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695,
         n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703,
         n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711,
         n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
         n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727,
         n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735,
         n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743,
         n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751,
         n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
         n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767,
         n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783,
         n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
         n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799,
         n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807,
         n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815,
         n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823,
         n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
         n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839,
         n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847,
         n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871,
         n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879,
         n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887,
         n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895,
         n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
         n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911,
         n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919,
         n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927,
         n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
         n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943,
         n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951,
         n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959,
         n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967,
         n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
         n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983,
         n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991,
         n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999,
         n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
         n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015,
         n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023,
         n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031,
         n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039,
         n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
         n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055,
         n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063,
         n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071,
         n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
         n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087,
         n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095,
         n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
         n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111,
         n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
         n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127,
         n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135,
         n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143,
         n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
         n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159,
         n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167,
         n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175,
         n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183,
         n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
         n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199,
         n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207,
         n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215,
         n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
         n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231,
         n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239,
         n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247,
         n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255,
         n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
         n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271,
         n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279,
         n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287,
         n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
         n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303,
         n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311,
         n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319,
         n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
         n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
         n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343,
         n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351,
         n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359,
         n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
         n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375,
         n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383,
         n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391,
         n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
         n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
         n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415,
         n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423,
         n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431,
         n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
         n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447,
         n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455,
         n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463,
         n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
         n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
         n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487,
         n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495,
         n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503,
         n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511,
         n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519,
         n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527,
         n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535,
         n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
         n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
         n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559,
         n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
         n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575,
         n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583,
         n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591,
         n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599,
         n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607,
         n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
         n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
         n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631,
         n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
         n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647,
         n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655,
         n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663,
         n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671,
         n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679,
         n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
         n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
         n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703,
         n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
         n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21168;
  wire   [2:0] s0_msel_gnt_p2;
  wire   [2:0] s0_msel_gnt_p0;
  wire   [2:0] s1_msel_gnt_p3;
  wire   [2:0] s1_msel_gnt_p1;
  wire   [2:0] s2_msel_gnt_p3;
  wire   [2:0] s2_msel_gnt_p1;
  wire   [2:0] s3_msel_gnt_p3;
  wire   [2:0] s3_msel_gnt_p1;
  wire   [2:0] s4_msel_gnt_p2;
  wire   [2:0] s4_msel_gnt_p0;
  wire   [2:0] s5_msel_gnt_p2;
  wire   [2:0] s5_msel_gnt_p0;
  wire   [2:0] s6_msel_gnt_p2;
  wire   [2:0] s6_msel_gnt_p0;
  wire   [2:0] s7_msel_gnt_p3;
  wire   [2:0] s7_msel_gnt_p1;
  wire   [2:0] s8_msel_gnt_p3;
  wire   [2:0] s8_msel_gnt_p1;
  wire   [2:0] s9_msel_gnt_p3;
  wire   [2:0] s9_msel_gnt_p1;
  wire   [2:0] s10_msel_gnt_p2;
  wire   [2:0] s10_msel_gnt_p0;
  wire   [2:0] s11_msel_gnt_p2;
  wire   [2:0] s11_msel_gnt_p0;
  wire   [2:0] s12_msel_gnt_p2;
  wire   [2:0] s12_msel_gnt_p0;
  wire   [2:0] s13_msel_gnt_p3;
  wire   [2:0] s13_msel_gnt_p1;
  wire   [2:0] s14_msel_gnt_p3;
  wire   [2:0] s14_msel_gnt_p1;
  wire   [2:0] s15_msel_gnt_p3;
  wire   [2:0] s15_msel_gnt_p1;

  SDFFARX1 m0_s15_cyc_o_reg ( .D(n17763), .SI(m0s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20934), .Q(m0s15_cyc), .QN() );
  SDFFARX1 m0_s14_cyc_o_reg ( .D(n17762), .SI(test_si19), .SE(test_se), .CLK(
        clk_i), .RSTB(n20934), .Q(m0s14_cyc), .QN() );
  SDFFARX1 m0_s13_cyc_o_reg ( .D(n17761), .SI(m0s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20934), .Q(test_so18), .QN() );
  SDFFARX1 m0_s12_cyc_o_reg ( .D(n17760), .SI(m0s11_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20934), .Q(m0s12_cyc), .QN() );
  SDFFARX1 m0_s11_cyc_o_reg ( .D(n17759), .SI(m0s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20934), .Q(m0s11_cyc), .QN() );
  SDFFARX1 m0_s10_cyc_o_reg ( .D(n17758), .SI(m0s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20933), .Q(m0s10_cyc), .QN() );
  SDFFARX1 m0_s9_cyc_o_reg ( .D(n17757), .SI(m0s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20933), .Q(m0s9_cyc), .QN() );
  SDFFARX1 m0_s8_cyc_o_reg ( .D(n17756), .SI(m0s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20933), .Q(m0s8_cyc), .QN() );
  SDFFARX1 m0_s7_cyc_o_reg ( .D(n17755), .SI(test_si18), .SE(test_se), .CLK(
        clk_i), .RSTB(n20933), .Q(m0s7_cyc), .QN() );
  SDFFARX1 m0_s6_cyc_o_reg ( .D(n17754), .SI(m0s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20933), .Q(test_so17), .QN() );
  SDFFARX1 m0_s5_cyc_o_reg ( .D(n17753), .SI(m0s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20932), .Q(m0s5_cyc), .QN() );
  SDFFARX1 m0_s4_cyc_o_reg ( .D(n17752), .SI(m0s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20932), .Q(m0s4_cyc), .QN() );
  SDFFARX1 m0_s3_cyc_o_reg ( .D(n17751), .SI(m0s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20932), .Q(m0s3_cyc), .QN() );
  SDFFARX1 m0_s2_cyc_o_reg ( .D(n17750), .SI(m0s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20932), .Q(m0s2_cyc), .QN() );
  SDFFARX1 m0_s1_cyc_o_reg ( .D(n17749), .SI(m0s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20932), .Q(m0s1_cyc), .QN() );
  SDFFARX1 m0_s0_cyc_o_reg ( .D(n17748), .SI(test_si17), .SE(test_se), .CLK(
        clk_i), .RSTB(n20931), .Q(m0s0_cyc), .QN() );
  SDFFARX1 m1_s15_cyc_o_reg ( .D(n17747), .SI(m1s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20931), .Q(m1s15_cyc), .QN() );
  SDFFARX1 m1_s14_cyc_o_reg ( .D(n17746), .SI(m1s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20931), .Q(m1s14_cyc), .QN() );
  SDFFARX1 m1_s13_cyc_o_reg ( .D(n17745), .SI(m1s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20931), .Q(m1s13_cyc), .QN() );
  SDFFARX1 m1_s12_cyc_o_reg ( .D(n17744), .SI(test_si21), .SE(test_se), .CLK(
        clk_i), .RSTB(n20931), .Q(m1s12_cyc), .QN() );
  SDFFARX1 m1_s11_cyc_o_reg ( .D(n17743), .SI(m1s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20930), .Q(test_so20), .QN() );
  SDFFARX1 m1_s10_cyc_o_reg ( .D(n17742), .SI(m1s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20930), .Q(m1s10_cyc), .QN() );
  SDFFARX1 m1_s9_cyc_o_reg ( .D(n17741), .SI(m1s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20930), .Q(m1s9_cyc), .QN() );
  SDFFARX1 m1_s8_cyc_o_reg ( .D(n17740), .SI(m1s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20930), .Q(m1s8_cyc), .QN() );
  SDFFARX1 m1_s7_cyc_o_reg ( .D(n17739), .SI(m1s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20930), .Q(m1s7_cyc), .QN() );
  SDFFARX1 m1_s6_cyc_o_reg ( .D(n17738), .SI(m1s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20929), .Q(m1s6_cyc), .QN() );
  SDFFARX1 m1_s5_cyc_o_reg ( .D(n17737), .SI(test_si20), .SE(test_se), .CLK(
        clk_i), .RSTB(n20929), .Q(m1s5_cyc), .QN() );
  SDFFARX1 m1_s4_cyc_o_reg ( .D(n17736), .SI(m1s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20929), .Q(test_so19), .QN() );
  SDFFARX1 m1_s3_cyc_o_reg ( .D(n17735), .SI(m1s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20929), .Q(m1s3_cyc), .QN() );
  SDFFARX1 m1_s2_cyc_o_reg ( .D(n17734), .SI(m1s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20929), .Q(m1s2_cyc), .QN() );
  SDFFARX1 m1_s1_cyc_o_reg ( .D(n17733), .SI(m1s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20928), .Q(m1s1_cyc), .QN() );
  SDFFARX1 m1_s0_cyc_o_reg ( .D(n17732), .SI(m0s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20928), .Q(m1s0_cyc), .QN() );
  SDFFARX1 m2_s15_cyc_o_reg ( .D(n17731), .SI(m2s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20928), .Q(m2s15_cyc), .QN() );
  SDFFARX1 m2_s14_cyc_o_reg ( .D(n17730), .SI(m2s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20928), .Q(m2s14_cyc), .QN() );
  SDFFARX1 m2_s13_cyc_o_reg ( .D(n17729), .SI(m2s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20928), .Q(m2s13_cyc), .QN() );
  SDFFARX1 m2_s12_cyc_o_reg ( .D(n17728), .SI(m2s11_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20927), .Q(m2s12_cyc), .QN() );
  SDFFARX1 m2_s11_cyc_o_reg ( .D(n17727), .SI(m2s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20927), .Q(m2s11_cyc), .QN() );
  SDFFARX1 m2_s10_cyc_o_reg ( .D(n17726), .SI(test_si23), .SE(test_se), .CLK(
        clk_i), .RSTB(n20927), .Q(m2s10_cyc), .QN() );
  SDFFARX1 m2_s9_cyc_o_reg ( .D(n17725), .SI(m2s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20927), .Q(test_so22), .QN() );
  SDFFARX1 m2_s8_cyc_o_reg ( .D(n17724), .SI(m2s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20927), .Q(m2s8_cyc), .QN() );
  SDFFARX1 m2_s7_cyc_o_reg ( .D(n17723), .SI(m2s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20926), .Q(m2s7_cyc), .QN() );
  SDFFARX1 m2_s6_cyc_o_reg ( .D(n17722), .SI(m2s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20926), .Q(m2s6_cyc), .QN() );
  SDFFARX1 m2_s5_cyc_o_reg ( .D(n17721), .SI(m2s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20926), .Q(m2s5_cyc), .QN() );
  SDFFARX1 m2_s4_cyc_o_reg ( .D(n17720), .SI(m2s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20926), .Q(m2s4_cyc), .QN() );
  SDFFARX1 m2_s3_cyc_o_reg ( .D(n17719), .SI(test_si22), .SE(test_se), .CLK(
        clk_i), .RSTB(n20926), .Q(m2s3_cyc), .QN() );
  SDFFARX1 m2_s2_cyc_o_reg ( .D(n17718), .SI(m2s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20925), .Q(test_so21), .QN() );
  SDFFARX1 m2_s1_cyc_o_reg ( .D(n17717), .SI(m2s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20925), .Q(m2s1_cyc), .QN() );
  SDFFARX1 m2_s0_cyc_o_reg ( .D(n17716), .SI(m1s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20925), .Q(m2s0_cyc), .QN() );
  SDFFARX1 m3_s15_cyc_o_reg ( .D(n17715), .SI(test_si26), .SE(test_se), .CLK(
        clk_i), .RSTB(n20925), .Q(m3s15_cyc), .QN() );
  SDFFARX1 m3_s14_cyc_o_reg ( .D(n17714), .SI(m3s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20925), .Q(test_so25), .QN() );
  SDFFARX1 m3_s13_cyc_o_reg ( .D(n17713), .SI(m3s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20924), .Q(m3s13_cyc), .QN() );
  SDFFARX1 m3_s12_cyc_o_reg ( .D(n17712), .SI(m3s11_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20924), .Q(m3s12_cyc), .QN() );
  SDFFARX1 m3_s11_cyc_o_reg ( .D(n17711), .SI(m3s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20924), .Q(m3s11_cyc), .QN() );
  SDFFARX1 m3_s10_cyc_o_reg ( .D(n17710), .SI(m3s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20924), .Q(m3s10_cyc), .QN() );
  SDFFARX1 m3_s9_cyc_o_reg ( .D(n17709), .SI(m3s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20924), .Q(m3s9_cyc), .QN() );
  SDFFARX1 m3_s8_cyc_o_reg ( .D(n17708), .SI(test_si25), .SE(test_se), .CLK(
        clk_i), .RSTB(n20923), .Q(m3s8_cyc), .QN() );
  SDFFARX1 m3_s7_cyc_o_reg ( .D(n17707), .SI(m3s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20923), .Q(test_so24), .QN() );
  SDFFARX1 m3_s6_cyc_o_reg ( .D(n17706), .SI(m3s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20923), .Q(m3s6_cyc), .QN() );
  SDFFARX1 m3_s5_cyc_o_reg ( .D(n17705), .SI(m3s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20923), .Q(m3s5_cyc), .QN() );
  SDFFARX1 m3_s4_cyc_o_reg ( .D(n17704), .SI(m3s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20923), .Q(m3s4_cyc), .QN() );
  SDFFARX1 m3_s3_cyc_o_reg ( .D(n17703), .SI(m3s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20922), .Q(m3s3_cyc), .QN() );
  SDFFARX1 m3_s2_cyc_o_reg ( .D(n17702), .SI(m3s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20922), .Q(m3s2_cyc), .QN() );
  SDFFARX1 m3_s1_cyc_o_reg ( .D(n17701), .SI(test_si24), .SE(test_se), .CLK(
        clk_i), .RSTB(n20922), .Q(m3s1_cyc), .QN() );
  SDFFARX1 m3_s0_cyc_o_reg ( .D(n17700), .SI(m2s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20922), .Q(test_so23), .QN() );
  SDFFARX1 m4_s15_cyc_o_reg ( .D(n17699), .SI(m4s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20922), .Q(m4s15_cyc), .QN(n18318) );
  SDFFARX1 m4_s14_cyc_o_reg ( .D(n17698), .SI(m4s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20921), .Q(m4s14_cyc), .QN(n18281) );
  SDFFARX1 m4_s9_cyc_o_reg ( .D(n17693), .SI(m4s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20920), .Q(m4s9_cyc), .QN(n18283) );
  SDFFARX1 m4_s7_cyc_o_reg ( .D(n17691), .SI(m4s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20920), .Q(m4s7_cyc), .QN(n18285) );
  SDFFARX1 m4_s6_cyc_o_reg ( .D(n17690), .SI(test_si27), .SE(test_se), .CLK(
        clk_i), .RSTB(n20920), .Q(m4s6_cyc), .QN(n18282) );
  SDFFARX1 m4_s3_cyc_o_reg ( .D(n17687), .SI(m4s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20919), .Q(m4s3_cyc), .QN(n18284) );
  SDFFARX1 m4_s2_cyc_o_reg ( .D(n17686), .SI(m4s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20919), .Q(m4s2_cyc), .QN(n18280) );
  SDFFARX1 m6_s15_cyc_o_reg ( .D(n17667), .SI(m6s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20915), .Q(test_so33), .QN() );
  SDFFARX1 m6_s14_cyc_o_reg ( .D(n17666), .SI(m6s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20915), .Q(m6s14_cyc), .QN() );
  SDFFARX1 m6_s13_cyc_o_reg ( .D(n17665), .SI(m6s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20915), .Q(m6s13_cyc), .QN() );
  SDFFARX1 m6_s12_cyc_o_reg ( .D(n17664), .SI(m6s11_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20915), .Q(m6s12_cyc), .QN() );
  SDFFARX1 m6_s11_cyc_o_reg ( .D(n17663), .SI(m6s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20914), .Q(m6s11_cyc), .QN() );
  SDFFARX1 m6_s10_cyc_o_reg ( .D(n17662), .SI(test_si33), .SE(test_se), .CLK(
        clk_i), .RSTB(n20914), .Q(m6s10_cyc), .QN() );
  SDFFARX1 m6_s9_cyc_o_reg ( .D(n17661), .SI(m6s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20914), .Q(test_so32), .QN() );
  SDFFARX1 m6_s8_cyc_o_reg ( .D(n17660), .SI(m6s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20914), .Q(m6s8_cyc), .QN() );
  SDFFARX1 m6_s7_cyc_o_reg ( .D(n17659), .SI(m6s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20914), .Q(m6s7_cyc), .QN() );
  SDFFARX1 m6_s6_cyc_o_reg ( .D(n17658), .SI(m6s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20913), .Q(m6s6_cyc), .QN() );
  SDFFARX1 m6_s5_cyc_o_reg ( .D(n17657), .SI(m6s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20913), .Q(m6s5_cyc), .QN() );
  SDFFARX1 m6_s4_cyc_o_reg ( .D(n17656), .SI(test_si32), .SE(test_se), .CLK(
        clk_i), .RSTB(n20913), .Q(m6s4_cyc), .QN() );
  SDFFARX1 m6_s3_cyc_o_reg ( .D(n17655), .SI(m6s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20913), .Q(test_so31), .QN() );
  SDFFARX1 m6_s2_cyc_o_reg ( .D(n17654), .SI(m6s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20913), .Q(m6s2_cyc), .QN() );
  SDFFARX1 m6_s1_cyc_o_reg ( .D(n17653), .SI(m6s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20912), .Q(m6s1_cyc), .QN() );
  SDFFARX1 m6_s0_cyc_o_reg ( .D(n17652), .SI(m5s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20912), .Q(m6s0_cyc), .QN() );
  SDFFARX1 m7_s15_cyc_o_reg ( .D(n17651), .SI(m7s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20912), .Q(m7s15_cyc), .QN() );
  SDFFARX1 m7_s14_cyc_o_reg ( .D(n17650), .SI(m7s13_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20912), .Q(m7s14_cyc), .QN() );
  SDFFARX1 m7_s13_cyc_o_reg ( .D(n17649), .SI(m7s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20912), .Q(m7s13_cyc), .QN() );
  SDFFARX1 m7_s12_cyc_o_reg ( .D(n17648), .SI(test_si36), .SE(test_se), .CLK(
        clk_i), .RSTB(n20911), .Q(m7s12_cyc), .QN() );
  SDFFARX1 m7_s11_cyc_o_reg ( .D(n17647), .SI(m7s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20911), .Q(test_so35), .QN() );
  SDFFARX1 m7_s10_cyc_o_reg ( .D(n17646), .SI(m7s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20911), .Q(m7s10_cyc), .QN() );
  SDFFARX1 m7_s9_cyc_o_reg ( .D(n17645), .SI(m7s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20911), .Q(m7s9_cyc), .QN() );
  SDFFARX1 m7_s8_cyc_o_reg ( .D(n17644), .SI(m7s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20911), .Q(m7s8_cyc), .QN() );
  SDFFARX1 m7_s7_cyc_o_reg ( .D(n17643), .SI(m7s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20910), .Q(m7s7_cyc), .QN() );
  SDFFARX1 m7_s6_cyc_o_reg ( .D(n17642), .SI(test_si35), .SE(test_se), .CLK(
        clk_i), .RSTB(n20910), .Q(m7s6_cyc), .QN() );
  SDFFARX1 m7_s5_cyc_o_reg ( .D(n17641), .SI(m7s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20910), .Q(test_so34), .QN() );
  SDFFARX1 m7_s4_cyc_o_reg ( .D(n17640), .SI(m7s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20910), .Q(m7s4_cyc), .QN() );
  SDFFARX1 m7_s3_cyc_o_reg ( .D(n17639), .SI(m7s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20910), .Q(m7s3_cyc), .QN() );
  SDFFARX1 m7_s2_cyc_o_reg ( .D(n17638), .SI(m7s1_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20909), .Q(m7s2_cyc), .QN() );
  SDFFARX1 m7_s1_cyc_o_reg ( .D(n17637), .SI(m7s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20909), .Q(m7s1_cyc), .QN() );
  SDFFARX1 m7_s0_cyc_o_reg ( .D(n17636), .SI(test_si34), .SE(test_se), .CLK(
        clk_i), .RSTB(n20909), .Q(m7s0_cyc), .QN() );
  SDFFX1 s0_m7_cyc_r_reg ( .D(m7s0_cyc), .SI(s0_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so40), .QN() );
  SDFFX1 s0_m6_cyc_r_reg ( .D(m6s0_cyc), .SI(s0_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s0_m6_cyc_r), .QN() );
  SDFFX1 s0_m5_cyc_r_reg ( .D(m5s0_cyc), .SI(s0_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s0_m5_cyc_r), .QN() );
  SDFFX1 s0_m4_cyc_r_reg ( .D(n18321), .SI(s0_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s0_m4_cyc_r), .QN() );
  SDFFX1 s0_m3_cyc_r_reg ( .D(test_so23), .SI(s0_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s0_m3_cyc_r), .QN() );
  SDFFX1 s0_m2_cyc_r_reg ( .D(m2s0_cyc), .SI(test_si40), .SE(test_se), .CLK(
        clk_i), .Q(s0_m2_cyc_r), .QN() );
  SDFFX1 s0_m1_cyc_r_reg ( .D(m1s0_cyc), .SI(s0_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so39), .QN() );
  SDFFX1 s0_m0_cyc_r_reg ( .D(m0s0_cyc), .SI(n21168), .SE(test_se), .CLK(clk_i), .Q(s0_m0_cyc_r), .QN() );
  SDFFX1 s1_m7_cyc_r_reg ( .D(m7s1_cyc), .SI(s1_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s1_m7_cyc_r), .QN() );
  SDFFX1 s1_m6_cyc_r_reg ( .D(m6s1_cyc), .SI(s1_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s1_m6_cyc_r), .QN() );
  SDFFX1 s1_m5_cyc_r_reg ( .D(test_so28), .SI(s1_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s1_m5_cyc_r), .QN() );
  SDFFX1 s1_m4_cyc_r_reg ( .D(n18322), .SI(s1_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s1_m4_cyc_r), .QN() );
  SDFFX1 s1_m3_cyc_r_reg ( .D(m3s1_cyc), .SI(test_si44), .SE(test_se), .CLK(
        clk_i), .Q(s1_m3_cyc_r), .QN() );
  SDFFX1 s1_m2_cyc_r_reg ( .D(m2s1_cyc), .SI(s1_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so43), .QN() );
  SDFFX1 s1_m1_cyc_r_reg ( .D(m1s1_cyc), .SI(s1_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s1_m1_cyc_r), .QN() );
  SDFFX1 s1_m0_cyc_r_reg ( .D(m0s1_cyc), .SI(s0_next), .SE(test_se), .CLK(
        clk_i), .Q(s1_m0_cyc_r), .QN() );
  SDFFX1 s2_m7_cyc_r_reg ( .D(m7s2_cyc), .SI(s2_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s2_m7_cyc_r), .QN() );
  SDFFX1 s2_m6_cyc_r_reg ( .D(m6s2_cyc), .SI(s2_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s2_m6_cyc_r), .QN() );
  SDFFX1 s2_m5_cyc_r_reg ( .D(m5s2_cyc), .SI(s2_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s2_m5_cyc_r), .QN() );
  SDFFX1 s2_m4_cyc_r_reg ( .D(n18325), .SI(test_si48), .SE(test_se), .CLK(
        clk_i), .Q(s2_m4_cyc_r), .QN() );
  SDFFX1 s2_m3_cyc_r_reg ( .D(m3s2_cyc), .SI(s2_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so47), .QN() );
  SDFFX1 s2_m2_cyc_r_reg ( .D(test_so21), .SI(s2_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s2_m2_cyc_r), .QN() );
  SDFFX1 s2_m1_cyc_r_reg ( .D(m1s2_cyc), .SI(s2_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s2_m1_cyc_r), .QN() );
  SDFFX1 s2_m0_cyc_r_reg ( .D(m0s2_cyc), .SI(s1_next), .SE(test_se), .CLK(
        clk_i), .Q(s2_m0_cyc_r), .QN() );
  SDFFX1 s3_m7_cyc_r_reg ( .D(m7s3_cyc), .SI(s3_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s3_m7_cyc_r), .QN() );
  SDFFX1 s3_m6_cyc_r_reg ( .D(test_so31), .SI(s3_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s3_m6_cyc_r), .QN() );
  SDFFX1 s3_m5_cyc_r_reg ( .D(m5s3_cyc), .SI(test_si52), .SE(test_se), .CLK(
        clk_i), .Q(s3_m5_cyc_r), .QN() );
  SDFFX1 s3_m4_cyc_r_reg ( .D(n18326), .SI(s3_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so51), .QN() );
  SDFFX1 s3_m3_cyc_r_reg ( .D(m3s3_cyc), .SI(s3_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s3_m3_cyc_r), .QN() );
  SDFFX1 s3_m2_cyc_r_reg ( .D(m2s3_cyc), .SI(s3_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s3_m2_cyc_r), .QN() );
  SDFFX1 s3_m1_cyc_r_reg ( .D(m1s3_cyc), .SI(s3_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s3_m1_cyc_r), .QN() );
  SDFFX1 s3_m0_cyc_r_reg ( .D(m0s3_cyc), .SI(s2_next), .SE(test_se), .CLK(
        clk_i), .Q(s3_m0_cyc_r), .QN() );
  SDFFX1 s4_m7_cyc_r_reg ( .D(m7s4_cyc), .SI(s4_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s4_m7_cyc_r), .QN() );
  SDFFX1 s4_m6_cyc_r_reg ( .D(m6s4_cyc), .SI(test_si56), .SE(test_se), .CLK(
        clk_i), .Q(s4_m6_cyc_r), .QN() );
  SDFFX1 s4_m5_cyc_r_reg ( .D(m5s4_cyc), .SI(s4_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so55), .QN() );
  SDFFX1 s4_m4_cyc_r_reg ( .D(n18329), .SI(s4_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s4_m4_cyc_r), .QN() );
  SDFFX1 s4_m3_cyc_r_reg ( .D(m3s4_cyc), .SI(s4_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s4_m3_cyc_r), .QN() );
  SDFFX1 s4_m2_cyc_r_reg ( .D(m2s4_cyc), .SI(s4_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s4_m2_cyc_r), .QN() );
  SDFFX1 s4_m1_cyc_r_reg ( .D(test_so19), .SI(s4_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s4_m1_cyc_r), .QN() );
  SDFFX1 s4_m0_cyc_r_reg ( .D(m0s4_cyc), .SI(test_si55), .SE(test_se), .CLK(
        clk_i), .Q(s4_m0_cyc_r), .QN() );
  SDFFX1 s5_m7_cyc_r_reg ( .D(test_so34), .SI(test_si60), .SE(test_se), .CLK(
        clk_i), .Q(s5_m7_cyc_r), .QN() );
  SDFFX1 s5_m6_cyc_r_reg ( .D(m6s5_cyc), .SI(s5_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so59), .QN() );
  SDFFX1 s5_m5_cyc_r_reg ( .D(m5s5_cyc), .SI(s5_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s5_m5_cyc_r), .QN() );
  SDFFX1 s5_m4_cyc_r_reg ( .D(n18330), .SI(s5_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s5_m4_cyc_r), .QN() );
  SDFFX1 s5_m3_cyc_r_reg ( .D(m3s5_cyc), .SI(s5_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s5_m3_cyc_r), .QN() );
  SDFFX1 s5_m2_cyc_r_reg ( .D(m2s5_cyc), .SI(s5_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s5_m2_cyc_r), .QN() );
  SDFFX1 s5_m1_cyc_r_reg ( .D(m1s5_cyc), .SI(test_si59), .SE(test_se), .CLK(
        clk_i), .Q(s5_m1_cyc_r), .QN() );
  SDFFX1 s5_m0_cyc_r_reg ( .D(m0s5_cyc), .SI(s4_next), .SE(test_se), .CLK(
        clk_i), .Q(test_so58), .QN() );
  SDFFX1 s6_m7_cyc_r_reg ( .D(m7s6_cyc), .SI(s6_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so63), .QN() );
  SDFFX1 s6_m6_cyc_r_reg ( .D(m6s6_cyc), .SI(s6_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s6_m6_cyc_r), .QN() );
  SDFFX1 s6_m5_cyc_r_reg ( .D(m5s6_cyc), .SI(s6_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s6_m5_cyc_r), .QN() );
  SDFFX1 s6_m4_cyc_r_reg ( .D(n18332), .SI(s6_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s6_m4_cyc_r), .QN() );
  SDFFX1 s6_m3_cyc_r_reg ( .D(m3s6_cyc), .SI(s6_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s6_m3_cyc_r), .QN() );
  SDFFX1 s6_m2_cyc_r_reg ( .D(m2s6_cyc), .SI(test_si63), .SE(test_se), .CLK(
        clk_i), .Q(s6_m2_cyc_r), .QN() );
  SDFFX1 s6_m1_cyc_r_reg ( .D(m1s6_cyc), .SI(s6_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so62), .QN() );
  SDFFX1 s6_m0_cyc_r_reg ( .D(test_so17), .SI(s5_next), .SE(test_se), .CLK(
        clk_i), .Q(s6_m0_cyc_r), .QN() );
  SDFFX1 s7_m7_cyc_r_reg ( .D(m7s7_cyc), .SI(s7_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s7_m7_cyc_r), .QN() );
  SDFFX1 s7_m6_cyc_r_reg ( .D(m6s7_cyc), .SI(s7_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s7_m6_cyc_r), .QN() );
  SDFFX1 s7_m5_cyc_r_reg ( .D(test_so29), .SI(s7_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s7_m5_cyc_r), .QN() );
  SDFFX1 s7_m4_cyc_r_reg ( .D(n18333), .SI(s7_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s7_m4_cyc_r), .QN() );
  SDFFX1 s7_m3_cyc_r_reg ( .D(test_so24), .SI(test_si67), .SE(test_se), .CLK(
        clk_i), .Q(s7_m3_cyc_r), .QN() );
  SDFFX1 s7_m2_cyc_r_reg ( .D(m2s7_cyc), .SI(s7_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so66), .QN() );
  SDFFX1 s7_m1_cyc_r_reg ( .D(m1s7_cyc), .SI(s7_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s7_m1_cyc_r), .QN() );
  SDFFX1 s7_m0_cyc_r_reg ( .D(m0s7_cyc), .SI(s6_next), .SE(test_se), .CLK(
        clk_i), .Q(s7_m0_cyc_r), .QN() );
  SDFFX1 s8_m7_cyc_r_reg ( .D(m7s8_cyc), .SI(s8_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s8_m7_cyc_r), .QN() );
  SDFFX1 s8_m6_cyc_r_reg ( .D(m6s8_cyc), .SI(s8_m5_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s8_m6_cyc_r), .QN() );
  SDFFX1 s8_m5_cyc_r_reg ( .D(m5s8_cyc), .SI(s8_m4_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s8_m5_cyc_r), .QN() );
  SDFFX1 s8_m4_cyc_r_reg ( .D(n18319), .SI(test_si71), .SE(test_se), .CLK(
        clk_i), .Q(s8_m4_cyc_r), .QN() );
  SDFFX1 s8_m3_cyc_r_reg ( .D(m3s8_cyc), .SI(s8_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so70), .QN() );
  SDFFX1 s8_m2_cyc_r_reg ( .D(m2s8_cyc), .SI(s8_m1_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s8_m2_cyc_r), .QN() );
  SDFFX1 s8_m1_cyc_r_reg ( .D(m1s8_cyc), .SI(s8_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s8_m1_cyc_r), .QN() );
  SDFFX1 s8_m0_cyc_r_reg ( .D(m0s8_cyc), .SI(s7_next), .SE(test_se), .CLK(
        clk_i), .Q(s8_m0_cyc_r), .QN() );
  SDFFX1 s9_m7_cyc_r_reg ( .D(m7s9_cyc), .SI(s9_m6_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s9_m7_cyc_r), .QN() );
  SDFFX1 s9_m6_cyc_r_reg ( .D(test_so32), .SI(s9_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s9_m6_cyc_r), .QN() );
  SDFFX1 s9_m5_cyc_r_reg ( .D(m5s9_cyc), .SI(test_si75), .SE(test_se), .CLK(
        clk_i), .Q(s9_m5_cyc_r), .QN() );
  SDFFX1 s9_m4_cyc_r_reg ( .D(n18320), .SI(s9_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(test_so74), .QN() );
  SDFFX1 s9_m3_cyc_r_reg ( .D(m3s9_cyc), .SI(s9_m2_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s9_m3_cyc_r), .QN() );
  SDFFX1 s9_m2_cyc_r_reg ( .D(test_so22), .SI(s9_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s9_m2_cyc_r), .QN() );
  SDFFX1 s9_m1_cyc_r_reg ( .D(m1s9_cyc), .SI(s9_m0_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s9_m1_cyc_r), .QN() );
  SDFFX1 s9_m0_cyc_r_reg ( .D(m0s9_cyc), .SI(s8_next), .SE(test_se), .CLK(
        clk_i), .Q(s9_m0_cyc_r), .QN() );
  SDFFX1 s10_m7_cyc_r_reg ( .D(m7s10_cyc), .SI(s10_m6_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s10_m7_cyc_r), .QN() );
  SDFFX1 s10_m6_cyc_r_reg ( .D(m6s10_cyc), .SI(test_si79), .SE(test_se), .CLK(
        clk_i), .Q(s10_m6_cyc_r), .QN() );
  SDFFX1 s10_m5_cyc_r_reg ( .D(m5s10_cyc), .SI(s10_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so78), .QN() );
  SDFFX1 s10_m4_cyc_r_reg ( .D(n18323), .SI(s10_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s10_m4_cyc_r), .QN() );
  SDFFX1 s10_m3_cyc_r_reg ( .D(m3s10_cyc), .SI(s10_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s10_m3_cyc_r), .QN() );
  SDFFX1 s10_m2_cyc_r_reg ( .D(m2s10_cyc), .SI(s10_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s10_m2_cyc_r), .QN() );
  SDFFX1 s10_m1_cyc_r_reg ( .D(m1s10_cyc), .SI(s10_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s10_m1_cyc_r), .QN() );
  SDFFX1 s10_m0_cyc_r_reg ( .D(m0s10_cyc), .SI(test_si78), .SE(test_se), .CLK(
        clk_i), .Q(s10_m0_cyc_r), .QN() );
  SDFFX1 s11_m7_cyc_r_reg ( .D(test_so35), .SI(test_si83), .SE(test_se), .CLK(
        clk_i), .Q(s11_m7_cyc_r), .QN() );
  SDFFX1 s11_m6_cyc_r_reg ( .D(m6s11_cyc), .SI(s11_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so82), .QN() );
  SDFFX1 s11_m5_cyc_r_reg ( .D(m5s11_cyc), .SI(s11_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s11_m5_cyc_r), .QN() );
  SDFFX1 s11_m4_cyc_r_reg ( .D(n18324), .SI(s11_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s11_m4_cyc_r), .QN() );
  SDFFX1 s11_m3_cyc_r_reg ( .D(m3s11_cyc), .SI(s11_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s11_m3_cyc_r), .QN() );
  SDFFX1 s11_m2_cyc_r_reg ( .D(m2s11_cyc), .SI(s11_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s11_m2_cyc_r), .QN() );
  SDFFX1 s11_m1_cyc_r_reg ( .D(test_so20), .SI(test_si82), .SE(test_se), .CLK(
        clk_i), .Q(s11_m1_cyc_r), .QN() );
  SDFFX1 s11_m0_cyc_r_reg ( .D(m0s11_cyc), .SI(s10_next), .SE(test_se), .CLK(
        clk_i), .Q(test_so81), .QN() );
  SDFFX1 s12_m7_cyc_r_reg ( .D(m7s12_cyc), .SI(s12_m6_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so86), .QN() );
  SDFFX1 s12_m6_cyc_r_reg ( .D(m6s12_cyc), .SI(s12_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s12_m6_cyc_r), .QN() );
  SDFFX1 s12_m5_cyc_r_reg ( .D(m5s12_cyc), .SI(s12_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s12_m5_cyc_r), .QN() );
  SDFFX1 s12_m4_cyc_r_reg ( .D(n18327), .SI(s12_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s12_m4_cyc_r), .QN() );
  SDFFX1 s12_m3_cyc_r_reg ( .D(m3s12_cyc), .SI(s12_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s12_m3_cyc_r), .QN() );
  SDFFX1 s12_m2_cyc_r_reg ( .D(m2s12_cyc), .SI(test_si86), .SE(test_se), .CLK(
        clk_i), .Q(s12_m2_cyc_r), .QN() );
  SDFFX1 s12_m1_cyc_r_reg ( .D(m1s12_cyc), .SI(s12_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so85), .QN() );
  SDFFX1 s12_m0_cyc_r_reg ( .D(m0s12_cyc), .SI(s11_next), .SE(test_se), .CLK(
        clk_i), .Q(s12_m0_cyc_r), .QN() );
  SDFFX1 s13_m7_cyc_r_reg ( .D(m7s13_cyc), .SI(s13_m6_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s13_m7_cyc_r), .QN() );
  SDFFX1 s13_m6_cyc_r_reg ( .D(m6s13_cyc), .SI(s13_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s13_m6_cyc_r), .QN() );
  SDFFX1 s13_m5_cyc_r_reg ( .D(test_so30), .SI(s13_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s13_m5_cyc_r), .QN() );
  SDFFX1 s13_m4_cyc_r_reg ( .D(n18328), .SI(s13_m3_cyc_r), .SE(test_se), .CLK(
        clk_i), .Q(s13_m4_cyc_r), .QN() );
  SDFFX1 s13_m3_cyc_r_reg ( .D(m3s13_cyc), .SI(test_si90), .SE(test_se), .CLK(
        clk_i), .Q(s13_m3_cyc_r), .QN() );
  SDFFX1 s13_m2_cyc_r_reg ( .D(m2s13_cyc), .SI(s13_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so89), .QN() );
  SDFFX1 s13_m1_cyc_r_reg ( .D(m1s13_cyc), .SI(s13_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s13_m1_cyc_r), .QN() );
  SDFFX1 s13_m0_cyc_r_reg ( .D(test_so18), .SI(s12_next), .SE(test_se), .CLK(
        clk_i), .Q(s13_m0_cyc_r), .QN() );
  SDFFX1 s14_m7_cyc_r_reg ( .D(m7s14_cyc), .SI(s14_m6_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s14_m7_cyc_r), .QN() );
  SDFFX1 s14_m6_cyc_r_reg ( .D(m6s14_cyc), .SI(s14_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s14_m6_cyc_r), .QN() );
  SDFFX1 s14_m5_cyc_r_reg ( .D(m5s14_cyc), .SI(s14_m4_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s14_m5_cyc_r), .QN() );
  SDFFX1 s14_m4_cyc_r_reg ( .D(n18331), .SI(test_si94), .SE(test_se), .CLK(
        clk_i), .Q(s14_m4_cyc_r), .QN() );
  SDFFX1 s14_m3_cyc_r_reg ( .D(test_so25), .SI(s14_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so93), .QN() );
  SDFFX1 s14_m2_cyc_r_reg ( .D(m2s14_cyc), .SI(s14_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s14_m2_cyc_r), .QN() );
  SDFFX1 s14_m1_cyc_r_reg ( .D(m1s14_cyc), .SI(s14_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s14_m1_cyc_r), .QN() );
  SDFFX1 s14_m0_cyc_r_reg ( .D(m0s14_cyc), .SI(s13_next), .SE(test_se), .CLK(
        clk_i), .Q(s14_m0_cyc_r), .QN() );
  SDFFX1 s15_m7_cyc_r_reg ( .D(m7s15_cyc), .SI(s15_m6_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s15_m7_cyc_r), .QN() );
  SDFFX1 s15_m6_cyc_r_reg ( .D(test_so33), .SI(s15_m5_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s15_m6_cyc_r), .QN() );
  SDFFX1 s15_m5_cyc_r_reg ( .D(m5s15_cyc), .SI(test_si98), .SE(test_se), .CLK(
        clk_i), .Q(s15_m5_cyc_r), .QN() );
  SDFFX1 s15_m4_cyc_r_reg ( .D(m4s15_cyc), .SI(s15_m3_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(test_so97), .QN() );
  SDFFX1 s15_m3_cyc_r_reg ( .D(m3s15_cyc), .SI(s15_m2_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s15_m3_cyc_r), .QN() );
  SDFFX1 s15_m2_cyc_r_reg ( .D(m2s15_cyc), .SI(s15_m1_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s15_m2_cyc_r), .QN() );
  SDFFX1 s15_m1_cyc_r_reg ( .D(m1s15_cyc), .SI(s15_m0_cyc_r), .SE(test_se), 
        .CLK(clk_i), .Q(s15_m1_cyc_r), .QN() );
  SDFFX1 s15_m0_cyc_r_reg ( .D(m0s15_cyc), .SI(s14_next), .SE(test_se), .CLK(
        clk_i), .Q(s15_m0_cyc_r), .QN() );
  SDFFX1 rf_rf_we_reg ( .D(rf_N18), .SI(rf_rf_dout_15_), .SE(test_se), .CLK(
        clk_i), .Q(n21168), .QN(n4502) );
  SDFFX1 s15_msel_pri_out_reg_1_ ( .D(n17634), .SI(s15_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s15_msel_pri_out_1_), .QN(n4213) );
  SDFFX1 s15_msel_pri_out_reg_0_ ( .D(n17633), .SI(s15_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s15_msel_pri_out_0_), .QN(n4212) );
  SDFFARX1 s15_msel_arb2_state_reg_2_ ( .D(n17612), .SI(s15_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20909), .Q(test_so99), .QN(n4237) );
  SDFFX1 s15_next_reg ( .D(n17764), .SI(s15_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(test_so100), .QN() );
  SDFFARX1 s15_msel_arb0_state_reg_2_ ( .D(n17609), .SI(s15_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20909), .Q(test_so98), .QN(n4221) );
  SDFFARX1 s15_msel_arb0_state_reg_0_ ( .D(n17611), .SI(s15_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20908), .Q(s15_msel_gnt_p0_0_), .QN(
        n4219) );
  SDFFARX1 s15_msel_arb0_state_reg_1_ ( .D(n17610), .SI(s15_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20908), .Q(s15_msel_gnt_p0_1_), .QN(
        n4220) );
  SDFFARX1 s15_msel_arb2_state_reg_0_ ( .D(n17614), .SI(s15_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20908), .Q(s15_msel_gnt_p2_0_), .QN(
        n4235) );
  SDFFARX1 s15_msel_arb2_state_reg_1_ ( .D(n17613), .SI(s15_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20908), .Q(s15_msel_gnt_p2_1_), .QN(
        n4236) );
  SDFFARX1 s15_msel_arb3_state_reg_0_ ( .D(n17617), .SI(test_si100), .SE(
        test_se), .CLK(clk_i), .RSTB(n20908), .Q(s15_msel_gnt_p3[0]), .QN(
        n4243) );
  SDFFARX1 s15_msel_arb3_state_reg_2_ ( .D(n17615), .SI(s15_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20907), .Q(s15_msel_gnt_p3[2]), .QN(
        n4245) );
  SDFFARX1 s15_msel_arb3_state_reg_1_ ( .D(n17616), .SI(s15_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20907), .Q(s15_msel_gnt_p3[1]), .QN(
        n4244) );
  SDFFARX1 s15_msel_arb1_state_reg_2_ ( .D(n17606), .SI(s15_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20907), .Q(s15_msel_gnt_p1[2]), .QN(
        n4229) );
  SDFFARX1 s15_msel_arb1_state_reg_0_ ( .D(n17608), .SI(test_si99), .SE(
        test_se), .CLK(clk_i), .RSTB(n20907), .Q(s15_msel_gnt_p1[0]), .QN(
        n4227) );
  SDFFARX1 s15_msel_arb1_state_reg_1_ ( .D(n17607), .SI(s15_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20907), .Q(s15_msel_gnt_p1[1]), .QN(
        n4228) );
  SDFFARX1 s8_msel_arb2_state_reg_2_ ( .D(n17158), .SI(test_si73), .SE(test_se), .CLK(clk_i), .RSTB(n20906), .Q(s8_msel_gnt_p2_2_), .QN(n3922) );
  SDFFARX1 s8_msel_arb2_state_reg_0_ ( .D(n17160), .SI(s8_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20906), .Q(s8_msel_gnt_p2_0_), .QN(
        n3920) );
  SDFFARX1 s8_msel_arb2_state_reg_1_ ( .D(n17159), .SI(s8_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20906), .Q(test_so72), .QN(n3921) );
  SDFFARX1 s8_msel_arb0_state_reg_2_ ( .D(n17161), .SI(test_si72), .SE(test_se), .CLK(clk_i), .RSTB(n20906), .Q(s8_msel_gnt_p0_2_), .QN(n3906) );
  SDFFARX1 s8_msel_arb0_state_reg_0_ ( .D(n17163), .SI(s8_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20906), .Q(s8_msel_gnt_p0_0_), .QN(n3904) );
  SDFFARX1 s8_msel_arb0_state_reg_1_ ( .D(n17162), .SI(s8_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20905), .Q(test_so71), .QN(n3905) );
  SDFFARX1 s8_msel_arb1_state_reg_2_ ( .D(n17164), .SI(s8_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20905), .Q(s8_msel_gnt_p1[2]), .QN(
        n3914) );
  SDFFARX1 s8_msel_arb1_state_reg_0_ ( .D(n17166), .SI(s8_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20905), .Q(s8_msel_gnt_p1[0]), .QN(
        n3912) );
  SDFFARX1 s8_msel_arb1_state_reg_1_ ( .D(n17165), .SI(s8_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20905), .Q(s8_msel_gnt_p1[1]), .QN(
        n3913) );
  SDFFARX1 s8_msel_arb3_state_reg_0_ ( .D(n17169), .SI(s8_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20905), .Q(s8_msel_gnt_p3[0]), .QN(
        n3928) );
  SDFFARX1 s8_msel_arb3_state_reg_2_ ( .D(n17167), .SI(s8_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20904), .Q(s8_msel_gnt_p3[2]), .QN(
        n3930) );
  SDFFARX1 s8_msel_arb3_state_reg_1_ ( .D(n17168), .SI(s8_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20904), .Q(s8_msel_gnt_p3[1]), .QN(
        n3929) );
  SDFFX1 s8_next_reg ( .D(n17771), .SI(test_si74), .SE(test_se), .CLK(clk_i), 
        .Q(s8_next), .QN() );
  SDFFX1 s8_msel_pri_out_reg_0_ ( .D(n17156), .SI(s8_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s8_msel_pri_out_0_), .QN(n3897) );
  SDFFX1 s8_msel_pri_out_reg_1_ ( .D(n17157), .SI(s8_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(test_so73), .QN(n3898) );
  SDFFARX1 s9_msel_arb2_state_reg_2_ ( .D(n17188), .SI(s9_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20904), .Q(test_so76), .QN(n3967) );
  SDFFARX1 s9_msel_arb2_state_reg_0_ ( .D(n17190), .SI(s9_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20904), .Q(s9_msel_gnt_p2_0_), .QN(
        n3965) );
  SDFFARX1 s9_msel_arb2_state_reg_1_ ( .D(n17189), .SI(s9_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20904), .Q(s9_msel_gnt_p2_1_), .QN(
        n3966) );
  SDFFARX1 s9_msel_arb0_state_reg_2_ ( .D(n17191), .SI(s9_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20903), .Q(test_so75), .QN(n3951) );
  SDFFARX1 s9_msel_arb0_state_reg_0_ ( .D(n17193), .SI(s9_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20903), .Q(s9_msel_gnt_p0_0_), .QN(n3949) );
  SDFFARX1 s9_msel_arb0_state_reg_1_ ( .D(n17192), .SI(s9_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20903), .Q(s9_msel_gnt_p0_1_), .QN(
        n3950) );
  SDFFARX1 s9_msel_arb1_state_reg_2_ ( .D(n17194), .SI(s9_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20903), .Q(s9_msel_gnt_p1[2]), .QN(
        n3959) );
  SDFFARX1 s9_msel_arb1_state_reg_0_ ( .D(n17196), .SI(test_si76), .SE(test_se), .CLK(clk_i), .RSTB(n20903), .Q(s9_msel_gnt_p1[0]), .QN(n3957) );
  SDFFARX1 s9_msel_arb1_state_reg_1_ ( .D(n17195), .SI(s9_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20902), .Q(s9_msel_gnt_p1[1]), .QN(
        n3958) );
  SDFFARX1 s9_msel_arb3_state_reg_0_ ( .D(n17199), .SI(test_si77), .SE(test_se), .CLK(clk_i), .RSTB(n20902), .Q(s9_msel_gnt_p3[0]), .QN(n3973) );
  SDFFARX1 s9_msel_arb3_state_reg_2_ ( .D(n17197), .SI(s9_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20902), .Q(s9_msel_gnt_p3[2]), .QN(
        n3975) );
  SDFFARX1 s9_msel_arb3_state_reg_1_ ( .D(n17198), .SI(s9_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20902), .Q(s9_msel_gnt_p3[1]), .QN(
        n3974) );
  SDFFX1 s9_next_reg ( .D(n17770), .SI(s9_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(test_so77), .QN() );
  SDFFX1 s9_msel_pri_out_reg_0_ ( .D(n17186), .SI(s9_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s9_msel_pri_out_0_), .QN(n3942) );
  SDFFX1 s9_msel_pri_out_reg_1_ ( .D(n17187), .SI(s9_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s9_msel_pri_out_1_), .QN(n3943) );
  SDFFARX1 s0_msel_arb2_state_reg_2_ ( .D(n17368), .SI(s0_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20902), .Q(s0_msel_gnt_p2[2]), .QN(
        n3562) );
  SDFFARX1 s0_msel_arb2_state_reg_0_ ( .D(n17370), .SI(test_si42), .SE(test_se), .CLK(clk_i), .RSTB(n20901), .Q(s0_msel_gnt_p2[0]), .QN(n3560) );
  SDFFARX1 s0_msel_arb2_state_reg_1_ ( .D(n17369), .SI(s0_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20901), .Q(s0_msel_gnt_p2[1]), .QN(
        n3561) );
  SDFFARX1 s0_msel_arb0_state_reg_2_ ( .D(n17371), .SI(s0_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20901), .Q(s0_msel_gnt_p0[2]), .QN(
        n3546) );
  SDFFARX1 s0_msel_arb0_state_reg_0_ ( .D(n17373), .SI(test_si41), .SE(test_se), .CLK(clk_i), .RSTB(n20901), .Q(s0_msel_gnt_p0[0]), .QN(n3544) );
  SDFFARX1 s0_msel_arb0_state_reg_1_ ( .D(n17372), .SI(s0_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20901), .Q(s0_msel_gnt_p0[1]), .QN(
        n3545) );
  SDFFARX1 s0_msel_arb1_state_reg_2_ ( .D(n17374), .SI(s0_msel_gnt_p1_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20900), .Q(test_so41), .QN(n3554) );
  SDFFARX1 s0_msel_arb1_state_reg_0_ ( .D(n17376), .SI(s0_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20900), .Q(s0_msel_gnt_p1_0_), .QN(
        n3552) );
  SDFFARX1 s0_msel_arb1_state_reg_1_ ( .D(n17375), .SI(s0_msel_gnt_p1_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20900), .Q(s0_msel_gnt_p1_1_), .QN(
        n3553) );
  SDFFARX1 s0_msel_arb3_state_reg_0_ ( .D(n17379), .SI(s0_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20900), .Q(s0_msel_gnt_p3_0_), .QN(
        n3568) );
  SDFFARX1 s0_msel_arb3_state_reg_2_ ( .D(n17377), .SI(s0_msel_gnt_p3_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20900), .Q(test_so42), .QN(n3570) );
  SDFFARX1 s0_msel_arb3_state_reg_1_ ( .D(n17378), .SI(s0_msel_gnt_p3_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20899), .Q(s0_msel_gnt_p3_1_), .QN(
        n3569) );
  SDFFX1 s0_next_reg ( .D(n17779), .SI(s0_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s0_next), .QN() );
  SDFFX1 s0_msel_pri_out_reg_0_ ( .D(n17366), .SI(test_si43), .SE(test_se), 
        .CLK(clk_i), .Q(s0_msel_pri_out_0_), .QN(n3537) );
  SDFFX1 s0_msel_pri_out_reg_1_ ( .D(n17367), .SI(s0_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s0_msel_pri_out_1_), .QN(n3538) );
  SDFFARX1 s1_msel_arb2_state_reg_2_ ( .D(n17398), .SI(s1_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20899), .Q(s1_msel_gnt_p2_2_), .QN(
        n3607) );
  SDFFARX1 s1_msel_arb2_state_reg_0_ ( .D(n17400), .SI(s1_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20899), .Q(test_so45), .QN(n3605) );
  SDFFARX1 s1_msel_arb2_state_reg_1_ ( .D(n17399), .SI(test_si46), .SE(test_se), .CLK(clk_i), .RSTB(n20899), .Q(s1_msel_gnt_p2_1_), .QN(n3606) );
  SDFFARX1 s1_msel_arb0_state_reg_2_ ( .D(n17401), .SI(s1_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20899), .Q(s1_msel_gnt_p0_2_), .QN(
        n3591) );
  SDFFARX1 s1_msel_arb0_state_reg_0_ ( .D(n17403), .SI(s1_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20898), .Q(test_so44), .QN(n3589) );
  SDFFARX1 s1_msel_arb0_state_reg_1_ ( .D(n17402), .SI(test_si45), .SE(test_se), .CLK(clk_i), .RSTB(n20898), .Q(s1_msel_gnt_p0_1_), .QN(n3590) );
  SDFFARX1 s1_msel_arb1_state_reg_2_ ( .D(n17404), .SI(s1_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20898), .Q(s1_msel_gnt_p1[2]), .QN(
        n3599) );
  SDFFARX1 s1_msel_arb1_state_reg_0_ ( .D(n17406), .SI(s1_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20898), .Q(s1_msel_gnt_p1[0]), .QN(
        n3597) );
  SDFFARX1 s1_msel_arb1_state_reg_1_ ( .D(n17405), .SI(s1_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20898), .Q(s1_msel_gnt_p1[1]), .QN(
        n3598) );
  SDFFARX1 s1_msel_arb3_state_reg_0_ ( .D(n17409), .SI(s1_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20897), .Q(s1_msel_gnt_p3[0]), .QN(
        n3613) );
  SDFFARX1 s1_msel_arb3_state_reg_2_ ( .D(n17407), .SI(s1_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20897), .Q(s1_msel_gnt_p3[2]), .QN(
        n3615) );
  SDFFARX1 s1_msel_arb3_state_reg_1_ ( .D(n17408), .SI(s1_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20897), .Q(s1_msel_gnt_p3[1]), .QN(
        n3614) );
  SDFFX1 s1_next_reg ( .D(n17778), .SI(s1_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s1_next), .QN() );
  SDFFX1 s1_msel_pri_out_reg_0_ ( .D(n17396), .SI(s1_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(test_so46), .QN(n3582) );
  SDFFX1 s1_msel_pri_out_reg_1_ ( .D(n17397), .SI(test_si47), .SE(test_se), 
        .CLK(clk_i), .Q(s1_msel_pri_out_1_), .QN(n3583) );
  SDFFARX1 s10_msel_arb2_state_reg_2_ ( .D(n17218), .SI(s10_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20897), .Q(s10_msel_gnt_p2[2]), .QN(
        n4012) );
  SDFFARX1 s10_msel_arb2_state_reg_0_ ( .D(n17220), .SI(s10_msel_gnt_p1_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20897), .Q(s10_msel_gnt_p2[0]), .QN(
        n4010) );
  SDFFARX1 s10_msel_arb2_state_reg_1_ ( .D(n17219), .SI(s10_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20896), .Q(s10_msel_gnt_p2[1]), .QN(
        n4011) );
  SDFFARX1 s10_msel_arb0_state_reg_2_ ( .D(n17221), .SI(s10_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20896), .Q(s10_msel_gnt_p0[2]), .QN(
        n3996) );
  SDFFARX1 s10_msel_arb0_state_reg_0_ ( .D(n17223), .SI(s10_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20896), .Q(s10_msel_gnt_p0[0]), .QN(
        n3994) );
  SDFFARX1 s10_msel_arb0_state_reg_1_ ( .D(n17222), .SI(s10_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20896), .Q(s10_msel_gnt_p0[1]), .QN(
        n3995) );
  SDFFARX1 s10_msel_arb1_state_reg_2_ ( .D(n17224), .SI(s10_msel_gnt_p1_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20896), .Q(s10_msel_gnt_p1_2_), .QN(
        n4004) );
  SDFFARX1 s10_msel_arb1_state_reg_0_ ( .D(n17226), .SI(s10_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20895), .Q(test_so79), .QN(n4002) );
  SDFFARX1 s10_msel_arb1_state_reg_1_ ( .D(n17225), .SI(test_si80), .SE(
        test_se), .CLK(clk_i), .RSTB(n20895), .Q(s10_msel_gnt_p1_1_), .QN(
        n4003) );
  SDFFARX1 s10_msel_arb3_state_reg_0_ ( .D(n17229), .SI(s10_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20895), .Q(test_so80), .QN(n4018) );
  SDFFARX1 s10_msel_arb3_state_reg_2_ ( .D(n17227), .SI(s10_msel_gnt_p3_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20895), .Q(s10_msel_gnt_p3_2_), .QN(
        n4020) );
  SDFFARX1 s10_msel_arb3_state_reg_1_ ( .D(n17228), .SI(test_si81), .SE(
        test_se), .CLK(clk_i), .RSTB(n20895), .Q(s10_msel_gnt_p3_1_), .QN(
        n4019) );
  SDFFX1 s10_next_reg ( .D(n17769), .SI(s10_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s10_next), .QN() );
  SDFFX1 s10_msel_pri_out_reg_0_ ( .D(n17216), .SI(s10_msel_gnt_p3_2_), .SE(
        test_se), .CLK(clk_i), .Q(s10_msel_pri_out_0_), .QN(n3987) );
  SDFFX1 s10_msel_pri_out_reg_1_ ( .D(n17217), .SI(s10_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s10_msel_pri_out_1_), .QN(n3988) );
  SDFFARX1 s11_msel_arb2_state_reg_2_ ( .D(n17248), .SI(s11_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20894), .Q(s11_msel_gnt_p2[2]), .QN(
        n4057) );
  SDFFARX1 s11_msel_arb2_state_reg_0_ ( .D(n17250), .SI(s11_msel_gnt_p1_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20894), .Q(s11_msel_gnt_p2[0]), .QN(
        n4055) );
  SDFFARX1 s11_msel_arb2_state_reg_1_ ( .D(n17249), .SI(s11_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20894), .Q(s11_msel_gnt_p2[1]), .QN(
        n4056) );
  SDFFARX1 s11_msel_arb0_state_reg_2_ ( .D(n17251), .SI(s11_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20894), .Q(s11_msel_gnt_p0[2]), .QN(
        n4041) );
  SDFFARX1 s11_msel_arb0_state_reg_0_ ( .D(n17253), .SI(s11_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20894), .Q(s11_msel_gnt_p0[0]), .QN(
        n4039) );
  SDFFARX1 s11_msel_arb0_state_reg_1_ ( .D(n17252), .SI(s11_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20893), .Q(s11_msel_gnt_p0[1]), .QN(
        n4040) );
  SDFFARX1 s11_msel_arb1_state_reg_2_ ( .D(n17254), .SI(test_si84), .SE(
        test_se), .CLK(clk_i), .RSTB(n20893), .Q(s11_msel_gnt_p1_2_), .QN(
        n4049) );
  SDFFARX1 s11_msel_arb1_state_reg_0_ ( .D(n17256), .SI(s11_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20893), .Q(s11_msel_gnt_p1_0_), .QN(
        n4047) );
  SDFFARX1 s11_msel_arb1_state_reg_1_ ( .D(n17255), .SI(s11_msel_gnt_p1_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20893), .Q(test_so83), .QN(n4048) );
  SDFFARX1 s11_msel_arb3_state_reg_0_ ( .D(n17259), .SI(s11_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20893), .Q(s11_msel_gnt_p3_0_), .QN(
        n4063) );
  SDFFARX1 s11_msel_arb3_state_reg_2_ ( .D(n17257), .SI(test_si85), .SE(
        test_se), .CLK(clk_i), .RSTB(n20892), .Q(s11_msel_gnt_p3_2_), .QN(
        n4065) );
  SDFFARX1 s11_msel_arb3_state_reg_1_ ( .D(n17258), .SI(s11_msel_gnt_p3_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20892), .Q(test_so84), .QN(n4064) );
  SDFFX1 s11_next_reg ( .D(n17768), .SI(s11_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s11_next), .QN() );
  SDFFX1 s11_msel_pri_out_reg_0_ ( .D(n17246), .SI(s11_msel_gnt_p3_2_), .SE(
        test_se), .CLK(clk_i), .Q(s11_msel_pri_out_0_), .QN(n4032) );
  SDFFX1 s11_msel_pri_out_reg_1_ ( .D(n17247), .SI(s11_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s11_msel_pri_out_1_), .QN(n4033) );
  SDFFARX1 s2_msel_arb2_state_reg_2_ ( .D(n17428), .SI(test_si50), .SE(test_se), .CLK(clk_i), .RSTB(n20892), .Q(s2_msel_gnt_p2_2_), .QN(n3652) );
  SDFFARX1 s2_msel_arb2_state_reg_0_ ( .D(n17430), .SI(s2_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20892), .Q(s2_msel_gnt_p2_0_), .QN(
        n3650) );
  SDFFARX1 s2_msel_arb2_state_reg_1_ ( .D(n17429), .SI(s2_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20892), .Q(test_so49), .QN(n3651) );
  SDFFARX1 s2_msel_arb0_state_reg_2_ ( .D(n17431), .SI(test_si49), .SE(test_se), .CLK(clk_i), .RSTB(n20891), .Q(s2_msel_gnt_p0_2_), .QN(n3636) );
  SDFFARX1 s2_msel_arb0_state_reg_0_ ( .D(n17433), .SI(s2_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20891), .Q(s2_msel_gnt_p0_0_), .QN(n3634) );
  SDFFARX1 s2_msel_arb0_state_reg_1_ ( .D(n17432), .SI(s2_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20891), .Q(test_so48), .QN(n3635) );
  SDFFARX1 s2_msel_arb1_state_reg_2_ ( .D(n17434), .SI(s2_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20891), .Q(s2_msel_gnt_p1[2]), .QN(
        n3644) );
  SDFFARX1 s2_msel_arb1_state_reg_0_ ( .D(n17436), .SI(s2_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20891), .Q(s2_msel_gnt_p1[0]), .QN(
        n3642) );
  SDFFARX1 s2_msel_arb1_state_reg_1_ ( .D(n17435), .SI(s2_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20890), .Q(s2_msel_gnt_p1[1]), .QN(
        n3643) );
  SDFFARX1 s2_msel_arb3_state_reg_0_ ( .D(n17439), .SI(s2_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20890), .Q(s2_msel_gnt_p3[0]), .QN(
        n3658) );
  SDFFARX1 s2_msel_arb3_state_reg_2_ ( .D(n17437), .SI(s2_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20890), .Q(s2_msel_gnt_p3[2]), .QN(
        n3660) );
  SDFFARX1 s2_msel_arb3_state_reg_1_ ( .D(n17438), .SI(s2_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20890), .Q(s2_msel_gnt_p3[1]), .QN(
        n3659) );
  SDFFX1 s2_next_reg ( .D(n17777), .SI(test_si51), .SE(test_se), .CLK(clk_i), 
        .Q(s2_next), .QN() );
  SDFFX1 s2_msel_pri_out_reg_0_ ( .D(n17426), .SI(s2_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s2_msel_pri_out_0_), .QN(n3627) );
  SDFFX1 s2_msel_pri_out_reg_1_ ( .D(n17427), .SI(s2_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(test_so50), .QN(n3628) );
  SDFFARX1 s3_msel_arb2_state_reg_2_ ( .D(n17458), .SI(s3_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20890), .Q(test_so53), .QN(n3697) );
  SDFFARX1 s3_msel_arb2_state_reg_0_ ( .D(n17460), .SI(s3_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20889), .Q(s3_msel_gnt_p2_0_), .QN(
        n3695) );
  SDFFARX1 s3_msel_arb2_state_reg_1_ ( .D(n17459), .SI(s3_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20889), .Q(s3_msel_gnt_p2_1_), .QN(
        n3696) );
  SDFFARX1 s3_msel_arb0_state_reg_2_ ( .D(n17461), .SI(s3_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20889), .Q(test_so52), .QN(n3681) );
  SDFFARX1 s3_msel_arb0_state_reg_0_ ( .D(n17463), .SI(s3_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20889), .Q(s3_msel_gnt_p0_0_), .QN(n3679) );
  SDFFARX1 s3_msel_arb0_state_reg_1_ ( .D(n17462), .SI(s3_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20889), .Q(s3_msel_gnt_p0_1_), .QN(
        n3680) );
  SDFFARX1 s3_msel_arb1_state_reg_2_ ( .D(n17464), .SI(s3_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20888), .Q(s3_msel_gnt_p1[2]), .QN(
        n3689) );
  SDFFARX1 s3_msel_arb1_state_reg_0_ ( .D(n17466), .SI(test_si53), .SE(test_se), .CLK(clk_i), .RSTB(n20888), .Q(s3_msel_gnt_p1[0]), .QN(n3687) );
  SDFFARX1 s3_msel_arb1_state_reg_1_ ( .D(n17465), .SI(s3_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20888), .Q(s3_msel_gnt_p1[1]), .QN(
        n3688) );
  SDFFARX1 s3_msel_arb3_state_reg_0_ ( .D(n17469), .SI(test_si54), .SE(test_se), .CLK(clk_i), .RSTB(n20888), .Q(s3_msel_gnt_p3[0]), .QN(n3703) );
  SDFFARX1 s3_msel_arb3_state_reg_2_ ( .D(n17467), .SI(s3_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20888), .Q(s3_msel_gnt_p3[2]), .QN(
        n3705) );
  SDFFARX1 s3_msel_arb3_state_reg_1_ ( .D(n17468), .SI(s3_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20887), .Q(s3_msel_gnt_p3[1]), .QN(
        n3704) );
  SDFFX1 s3_next_reg ( .D(n17776), .SI(s3_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(test_so54), .QN() );
  SDFFX1 s3_msel_pri_out_reg_0_ ( .D(n17456), .SI(s3_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s3_msel_pri_out_0_), .QN(n3672) );
  SDFFX1 s3_msel_pri_out_reg_1_ ( .D(n17457), .SI(s3_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s3_msel_pri_out_1_), .QN(n3673) );
  SDFFARX1 s12_msel_arb2_state_reg_2_ ( .D(n17278), .SI(s12_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20887), .Q(s12_msel_gnt_p2[2]), .QN(
        n4102) );
  SDFFARX1 s12_msel_arb2_state_reg_0_ ( .D(n17280), .SI(test_si88), .SE(
        test_se), .CLK(clk_i), .RSTB(n20887), .Q(s12_msel_gnt_p2[0]), .QN(
        n4100) );
  SDFFARX1 s12_msel_arb2_state_reg_1_ ( .D(n17279), .SI(s12_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20887), .Q(s12_msel_gnt_p2[1]), .QN(
        n4101) );
  SDFFARX1 s12_msel_arb0_state_reg_2_ ( .D(n17281), .SI(s12_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20887), .Q(s12_msel_gnt_p0[2]), .QN(
        n4086) );
  SDFFARX1 s12_msel_arb0_state_reg_0_ ( .D(n17283), .SI(test_si87), .SE(
        test_se), .CLK(clk_i), .RSTB(n20886), .Q(s12_msel_gnt_p0[0]), .QN(
        n4084) );
  SDFFARX1 s12_msel_arb0_state_reg_1_ ( .D(n17282), .SI(s12_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20886), .Q(s12_msel_gnt_p0[1]), .QN(
        n4085) );
  SDFFARX1 s12_msel_arb1_state_reg_2_ ( .D(n17284), .SI(s12_msel_gnt_p1_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20886), .Q(test_so87), .QN(n4094) );
  SDFFARX1 s12_msel_arb1_state_reg_0_ ( .D(n17286), .SI(s12_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20886), .Q(s12_msel_gnt_p1_0_), .QN(
        n4092) );
  SDFFARX1 s12_msel_arb1_state_reg_1_ ( .D(n17285), .SI(s12_msel_gnt_p1_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20886), .Q(s12_msel_gnt_p1_1_), .QN(
        n4093) );
  SDFFARX1 s12_msel_arb3_state_reg_0_ ( .D(n17289), .SI(s12_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20885), .Q(s12_msel_gnt_p3_0_), .QN(
        n4108) );
  SDFFARX1 s12_msel_arb3_state_reg_2_ ( .D(n17287), .SI(s12_msel_gnt_p3_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20885), .Q(test_so88), .QN(n4110) );
  SDFFARX1 s12_msel_arb3_state_reg_1_ ( .D(n17288), .SI(s12_msel_gnt_p3_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20885), .Q(s12_msel_gnt_p3_1_), .QN(
        n4109) );
  SDFFX1 s12_next_reg ( .D(n17767), .SI(s12_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s12_next), .QN() );
  SDFFX1 s12_msel_pri_out_reg_0_ ( .D(n17276), .SI(test_si89), .SE(test_se), 
        .CLK(clk_i), .Q(s12_msel_pri_out_0_), .QN(n4077) );
  SDFFX1 s12_msel_pri_out_reg_1_ ( .D(n17277), .SI(s12_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s12_msel_pri_out_1_), .QN(n4078) );
  SDFFARX1 s13_msel_arb2_state_reg_2_ ( .D(n17308), .SI(s13_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20885), .Q(s13_msel_gnt_p2_2_), .QN(
        n4147) );
  SDFFARX1 s13_msel_arb2_state_reg_0_ ( .D(n17310), .SI(s13_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20885), .Q(test_so91), .QN(n4145) );
  SDFFARX1 s13_msel_arb2_state_reg_1_ ( .D(n17309), .SI(test_si92), .SE(
        test_se), .CLK(clk_i), .RSTB(n20884), .Q(s13_msel_gnt_p2_1_), .QN(
        n4146) );
  SDFFARX1 s13_msel_arb0_state_reg_2_ ( .D(n17311), .SI(s13_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20884), .Q(s13_msel_gnt_p0_2_), .QN(
        n4131) );
  SDFFARX1 s13_msel_arb0_state_reg_0_ ( .D(n17313), .SI(s13_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20884), .Q(test_so90), .QN(n4129) );
  SDFFARX1 s13_msel_arb0_state_reg_1_ ( .D(n17312), .SI(test_si91), .SE(
        test_se), .CLK(clk_i), .RSTB(n20884), .Q(s13_msel_gnt_p0_1_), .QN(
        n4130) );
  SDFFARX1 s13_msel_arb1_state_reg_2_ ( .D(n17314), .SI(s13_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20884), .Q(s13_msel_gnt_p1[2]), .QN(
        n4139) );
  SDFFARX1 s13_msel_arb1_state_reg_0_ ( .D(n17316), .SI(s13_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20883), .Q(s13_msel_gnt_p1[0]), .QN(
        n4137) );
  SDFFARX1 s13_msel_arb1_state_reg_1_ ( .D(n17315), .SI(s13_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20883), .Q(s13_msel_gnt_p1[1]), .QN(
        n4138) );
  SDFFARX1 s13_msel_arb3_state_reg_0_ ( .D(n17319), .SI(s13_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20883), .Q(s13_msel_gnt_p3[0]), .QN(
        n4153) );
  SDFFARX1 s13_msel_arb3_state_reg_2_ ( .D(n17317), .SI(s13_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20883), .Q(s13_msel_gnt_p3[2]), .QN(
        n4155) );
  SDFFARX1 s13_msel_arb3_state_reg_1_ ( .D(n17318), .SI(s13_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20883), .Q(s13_msel_gnt_p3[1]), .QN(
        n4154) );
  SDFFX1 s13_next_reg ( .D(n17766), .SI(s13_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s13_next), .QN() );
  SDFFX1 s13_msel_pri_out_reg_0_ ( .D(n17306), .SI(s13_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(test_so92), .QN(n4122) );
  SDFFX1 s13_msel_pri_out_reg_1_ ( .D(n17307), .SI(test_si93), .SE(test_se), 
        .CLK(clk_i), .Q(s13_msel_pri_out_1_), .QN(n4123) );
  SDFFARX1 s4_msel_arb2_state_reg_2_ ( .D(n17488), .SI(s4_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20882), .Q(s4_msel_gnt_p2[2]), .QN(
        n3742) );
  SDFFARX1 s4_msel_arb2_state_reg_0_ ( .D(n17490), .SI(s4_msel_gnt_p1_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20882), .Q(s4_msel_gnt_p2[0]), .QN(
        n3740) );
  SDFFARX1 s4_msel_arb2_state_reg_1_ ( .D(n17489), .SI(s4_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20882), .Q(s4_msel_gnt_p2[1]), .QN(
        n3741) );
  SDFFARX1 s4_msel_arb0_state_reg_2_ ( .D(n17491), .SI(s4_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20882), .Q(s4_msel_gnt_p0[2]), .QN(
        n3726) );
  SDFFARX1 s4_msel_arb0_state_reg_0_ ( .D(n17493), .SI(s4_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20882), .Q(s4_msel_gnt_p0[0]), .QN(n3724) );
  SDFFARX1 s4_msel_arb0_state_reg_1_ ( .D(n17492), .SI(s4_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20881), .Q(s4_msel_gnt_p0[1]), .QN(
        n3725) );
  SDFFARX1 s4_msel_arb1_state_reg_2_ ( .D(n17494), .SI(s4_msel_gnt_p1_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20881), .Q(s4_msel_gnt_p1_2_), .QN(
        n3734) );
  SDFFARX1 s4_msel_arb1_state_reg_0_ ( .D(n17496), .SI(s4_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20881), .Q(test_so56), .QN(n3732) );
  SDFFARX1 s4_msel_arb1_state_reg_1_ ( .D(n17495), .SI(test_si57), .SE(test_se), .CLK(clk_i), .RSTB(n20881), .Q(s4_msel_gnt_p1_1_), .QN(n3733) );
  SDFFARX1 s4_msel_arb3_state_reg_0_ ( .D(n17499), .SI(s4_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20881), .Q(test_so57), .QN(n3748) );
  SDFFARX1 s4_msel_arb3_state_reg_2_ ( .D(n17497), .SI(s4_msel_gnt_p3_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20880), .Q(s4_msel_gnt_p3_2_), .QN(
        n3750) );
  SDFFARX1 s4_msel_arb3_state_reg_1_ ( .D(n17498), .SI(test_si58), .SE(test_se), .CLK(clk_i), .RSTB(n20880), .Q(s4_msel_gnt_p3_1_), .QN(n3749) );
  SDFFX1 s4_next_reg ( .D(n17775), .SI(s4_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s4_next), .QN() );
  SDFFX1 s4_msel_pri_out_reg_0_ ( .D(n17486), .SI(s4_msel_gnt_p3_2_), .SE(
        test_se), .CLK(clk_i), .Q(s4_msel_pri_out_0_), .QN(n3717) );
  SDFFX1 s4_msel_pri_out_reg_1_ ( .D(n17487), .SI(s4_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s4_msel_pri_out_1_), .QN(n3718) );
  SDFFARX1 s5_msel_arb2_state_reg_2_ ( .D(n17518), .SI(s5_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20880), .Q(s5_msel_gnt_p2[2]), .QN(
        n3787) );
  SDFFARX1 s5_msel_arb2_state_reg_0_ ( .D(n17520), .SI(s5_msel_gnt_p1_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20880), .Q(s5_msel_gnt_p2[0]), .QN(
        n3785) );
  SDFFARX1 s5_msel_arb2_state_reg_1_ ( .D(n17519), .SI(s5_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20880), .Q(s5_msel_gnt_p2[1]), .QN(
        n3786) );
  SDFFARX1 s5_msel_arb0_state_reg_2_ ( .D(n17521), .SI(s5_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20879), .Q(s5_msel_gnt_p0[2]), .QN(
        n3771) );
  SDFFARX1 s5_msel_arb0_state_reg_0_ ( .D(n17523), .SI(s5_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20879), .Q(s5_msel_gnt_p0[0]), .QN(n3769) );
  SDFFARX1 s5_msel_arb0_state_reg_1_ ( .D(n17522), .SI(s5_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20879), .Q(s5_msel_gnt_p0[1]), .QN(
        n3770) );
  SDFFARX1 s5_msel_arb1_state_reg_2_ ( .D(n17524), .SI(test_si61), .SE(test_se), .CLK(clk_i), .RSTB(n20879), .Q(s5_msel_gnt_p1_2_), .QN(n3779) );
  SDFFARX1 s5_msel_arb1_state_reg_0_ ( .D(n17526), .SI(s5_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20879), .Q(s5_msel_gnt_p1_0_), .QN(
        n3777) );
  SDFFARX1 s5_msel_arb1_state_reg_1_ ( .D(n17525), .SI(s5_msel_gnt_p1_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20878), .Q(test_so60), .QN(n3778) );
  SDFFARX1 s5_msel_arb3_state_reg_0_ ( .D(n17529), .SI(s5_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20878), .Q(s5_msel_gnt_p3_0_), .QN(
        n3793) );
  SDFFARX1 s5_msel_arb3_state_reg_2_ ( .D(n17527), .SI(test_si62), .SE(test_se), .CLK(clk_i), .RSTB(n20878), .Q(s5_msel_gnt_p3_2_), .QN(n3795) );
  SDFFARX1 s5_msel_arb3_state_reg_1_ ( .D(n17528), .SI(s5_msel_gnt_p3_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20878), .Q(test_so61), .QN(n3794) );
  SDFFX1 s5_next_reg ( .D(n17774), .SI(s5_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s5_next), .QN() );
  SDFFX1 s5_msel_pri_out_reg_0_ ( .D(n17516), .SI(s5_msel_gnt_p3_2_), .SE(
        test_se), .CLK(clk_i), .Q(s5_msel_pri_out_0_), .QN(n3762) );
  SDFFX1 s5_msel_pri_out_reg_1_ ( .D(n17517), .SI(s5_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s5_msel_pri_out_1_), .QN(n3763) );
  SDFFARX1 s14_msel_arb2_state_reg_2_ ( .D(n17338), .SI(test_si96), .SE(
        test_se), .CLK(clk_i), .RSTB(n20878), .Q(s14_msel_gnt_p2_2_), .QN(
        n4192) );
  SDFFARX1 s14_msel_arb2_state_reg_0_ ( .D(n17340), .SI(s14_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20877), .Q(s14_msel_gnt_p2_0_), .QN(
        n4190) );
  SDFFARX1 s14_msel_arb2_state_reg_1_ ( .D(n17339), .SI(s14_msel_gnt_p2_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20877), .Q(test_so95), .QN(n4191) );
  SDFFARX1 s14_msel_arb0_state_reg_2_ ( .D(n17341), .SI(test_si95), .SE(
        test_se), .CLK(clk_i), .RSTB(n20877), .Q(s14_msel_gnt_p0_2_), .QN(
        n4176) );
  SDFFARX1 s14_msel_arb0_state_reg_0_ ( .D(n17343), .SI(s14_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20877), .Q(s14_msel_gnt_p0_0_), .QN(
        n4174) );
  SDFFARX1 s14_msel_arb0_state_reg_1_ ( .D(n17342), .SI(s14_msel_gnt_p0_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20877), .Q(test_so94), .QN(n4175) );
  SDFFARX1 s14_msel_arb1_state_reg_2_ ( .D(n17344), .SI(s14_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20876), .Q(s14_msel_gnt_p1[2]), .QN(
        n4184) );
  SDFFARX1 s14_msel_arb1_state_reg_0_ ( .D(n17346), .SI(s14_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20876), .Q(s14_msel_gnt_p1[0]), .QN(
        n4182) );
  SDFFARX1 s14_msel_arb1_state_reg_1_ ( .D(n17345), .SI(s14_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20876), .Q(s14_msel_gnt_p1[1]), .QN(
        n4183) );
  SDFFARX1 s14_msel_arb3_state_reg_0_ ( .D(n17349), .SI(s14_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20876), .Q(s14_msel_gnt_p3[0]), .QN(
        n4198) );
  SDFFARX1 s14_msel_arb3_state_reg_2_ ( .D(n17347), .SI(s14_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20876), .Q(s14_msel_gnt_p3[2]), .QN(
        n4200) );
  SDFFARX1 s14_msel_arb3_state_reg_1_ ( .D(n17348), .SI(s14_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20875), .Q(s14_msel_gnt_p3[1]), .QN(
        n4199) );
  SDFFX1 s14_next_reg ( .D(n17765), .SI(test_si97), .SE(test_se), .CLK(clk_i), 
        .Q(s14_next), .QN() );
  SDFFX1 s14_msel_pri_out_reg_0_ ( .D(n17336), .SI(s14_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(s14_msel_pri_out_0_), .QN(n4167) );
  SDFFX1 s14_msel_pri_out_reg_1_ ( .D(n17337), .SI(s14_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(test_so96), .QN(n4168) );
  SDFFARX1 s6_msel_arb2_state_reg_2_ ( .D(n17548), .SI(s6_msel_gnt_p2[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20875), .Q(s6_msel_gnt_p2[2]), .QN(
        n3832) );
  SDFFARX1 s6_msel_arb2_state_reg_0_ ( .D(n17550), .SI(test_si65), .SE(test_se), .CLK(clk_i), .RSTB(n20875), .Q(s6_msel_gnt_p2[0]), .QN(n3830) );
  SDFFARX1 s6_msel_arb2_state_reg_1_ ( .D(n17549), .SI(s6_msel_gnt_p2[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20875), .Q(s6_msel_gnt_p2[1]), .QN(
        n3831) );
  SDFFARX1 s6_msel_arb0_state_reg_2_ ( .D(n17551), .SI(s6_msel_gnt_p0[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20875), .Q(s6_msel_gnt_p0[2]), .QN(
        n3816) );
  SDFFARX1 s6_msel_arb0_state_reg_0_ ( .D(n17553), .SI(test_si64), .SE(test_se), .CLK(clk_i), .RSTB(n20874), .Q(s6_msel_gnt_p0[0]), .QN(n3814) );
  SDFFARX1 s6_msel_arb0_state_reg_1_ ( .D(n17552), .SI(s6_msel_gnt_p0[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20874), .Q(s6_msel_gnt_p0[1]), .QN(
        n3815) );
  SDFFARX1 s6_msel_arb1_state_reg_2_ ( .D(n17554), .SI(s6_msel_gnt_p1_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20874), .Q(test_so64), .QN(n3824) );
  SDFFARX1 s6_msel_arb1_state_reg_0_ ( .D(n17556), .SI(s6_msel_gnt_p0[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20874), .Q(s6_msel_gnt_p1_0_), .QN(
        n3822) );
  SDFFARX1 s6_msel_arb1_state_reg_1_ ( .D(n17555), .SI(s6_msel_gnt_p1_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20874), .Q(s6_msel_gnt_p1_1_), .QN(
        n3823) );
  SDFFARX1 s6_msel_arb3_state_reg_0_ ( .D(n17559), .SI(s6_msel_gnt_p2[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20873), .Q(s6_msel_gnt_p3_0_), .QN(
        n3838) );
  SDFFARX1 s6_msel_arb3_state_reg_2_ ( .D(n17557), .SI(s6_msel_gnt_p3_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20873), .Q(test_so65), .QN(n3840) );
  SDFFARX1 s6_msel_arb3_state_reg_1_ ( .D(n17558), .SI(s6_msel_gnt_p3_0_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20873), .Q(s6_msel_gnt_p3_1_), .QN(
        n3839) );
  SDFFX1 s6_next_reg ( .D(n17773), .SI(s6_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s6_next), .QN() );
  SDFFX1 s6_msel_pri_out_reg_0_ ( .D(n17546), .SI(test_si66), .SE(test_se), 
        .CLK(clk_i), .Q(s6_msel_pri_out_0_), .QN(n3807) );
  SDFFX1 s6_msel_pri_out_reg_1_ ( .D(n17547), .SI(s6_msel_pri_out_0_), .SE(
        test_se), .CLK(clk_i), .Q(s6_msel_pri_out_1_), .QN(n3808) );
  SDFFARX1 s7_msel_arb2_state_reg_2_ ( .D(n17578), .SI(s7_msel_gnt_p2_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20873), .Q(s7_msel_gnt_p2_2_), .QN(
        n3877) );
  SDFFARX1 s7_msel_arb2_state_reg_0_ ( .D(n17580), .SI(s7_msel_gnt_p1[2]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20873), .Q(test_so68), .QN(n3875) );
  SDFFARX1 s7_msel_arb2_state_reg_1_ ( .D(n17579), .SI(test_si69), .SE(test_se), .CLK(clk_i), .RSTB(n20872), .Q(s7_msel_gnt_p2_1_), .QN(n3876) );
  SDFFARX1 s7_msel_arb0_state_reg_2_ ( .D(n17581), .SI(s7_msel_gnt_p0_1_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20872), .Q(s7_msel_gnt_p0_2_), .QN(
        n3861) );
  SDFFARX1 s7_msel_arb0_state_reg_0_ ( .D(n17583), .SI(s7_m7_cyc_r), .SE(
        test_se), .CLK(clk_i), .RSTB(n20872), .Q(test_so67), .QN(n3859) );
  SDFFARX1 s7_msel_arb0_state_reg_1_ ( .D(n17582), .SI(test_si68), .SE(test_se), .CLK(clk_i), .RSTB(n20872), .Q(s7_msel_gnt_p0_1_), .QN(n3860) );
  SDFFARX1 s7_msel_arb1_state_reg_2_ ( .D(n17584), .SI(s7_msel_gnt_p1[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20872), .Q(s7_msel_gnt_p1[2]), .QN(
        n3869) );
  SDFFARX1 s7_msel_arb1_state_reg_0_ ( .D(n17586), .SI(s7_msel_gnt_p0_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20871), .Q(s7_msel_gnt_p1[0]), .QN(
        n3867) );
  SDFFARX1 s7_msel_arb1_state_reg_1_ ( .D(n17585), .SI(s7_msel_gnt_p1[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20871), .Q(s7_msel_gnt_p1[1]), .QN(
        n3868) );
  SDFFARX1 s7_msel_arb3_state_reg_0_ ( .D(n17589), .SI(s7_msel_gnt_p2_2_), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20871), .Q(s7_msel_gnt_p3[0]), .QN(
        n3883) );
  SDFFARX1 s7_msel_arb3_state_reg_2_ ( .D(n17587), .SI(s7_msel_gnt_p3[1]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20871), .Q(s7_msel_gnt_p3[2]), .QN(
        n3885) );
  SDFFARX1 s7_msel_arb3_state_reg_1_ ( .D(n17588), .SI(s7_msel_gnt_p3[0]), 
        .SE(test_se), .CLK(clk_i), .RSTB(n20871), .Q(s7_msel_gnt_p3[1]), .QN(
        n3884) );
  SDFFX1 s7_next_reg ( .D(n17772), .SI(s7_msel_pri_out_1_), .SE(test_se), 
        .CLK(clk_i), .Q(s7_next), .QN() );
  SDFFX1 s7_msel_pri_out_reg_0_ ( .D(n17576), .SI(s7_msel_gnt_p3[2]), .SE(
        test_se), .CLK(clk_i), .Q(test_so69), .QN(n3852) );
  SDFFX1 s7_msel_pri_out_reg_1_ ( .D(n17577), .SI(test_si70), .SE(test_se), 
        .CLK(clk_i), .Q(s7_msel_pri_out_1_), .QN(n3853) );
  SDFFX1 rf_rf_ack_reg ( .D(rf_N19), .SI(m7s15_cyc), .SE(test_se), .CLK(clk_i), 
        .Q(rf_rf_ack), .QN() );
  SDFFX1 rf_rf_dout_reg_15_ ( .D(rf_N130), .SI(rf_rf_dout_14_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_15_), .QN() );
  SDFFX1 rf_rf_dout_reg_14_ ( .D(rf_N129), .SI(rf_rf_dout_13_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_14_), .QN() );
  SDFFX1 rf_rf_dout_reg_13_ ( .D(rf_N128), .SI(test_si39), .SE(test_se), .CLK(
        clk_i), .Q(rf_rf_dout_13_), .QN() );
  SDFFX1 rf_rf_dout_reg_12_ ( .D(rf_N127), .SI(rf_rf_dout_11_), .SE(test_se), 
        .CLK(clk_i), .Q(test_so38), .QN() );
  SDFFX1 rf_rf_dout_reg_11_ ( .D(rf_N126), .SI(rf_rf_dout_10_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_11_), .QN() );
  SDFFX1 rf_rf_dout_reg_10_ ( .D(rf_N125), .SI(rf_rf_dout_9_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_10_), .QN() );
  SDFFX1 rf_rf_dout_reg_9_ ( .D(rf_N124), .SI(rf_rf_dout_8_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_9_), .QN() );
  SDFFX1 rf_rf_dout_reg_8_ ( .D(rf_N123), .SI(rf_rf_dout_7_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_8_), .QN() );
  SDFFX1 rf_rf_dout_reg_7_ ( .D(rf_N122), .SI(test_si38), .SE(test_se), .CLK(
        clk_i), .Q(rf_rf_dout_7_), .QN() );
  SDFFX1 rf_rf_dout_reg_6_ ( .D(rf_N121), .SI(rf_rf_dout_5_), .SE(test_se), 
        .CLK(clk_i), .Q(test_so37), .QN() );
  SDFFX1 rf_rf_dout_reg_5_ ( .D(rf_N120), .SI(rf_rf_dout_4_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_5_), .QN() );
  SDFFX1 rf_rf_dout_reg_4_ ( .D(rf_N119), .SI(rf_rf_dout_3_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_4_), .QN() );
  SDFFX1 rf_rf_dout_reg_3_ ( .D(rf_N118), .SI(rf_rf_dout_2_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_3_), .QN() );
  SDFFX1 rf_rf_dout_reg_2_ ( .D(rf_N117), .SI(rf_rf_dout_1_), .SE(test_se), 
        .CLK(clk_i), .Q(rf_rf_dout_2_), .QN() );
  SDFFX1 rf_rf_dout_reg_1_ ( .D(rf_N116), .SI(test_si37), .SE(test_se), .CLK(
        clk_i), .Q(rf_rf_dout_1_), .QN() );
  SDFFX1 rf_rf_dout_reg_0_ ( .D(rf_N115), .SI(rf_rf_ack), .SE(test_se), .CLK(
        clk_i), .Q(test_so36), .QN() );
  LSDNENX1 U18063 ( .D(n9415), .ENB(n9450), .Q(n9447) );
  LSDNENX1 U18070 ( .D(n9726), .ENB(n9761), .Q(n9758) );
  LSDNENX1 U18077 ( .D(n10036), .ENB(n10071), .Q(n10068) );
  LSDNENX1 U18084 ( .D(n10346), .ENB(n10381), .Q(n10378) );
  LSDNENX1 U18091 ( .D(n10655), .ENB(n10690), .Q(n10687) );
  LSDNENX1 U18098 ( .D(n10965), .ENB(n11000), .Q(n10997) );
  LSDNENX1 U18105 ( .D(n11274), .ENB(n11309), .Q(n11306) );
  LSDNENX1 U18112 ( .D(n11584), .ENB(n11619), .Q(n11616) );
  LSDNENX1 U18119 ( .D(n11894), .ENB(n11929), .Q(n11926) );
  LSDNENX1 U18126 ( .D(n12204), .ENB(n12239), .Q(n12236) );
  LSDNENX1 U18133 ( .D(n12513), .ENB(n12548), .Q(n12545) );
  LSDNENX1 U18140 ( .D(n12822), .ENB(n12857), .Q(n12854) );
  LSDNENX1 U18147 ( .D(n13131), .ENB(n13166), .Q(n13163) );
  LSDNENX1 U18154 ( .D(n13440), .ENB(n13475), .Q(n13472) );
  LSDNENX1 U18161 ( .D(n13749), .ENB(n13784), .Q(n13781) );
  LSDNENX1 U18166 ( .D(n14013), .ENB(n14048), .Q(n14045) );
  SDFFARX1 rf_conf0_reg_15_ ( .D(n1586), .SI(test_si1), .SE(test_se), .CLK(
        clk_i), .RSTB(n21079), .Q(conf0_15_), .QN(n18056) );
  SDFFARX1 rf_conf0_reg_13_ ( .D(n1584), .SI(conf0_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20985), .Q(conf0_13_), .QN(n18060) );
  SDFFARX1 rf_conf1_reg_15_ ( .D(n1536), .SI(test_si2), .SE(test_se), .CLK(
        clk_i), .RSTB(n20982), .Q(conf1_15_), .QN(n18208) );
  SDFFARX1 rf_conf1_reg_13_ ( .D(n1534), .SI(conf1_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20982), .Q(conf1_13_), .QN(n18212) );
  SDFFARX1 rf_conf2_reg_15_ ( .D(n1486), .SI(test_si3), .SE(test_se), .CLK(
        clk_i), .RSTB(n20979), .Q(conf2_15_), .QN(n18039) );
  SDFFARX1 rf_conf2_reg_13_ ( .D(n1484), .SI(conf2_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20979), .Q(conf2_13_), .QN(n18043) );
  SDFFARX1 rf_conf3_reg_15_ ( .D(n1436), .SI(test_si4), .SE(test_se), .CLK(
        clk_i), .RSTB(n20976), .Q(conf3_15_), .QN(n18192) );
  SDFFARX1 rf_conf3_reg_13_ ( .D(n1434), .SI(conf3_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20976), .Q(conf3_13_), .QN(n18195) );
  SDFFARX1 rf_conf4_reg_15_ ( .D(n1386), .SI(test_si5), .SE(test_se), .CLK(
        clk_i), .RSTB(n20973), .Q(conf4_15_), .QN(n18053) );
  SDFFARX1 rf_conf4_reg_13_ ( .D(n1384), .SI(conf4_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20972), .Q(conf4_13_), .QN(n18057) );
  SDFFARX1 rf_conf5_reg_15_ ( .D(n1336), .SI(test_si6), .SE(test_se), .CLK(
        clk_i), .RSTB(n20970), .Q(conf5_15_), .QN(n18205) );
  SDFFARX1 rf_conf5_reg_13_ ( .D(n1334), .SI(conf5_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20969), .Q(conf5_13_), .QN(n18209) );
  SDFFARX1 rf_conf6_reg_15_ ( .D(n1286), .SI(test_si7), .SE(test_se), .CLK(
        clk_i), .RSTB(n20966), .Q(conf6_15_), .QN(n18037) );
  SDFFARX1 rf_conf6_reg_13_ ( .D(n1284), .SI(conf6_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20966), .Q(conf6_13_), .QN(n18041) );
  SDFFARX1 rf_conf7_reg_15_ ( .D(n1236), .SI(test_si8), .SE(test_se), .CLK(
        clk_i), .RSTB(n20963), .Q(conf7_15_), .QN(n18191) );
  SDFFARX1 rf_conf7_reg_13_ ( .D(n1234), .SI(conf7_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20963), .Q(conf7_13_), .QN(n18194) );
  SDFFARX1 rf_conf8_reg_15_ ( .D(n1186), .SI(test_si9), .SE(test_se), .CLK(
        clk_i), .RSTB(n20960), .Q(conf8_15_), .QN(n18040) );
  SDFFARX1 rf_conf8_reg_13_ ( .D(n1184), .SI(conf8_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20960), .Q(conf8_13_), .QN(n18044) );
  SDFFARX1 rf_conf9_reg_15_ ( .D(n1136), .SI(test_si10), .SE(test_se), .CLK(
        clk_i), .RSTB(n20957), .Q(conf9_15_), .QN(n18193) );
  SDFFARX1 rf_conf9_reg_13_ ( .D(n1134), .SI(conf9_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20956), .Q(conf9_13_), .QN(n18196) );
  SDFFARX1 rf_conf10_reg_15_ ( .D(n1086), .SI(test_si11), .SE(test_se), .CLK(
        clk_i), .RSTB(n20954), .Q(conf10_15_), .QN(n18055) );
  SDFFARX1 rf_conf10_reg_13_ ( .D(n1084), .SI(conf10_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20953), .Q(conf10_13_), .QN(n18059) );
  SDFFARX1 rf_conf11_reg_15_ ( .D(n1036), .SI(test_si12), .SE(test_se), .CLK(
        clk_i), .RSTB(n20950), .Q(conf11_15_), .QN(n18207) );
  SDFFARX1 rf_conf11_reg_13_ ( .D(n1034), .SI(conf11_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20950), .Q(conf11_13_), .QN(n18211) );
  SDFFARX1 rf_conf12_reg_15_ ( .D(n986), .SI(test_si13), .SE(test_se), .CLK(
        clk_i), .RSTB(n20947), .Q(conf12_15_), .QN(n18054) );
  SDFFARX1 rf_conf12_reg_13_ ( .D(n984), .SI(conf12_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20947), .Q(conf12_13_), .QN(n18058) );
  SDFFARX1 rf_conf13_reg_15_ ( .D(n936), .SI(test_si14), .SE(test_se), .CLK(
        clk_i), .RSTB(n20944), .Q(conf13_15_), .QN(n18206) );
  SDFFARX1 rf_conf13_reg_13_ ( .D(n934), .SI(conf13_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20944), .Q(conf13_13_), .QN(n18210) );
  SDFFARX1 rf_conf14_reg_15_ ( .D(n886), .SI(test_si15), .SE(test_se), .CLK(
        clk_i), .RSTB(n20941), .Q(conf14_15_), .QN(n18038) );
  SDFFARX1 rf_conf14_reg_13_ ( .D(n884), .SI(conf14_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20940), .Q(conf14_13_), .QN(n18042) );
  SDFFARX1 rf_conf15_reg_15_ ( .D(n836), .SI(test_si16), .SE(test_se), .CLK(
        clk_i), .RSTB(n20938), .Q(conf15_15_), .QN(n18189) );
  SDFFARX1 rf_conf15_reg_13_ ( .D(n834), .SI(conf15_14_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20937), .Q(conf15_13_), .QN(n18190) );
  SDFFARX1 rf_conf0_reg_14_ ( .D(n1585), .SI(conf0_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20985), .Q(conf0_14_), .QN(n18220) );
  SDFFARX1 rf_conf1_reg_14_ ( .D(n1535), .SI(conf1_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20982), .Q(conf1_14_), .QN(n18052) );
  SDFFARX1 rf_conf2_reg_14_ ( .D(n1485), .SI(conf2_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20979), .Q(conf2_14_), .QN(n18203) );
  SDFFARX1 rf_conf3_reg_14_ ( .D(n1435), .SI(conf3_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20976), .Q(conf3_14_), .QN(n18033) );
  SDFFARX1 rf_conf4_reg_14_ ( .D(n1385), .SI(conf4_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20973), .Q(conf4_14_), .QN(n18217) );
  SDFFARX1 rf_conf5_reg_14_ ( .D(n1335), .SI(conf5_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20969), .Q(conf5_14_), .QN(n18049) );
  SDFFARX1 rf_conf6_reg_14_ ( .D(n1285), .SI(conf6_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20966), .Q(conf6_14_), .QN(n18201) );
  SDFFARX1 rf_conf7_reg_14_ ( .D(n1235), .SI(conf7_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20963), .Q(conf7_14_), .QN(n18032) );
  SDFFARX1 rf_conf8_reg_14_ ( .D(n1185), .SI(conf8_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20960), .Q(conf8_14_), .QN(n18204) );
  SDFFARX1 rf_conf9_reg_14_ ( .D(n1135), .SI(conf9_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20957), .Q(conf9_14_), .QN(n18034) );
  SDFFARX1 rf_conf10_reg_14_ ( .D(n1085), .SI(conf10_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20953), .Q(conf10_14_), .QN(n18219) );
  SDFFARX1 rf_conf11_reg_14_ ( .D(n1035), .SI(conf11_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20950), .Q(conf11_14_), .QN(n18051) );
  SDFFARX1 rf_conf12_reg_14_ ( .D(n985), .SI(conf12_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20947), .Q(conf12_14_), .QN(n18218) );
  SDFFARX1 rf_conf13_reg_14_ ( .D(n935), .SI(conf13_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20944), .Q(conf13_14_), .QN(n18050) );
  SDFFARX1 rf_conf14_reg_14_ ( .D(n885), .SI(conf14_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20941), .Q(conf14_14_), .QN(n18202) );
  SDFFARX1 rf_conf15_reg_14_ ( .D(n835), .SI(conf15_15_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20937), .Q(conf15_14_), .QN(n18036) );
  SDFFARX1 rf_conf15_reg_12_ ( .D(n833), .SI(conf15_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20937), .Q(conf15_12_), .QN(n18035) );
  SDFFARX1 rf_conf0_reg_12_ ( .D(n1583), .SI(conf0_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20985), .Q(conf0_12_), .QN(n18216) );
  SDFFARX1 rf_conf1_reg_12_ ( .D(n1533), .SI(conf1_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20982), .Q(conf1_12_), .QN(n18048) );
  SDFFARX1 rf_conf2_reg_12_ ( .D(n1483), .SI(conf2_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20979), .Q(conf2_12_), .QN(n18199) );
  SDFFARX1 rf_conf3_reg_12_ ( .D(n1433), .SI(conf3_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20975), .Q(conf3_12_), .QN(n18030) );
  SDFFARX1 rf_conf4_reg_12_ ( .D(n1383), .SI(conf4_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20972), .Q(conf4_12_), .QN(n18213) );
  SDFFARX1 rf_conf5_reg_12_ ( .D(n1333), .SI(conf5_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20969), .Q(conf5_12_), .QN(n18045) );
  SDFFARX1 rf_conf6_reg_12_ ( .D(n1283), .SI(conf6_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20966), .Q(conf6_12_), .QN(n18197) );
  SDFFARX1 rf_conf7_reg_12_ ( .D(n1233), .SI(conf7_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20963), .Q(conf7_12_), .QN(n18029) );
  SDFFARX1 rf_conf8_reg_12_ ( .D(n1183), .SI(conf8_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20959), .Q(conf8_12_), .QN(n18200) );
  SDFFARX1 rf_conf9_reg_12_ ( .D(n1133), .SI(conf9_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20956), .Q(conf9_12_), .QN(n18031) );
  SDFFARX1 rf_conf10_reg_12_ ( .D(n1083), .SI(conf10_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20953), .Q(conf10_12_), .QN(n18215) );
  SDFFARX1 rf_conf11_reg_12_ ( .D(n1033), .SI(conf11_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20950), .Q(conf11_12_), .QN(n18047) );
  SDFFARX1 rf_conf12_reg_12_ ( .D(n983), .SI(conf12_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20947), .Q(conf12_12_), .QN(n18214) );
  SDFFARX1 rf_conf13_reg_12_ ( .D(n933), .SI(conf13_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20943), .Q(conf13_12_), .QN(n18046) );
  SDFFARX1 rf_conf14_reg_12_ ( .D(n883), .SI(conf14_13_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20940), .Q(conf14_12_), .QN(n18198) );
  SDFFARX1 rf_conf0_reg_7_ ( .D(n1578), .SI(conf0_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20984), .Q(conf0_7_), .QN(n18012) );
  SDFFARX1 rf_conf0_reg_5_ ( .D(n1576), .SI(conf0_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20984), .Q(conf0_5_), .QN(n18011) );
  SDFFARX1 rf_conf1_reg_7_ ( .D(n1528), .SI(conf1_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20981), .Q(conf1_7_), .QN(n18121) );
  SDFFARX1 rf_conf1_reg_5_ ( .D(n1526), .SI(conf1_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20980), .Q(conf1_5_), .QN(n18120) );
  SDFFARX1 rf_conf2_reg_7_ ( .D(n1478), .SI(conf2_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20978), .Q(conf2_7_), .QN(n17982) );
  SDFFARX1 rf_conf2_reg_5_ ( .D(n1476), .SI(conf2_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20977), .Q(conf2_5_), .QN(n17981) );
  SDFFARX1 rf_conf3_reg_7_ ( .D(n1428), .SI(conf3_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20974), .Q(conf3_7_), .QN(n18092) );
  SDFFARX1 rf_conf3_reg_5_ ( .D(n1426), .SI(conf3_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20974), .Q(conf3_5_), .QN(n18091) );
  SDFFARX1 rf_conf4_reg_7_ ( .D(n1378), .SI(conf4_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20971), .Q(conf4_7_), .QN(n18006) );
  SDFFARX1 rf_conf4_reg_5_ ( .D(n1376), .SI(conf4_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20971), .Q(conf4_5_), .QN(n18005) );
  SDFFARX1 rf_conf5_reg_7_ ( .D(n1328), .SI(conf5_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20968), .Q(conf5_7_), .QN(n18115) );
  SDFFARX1 rf_conf5_reg_5_ ( .D(n1326), .SI(conf5_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20968), .Q(conf5_5_), .QN(n18114) );
  SDFFARX1 rf_conf6_reg_7_ ( .D(n1278), .SI(conf6_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20965), .Q(conf6_7_), .QN(n17978) );
  SDFFARX1 rf_conf7_reg_7_ ( .D(n1228), .SI(conf7_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20962), .Q(conf7_7_), .QN(n18090) );
  SDFFARX1 rf_conf7_reg_5_ ( .D(n1226), .SI(conf7_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20961), .Q(conf7_5_), .QN(n18089) );
  SDFFARX1 rf_conf8_reg_7_ ( .D(n1178), .SI(conf8_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20958), .Q(conf8_7_), .QN(n17984) );
  SDFFARX1 rf_conf8_reg_5_ ( .D(n1176), .SI(conf8_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20958), .Q(conf8_5_), .QN(n17983) );
  SDFFARX1 rf_conf9_reg_7_ ( .D(n1128), .SI(conf9_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20955), .Q(conf9_7_), .QN(n18094) );
  SDFFARX1 rf_conf10_reg_7_ ( .D(n1078), .SI(conf10_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20952), .Q(conf10_7_), .QN(n18010) );
  SDFFARX1 rf_conf10_reg_5_ ( .D(n1076), .SI(conf10_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20952), .Q(conf10_5_), .QN(n18009) );
  SDFFARX1 rf_conf11_reg_7_ ( .D(n1028), .SI(conf11_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20949), .Q(conf11_7_), .QN(n18119) );
  SDFFARX1 rf_conf12_reg_7_ ( .D(n978), .SI(conf12_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20946), .Q(conf12_7_), .QN(n18008) );
  SDFFARX1 rf_conf12_reg_5_ ( .D(n976), .SI(conf12_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20945), .Q(conf12_5_), .QN(n18007) );
  SDFFARX1 rf_conf13_reg_7_ ( .D(n928), .SI(conf13_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20942), .Q(conf13_7_), .QN(n18117) );
  SDFFARX1 rf_conf14_reg_7_ ( .D(n878), .SI(conf14_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20939), .Q(conf14_7_), .QN(n17980) );
  SDFFARX1 rf_conf14_reg_5_ ( .D(n876), .SI(conf14_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20939), .Q(conf14_5_), .QN(n17979) );
  SDFFARX1 rf_conf15_reg_7_ ( .D(n828), .SI(conf15_8_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20936), .Q(conf15_7_), .QN(n18087) );
  SDFFARX1 rf_conf15_reg_5_ ( .D(n826), .SI(conf15_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20936), .Q(conf15_5_), .QN(n18086) );
  SDFFARX1 rf_conf0_reg_6_ ( .D(n1577), .SI(conf0_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20984), .Q(conf0_6_), .QN(n18133) );
  SDFFARX1 rf_conf1_reg_6_ ( .D(n1527), .SI(conf1_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20981), .Q(conf1_6_), .QN(n17996) );
  SDFFARX1 rf_conf2_reg_6_ ( .D(n1477), .SI(conf2_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20977), .Q(conf2_6_), .QN(n18104) );
  SDFFARX1 rf_conf3_reg_6_ ( .D(n1427), .SI(conf3_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20974), .Q(conf3_6_), .QN(n17966) );
  SDFFARX1 rf_conf4_reg_6_ ( .D(n1377), .SI(conf4_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20971), .Q(conf4_6_), .QN(n18130) );
  SDFFARX1 rf_conf5_reg_6_ ( .D(n1327), .SI(conf5_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20968), .Q(conf5_6_), .QN(n17993) );
  SDFFARX1 rf_conf6_reg_6_ ( .D(n1277), .SI(conf6_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20965), .Q(conf6_6_), .QN(n18102) );
  SDFFARX1 rf_conf7_reg_6_ ( .D(n1227), .SI(conf7_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20961), .Q(conf7_6_), .QN(n17965) );
  SDFFARX1 rf_conf8_reg_6_ ( .D(n1177), .SI(conf8_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20958), .Q(conf8_6_), .QN(n18105) );
  SDFFARX1 rf_conf9_reg_6_ ( .D(n1127), .SI(conf9_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20955), .Q(conf9_6_), .QN(n17967) );
  SDFFARX1 rf_conf10_reg_6_ ( .D(n1077), .SI(conf10_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20952), .Q(conf10_6_), .QN(n18132) );
  SDFFARX1 rf_conf11_reg_6_ ( .D(n1027), .SI(conf11_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20949), .Q(conf11_6_), .QN(n17995) );
  SDFFARX1 rf_conf12_reg_6_ ( .D(n977), .SI(conf12_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20945), .Q(conf12_6_), .QN(n18131) );
  SDFFARX1 rf_conf13_reg_6_ ( .D(n927), .SI(conf13_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20942), .Q(conf13_6_), .QN(n17994) );
  SDFFARX1 rf_conf14_reg_6_ ( .D(n877), .SI(conf14_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20939), .Q(conf14_6_), .QN(n18103) );
  SDFFARX1 rf_conf15_reg_6_ ( .D(n827), .SI(conf15_7_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20936), .Q(conf15_6_), .QN(n17976) );
  SDFFARX1 rf_conf0_reg_11_ ( .D(n1582), .SI(conf0_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20985), .Q(conf0_11_), .QN(n18082) );
  SDFFARX1 rf_conf1_reg_11_ ( .D(n1532), .SI(conf1_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20982), .Q(conf1_11_), .QN(n17963) );
  SDFFARX1 rf_conf2_reg_11_ ( .D(n1482), .SI(conf2_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20978), .Q(conf2_11_), .QN(n18077) );
  SDFFARX1 rf_conf3_reg_11_ ( .D(n1432), .SI(conf3_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20975), .Q(conf3_11_), .QN(n17951) );
  SDFFARX1 rf_conf4_reg_11_ ( .D(n1382), .SI(conf4_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20972), .Q(conf4_11_), .QN(n18079) );
  SDFFARX1 rf_conf5_reg_11_ ( .D(n1332), .SI(conf5_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20969), .Q(conf5_11_), .QN(n17960) );
  SDFFARX1 rf_conf6_reg_11_ ( .D(n1282), .SI(conf6_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20966), .Q(conf6_11_), .QN(n18075) );
  SDFFARX1 rf_conf7_reg_11_ ( .D(n1232), .SI(conf7_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20962), .Q(conf7_11_), .QN(n17950) );
  SDFFARX1 rf_conf8_reg_11_ ( .D(n1182), .SI(conf8_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20959), .Q(conf8_11_), .QN(n18078) );
  SDFFARX1 rf_conf9_reg_11_ ( .D(n1132), .SI(conf9_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20956), .Q(conf9_11_), .QN(n17952) );
  SDFFARX1 rf_conf10_reg_11_ ( .D(n1082), .SI(conf10_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20953), .Q(conf10_11_), .QN(n18081) );
  SDFFARX1 rf_conf11_reg_11_ ( .D(n1032), .SI(conf11_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20950), .Q(conf11_11_), .QN(n17962) );
  SDFFARX1 rf_conf12_reg_11_ ( .D(n982), .SI(conf12_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20946), .Q(conf12_11_), .QN(n18080) );
  SDFFARX1 rf_conf13_reg_11_ ( .D(n932), .SI(conf13_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20943), .Q(conf13_11_), .QN(n17961) );
  SDFFARX1 rf_conf14_reg_11_ ( .D(n882), .SI(conf14_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20940), .Q(conf14_11_), .QN(n18076) );
  SDFFARX1 rf_conf15_reg_11_ ( .D(n832), .SI(conf15_12_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20937), .Q(conf15_11_), .QN(n17949) );
  SDFFARX1 rf_conf0_reg_10_ ( .D(n1581), .SI(conf0_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20985), .Q(conf0_10_), .QN(n17956) );
  SDFFARX1 rf_conf1_reg_10_ ( .D(n1531), .SI(conf1_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20981), .Q(conf1_10_), .QN(n18074) );
  SDFFARX1 rf_conf2_reg_10_ ( .D(n1481), .SI(conf2_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20978), .Q(conf2_10_), .QN(n17943) );
  SDFFARX1 rf_conf3_reg_10_ ( .D(n1431), .SI(conf3_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20975), .Q(conf3_10_), .QN(n18067) );
  SDFFARX1 rf_conf4_reg_10_ ( .D(n1381), .SI(conf4_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20972), .Q(conf4_10_), .QN(n17953) );
  SDFFARX1 rf_conf5_reg_10_ ( .D(n1331), .SI(conf5_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20969), .Q(conf5_10_), .QN(n18071) );
  SDFFARX1 rf_conf6_reg_10_ ( .D(n1281), .SI(conf6_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20965), .Q(conf6_10_), .QN(n17941) );
  SDFFARX1 rf_conf7_reg_10_ ( .D(n1231), .SI(conf7_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20962), .Q(conf7_10_), .QN(n18069) );
  SDFFARX1 rf_conf8_reg_10_ ( .D(n1181), .SI(conf8_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20959), .Q(conf8_10_), .QN(n17944) );
  SDFFARX1 rf_conf9_reg_10_ ( .D(n1131), .SI(conf9_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20956), .Q(conf9_10_), .QN(n18068) );
  SDFFARX1 rf_conf10_reg_10_ ( .D(n1081), .SI(conf10_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20953), .Q(conf10_10_), .QN(n17955) );
  SDFFARX1 rf_conf11_reg_10_ ( .D(n1031), .SI(conf11_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20949), .Q(conf11_10_), .QN(n18073) );
  SDFFARX1 rf_conf12_reg_10_ ( .D(n981), .SI(conf12_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20946), .Q(conf12_10_), .QN(n17954) );
  SDFFARX1 rf_conf13_reg_10_ ( .D(n931), .SI(conf13_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20943), .Q(conf13_10_), .QN(n18072) );
  SDFFARX1 rf_conf14_reg_10_ ( .D(n881), .SI(conf14_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20940), .Q(conf14_10_), .QN(n17942) );
  SDFFARX1 rf_conf15_reg_10_ ( .D(n831), .SI(conf15_11_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20937), .Q(conf15_10_), .QN(n18070) );
  SDFFARX1 rf_conf0_reg_0_ ( .D(n1571), .SI(conf0_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20983), .Q(test_so1), .QN(n18149) );
  SDFFARX1 rf_conf1_reg_0_ ( .D(n1521), .SI(conf1_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20979), .Q(test_so2), .QN(n18028) );
  SDFFARX1 rf_conf2_reg_0_ ( .D(n1471), .SI(conf2_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20976), .Q(test_so3), .QN(n18144) );
  SDFFARX1 rf_conf3_reg_0_ ( .D(n1421), .SI(conf3_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20973), .Q(test_so4), .QN(n18022) );
  SDFFARX1 rf_conf4_reg_0_ ( .D(n1371), .SI(conf4_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20970), .Q(test_so5), .QN(n18146) );
  SDFFARX1 rf_conf5_reg_0_ ( .D(n1321), .SI(conf5_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20967), .Q(test_so6), .QN(n18025) );
  SDFFARX1 rf_conf6_reg_0_ ( .D(n1271), .SI(conf6_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20963), .Q(test_so7), .QN(n18142) );
  SDFFARX1 rf_conf7_reg_0_ ( .D(n1221), .SI(conf7_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20960), .Q(test_so8), .QN(n18021) );
  SDFFARX1 rf_conf8_reg_0_ ( .D(n1171), .SI(conf8_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20957), .Q(test_so9), .QN(n18145) );
  SDFFARX1 rf_conf9_reg_0_ ( .D(n1121), .SI(conf9_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20954), .Q(test_so10), .QN(n18023) );
  SDFFARX1 rf_conf10_reg_0_ ( .D(n1071), .SI(conf10_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20951), .Q(test_so11), .QN(n18148) );
  SDFFARX1 rf_conf11_reg_0_ ( .D(n1021), .SI(conf11_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20947), .Q(test_so12), .QN(n18027) );
  SDFFARX1 rf_conf12_reg_0_ ( .D(n971), .SI(conf12_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20944), .Q(test_so13), .QN(n18147) );
  SDFFARX1 rf_conf13_reg_0_ ( .D(n921), .SI(conf13_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20941), .Q(test_so14), .QN(n18026) );
  SDFFARX1 rf_conf14_reg_0_ ( .D(n871), .SI(conf14_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20938), .Q(test_so15), .QN(n18143) );
  SDFFARX1 rf_conf15_reg_0_ ( .D(n821), .SI(conf15_1_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20935), .Q(test_so16), .QN(n18024) );
  SDFFARX1 rf_conf0_reg_3_ ( .D(n1574), .SI(conf0_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20983), .Q(conf0_3_), .QN(n18016) );
  SDFFARX1 rf_conf0_reg_1_ ( .D(n1572), .SI(conf0_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20983), .Q(conf0_1_), .QN(n18020) );
  SDFFARX1 rf_conf1_reg_3_ ( .D(n1524), .SI(conf1_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20980), .Q(conf1_3_), .QN(n18125) );
  SDFFARX1 rf_conf1_reg_1_ ( .D(n1522), .SI(conf1_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20980), .Q(conf1_1_), .QN(n18129) );
  SDFFARX1 rf_conf2_reg_3_ ( .D(n1474), .SI(conf2_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20977), .Q(conf2_3_), .QN(n17987) );
  SDFFARX1 rf_conf2_reg_1_ ( .D(n1472), .SI(conf2_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20976), .Q(conf2_1_), .QN(n17991) );
  SDFFARX1 rf_conf3_reg_3_ ( .D(n1424), .SI(conf3_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20974), .Q(conf3_3_), .QN(n18096) );
  SDFFARX1 rf_conf3_reg_1_ ( .D(n1422), .SI(conf3_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20973), .Q(conf3_1_), .QN(n18100) );
  SDFFARX1 rf_conf4_reg_3_ ( .D(n1374), .SI(conf4_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20970), .Q(conf4_3_), .QN(n18013) );
  SDFFARX1 rf_conf4_reg_1_ ( .D(n1372), .SI(conf4_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20970), .Q(conf4_1_), .QN(n18017) );
  SDFFARX1 rf_conf5_reg_3_ ( .D(n1324), .SI(conf5_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20967), .Q(conf5_3_), .QN(n18122) );
  SDFFARX1 rf_conf5_reg_1_ ( .D(n1322), .SI(conf5_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20967), .Q(conf5_1_), .QN(n18126) );
  SDFFARX1 rf_conf6_reg_5_ ( .D(n1276), .SI(conf6_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20964), .Q(conf6_5_), .QN(n17977) );
  SDFFARX1 rf_conf6_reg_3_ ( .D(n1274), .SI(conf6_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20964), .Q(conf6_3_), .QN(n17985) );
  SDFFARX1 rf_conf6_reg_1_ ( .D(n1272), .SI(conf6_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20964), .Q(conf6_1_), .QN(n17989) );
  SDFFARX1 rf_conf7_reg_3_ ( .D(n1224), .SI(conf7_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20961), .Q(conf7_3_), .QN(n18095) );
  SDFFARX1 rf_conf7_reg_1_ ( .D(n1222), .SI(conf7_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20960), .Q(conf7_1_), .QN(n18099) );
  SDFFARX1 rf_conf8_reg_3_ ( .D(n1174), .SI(conf8_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20958), .Q(conf8_3_), .QN(n17988) );
  SDFFARX1 rf_conf8_reg_1_ ( .D(n1172), .SI(conf8_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20957), .Q(conf8_1_), .QN(n17992) );
  SDFFARX1 rf_conf9_reg_5_ ( .D(n1126), .SI(conf9_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20955), .Q(conf9_5_), .QN(n18093) );
  SDFFARX1 rf_conf9_reg_3_ ( .D(n1124), .SI(conf9_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20954), .Q(conf9_3_), .QN(n18097) );
  SDFFARX1 rf_conf9_reg_1_ ( .D(n1122), .SI(conf9_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20954), .Q(conf9_1_), .QN(n18101) );
  SDFFARX1 rf_conf10_reg_3_ ( .D(n1074), .SI(conf10_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20951), .Q(conf10_3_), .QN(n18015) );
  SDFFARX1 rf_conf10_reg_1_ ( .D(n1072), .SI(conf10_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20951), .Q(conf10_1_), .QN(n18019) );
  SDFFARX1 rf_conf11_reg_5_ ( .D(n1026), .SI(conf11_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20948), .Q(conf11_5_), .QN(n18118) );
  SDFFARX1 rf_conf11_reg_3_ ( .D(n1024), .SI(conf11_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20948), .Q(conf11_3_), .QN(n18124) );
  SDFFARX1 rf_conf11_reg_1_ ( .D(n1022), .SI(conf11_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20948), .Q(conf11_1_), .QN(n18128) );
  SDFFARX1 rf_conf12_reg_3_ ( .D(n974), .SI(conf12_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20945), .Q(conf12_3_), .QN(n18014) );
  SDFFARX1 rf_conf12_reg_1_ ( .D(n972), .SI(conf12_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20944), .Q(conf12_1_), .QN(n18018) );
  SDFFARX1 rf_conf13_reg_5_ ( .D(n926), .SI(conf13_6_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20942), .Q(conf13_5_), .QN(n18116) );
  SDFFARX1 rf_conf13_reg_3_ ( .D(n924), .SI(conf13_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20942), .Q(conf13_3_), .QN(n18123) );
  SDFFARX1 rf_conf13_reg_1_ ( .D(n922), .SI(conf13_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20941), .Q(conf13_1_), .QN(n18127) );
  SDFFARX1 rf_conf14_reg_3_ ( .D(n874), .SI(conf14_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20938), .Q(conf14_3_), .QN(n17986) );
  SDFFARX1 rf_conf14_reg_1_ ( .D(n872), .SI(conf14_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20938), .Q(conf14_1_), .QN(n17990) );
  SDFFARX1 rf_conf15_reg_9_ ( .D(n830), .SI(conf15_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20936), .Q(conf15_9_), .QN(n17939) );
  SDFFARX1 rf_conf15_reg_3_ ( .D(n824), .SI(conf15_4_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20935), .Q(conf15_3_), .QN(n18088) );
  SDFFARX1 rf_conf15_reg_1_ ( .D(n822), .SI(conf15_2_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20935), .Q(conf15_1_), .QN(n18098) );
  SDFFARX1 rf_conf0_reg_4_ ( .D(n1575), .SI(conf0_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20983), .Q(conf0_4_), .QN(n18141) );
  SDFFARX1 rf_conf0_reg_2_ ( .D(n1573), .SI(conf0_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20983), .Q(conf0_2_), .QN(n18140) );
  SDFFARX1 rf_conf1_reg_4_ ( .D(n1525), .SI(conf1_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20980), .Q(conf1_4_), .QN(n18004) );
  SDFFARX1 rf_conf1_reg_2_ ( .D(n1523), .SI(conf1_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20980), .Q(conf1_2_), .QN(n18003) );
  SDFFARX1 rf_conf2_reg_4_ ( .D(n1475), .SI(conf2_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20977), .Q(conf2_4_), .QN(n18111) );
  SDFFARX1 rf_conf2_reg_2_ ( .D(n1473), .SI(conf2_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20977), .Q(conf2_2_), .QN(n18110) );
  SDFFARX1 rf_conf3_reg_4_ ( .D(n1425), .SI(conf3_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20974), .Q(conf3_4_), .QN(n17971) );
  SDFFARX1 rf_conf3_reg_2_ ( .D(n1423), .SI(conf3_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20973), .Q(conf3_2_), .QN(n17970) );
  SDFFARX1 rf_conf4_reg_4_ ( .D(n1375), .SI(conf4_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20971), .Q(conf4_4_), .QN(n18135) );
  SDFFARX1 rf_conf4_reg_2_ ( .D(n1373), .SI(conf4_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20970), .Q(conf4_2_), .QN(n18134) );
  SDFFARX1 rf_conf5_reg_4_ ( .D(n1325), .SI(conf5_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20967), .Q(conf5_4_), .QN(n17998) );
  SDFFARX1 rf_conf5_reg_2_ ( .D(n1323), .SI(conf5_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20967), .Q(conf5_2_), .QN(n17997) );
  SDFFARX1 rf_conf6_reg_4_ ( .D(n1275), .SI(conf6_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20964), .Q(conf6_4_), .QN(n18107) );
  SDFFARX1 rf_conf6_reg_2_ ( .D(n1273), .SI(conf6_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20964), .Q(conf6_2_), .QN(n18106) );
  SDFFARX1 rf_conf7_reg_4_ ( .D(n1225), .SI(conf7_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20961), .Q(conf7_4_), .QN(n17969) );
  SDFFARX1 rf_conf7_reg_2_ ( .D(n1223), .SI(conf7_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20961), .Q(conf7_2_), .QN(n17968) );
  SDFFARX1 rf_conf8_reg_4_ ( .D(n1175), .SI(conf8_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20958), .Q(conf8_4_), .QN(n18113) );
  SDFFARX1 rf_conf8_reg_2_ ( .D(n1173), .SI(conf8_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20957), .Q(conf8_2_), .QN(n18112) );
  SDFFARX1 rf_conf9_reg_4_ ( .D(n1125), .SI(conf9_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20955), .Q(conf9_4_), .QN(n17973) );
  SDFFARX1 rf_conf9_reg_2_ ( .D(n1123), .SI(conf9_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20954), .Q(conf9_2_), .QN(n17972) );
  SDFFARX1 rf_conf10_reg_4_ ( .D(n1075), .SI(conf10_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20951), .Q(conf10_4_), .QN(n18139) );
  SDFFARX1 rf_conf10_reg_2_ ( .D(n1073), .SI(conf10_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20951), .Q(conf10_2_), .QN(n18138) );
  SDFFARX1 rf_conf11_reg_4_ ( .D(n1025), .SI(conf11_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20948), .Q(conf11_4_), .QN(n18002) );
  SDFFARX1 rf_conf11_reg_2_ ( .D(n1023), .SI(conf11_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20948), .Q(conf11_2_), .QN(n18001) );
  SDFFARX1 rf_conf12_reg_4_ ( .D(n975), .SI(conf12_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20945), .Q(conf12_4_), .QN(n18137) );
  SDFFARX1 rf_conf12_reg_2_ ( .D(n973), .SI(conf12_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20945), .Q(conf12_2_), .QN(n18136) );
  SDFFARX1 rf_conf13_reg_4_ ( .D(n925), .SI(conf13_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20942), .Q(conf13_4_), .QN(n18000) );
  SDFFARX1 rf_conf13_reg_2_ ( .D(n923), .SI(conf13_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20941), .Q(conf13_2_), .QN(n17999) );
  SDFFARX1 rf_conf14_reg_4_ ( .D(n875), .SI(conf14_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20939), .Q(conf14_4_), .QN(n18109) );
  SDFFARX1 rf_conf14_reg_2_ ( .D(n873), .SI(conf14_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20938), .Q(conf14_2_), .QN(n18108) );
  SDFFARX1 rf_conf15_reg_8_ ( .D(n829), .SI(conf15_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20936), .Q(conf15_8_), .QN(n18150) );
  SDFFARX1 rf_conf15_reg_4_ ( .D(n825), .SI(conf15_5_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20935), .Q(conf15_4_), .QN(n17974) );
  SDFFARX1 rf_conf15_reg_2_ ( .D(n823), .SI(conf15_3_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20935), .Q(conf15_2_), .QN(n17975) );
  SDFFARX1 rf_conf0_reg_9_ ( .D(n1580), .SI(conf0_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20984), .Q(conf0_9_), .QN(n17959) );
  SDFFARX1 rf_conf1_reg_9_ ( .D(n1530), .SI(conf1_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20981), .Q(conf1_9_), .QN(n18064) );
  SDFFARX1 rf_conf2_reg_9_ ( .D(n1480), .SI(conf2_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20978), .Q(conf2_9_), .QN(n18154) );
  SDFFARX1 rf_conf3_reg_9_ ( .D(n1430), .SI(conf3_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20975), .Q(conf3_9_), .QN(n17945) );
  SDFFARX1 rf_conf4_reg_9_ ( .D(n1380), .SI(conf4_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20972), .Q(conf4_9_), .QN(n17934) );
  SDFFARX1 rf_conf5_reg_9_ ( .D(n1330), .SI(conf5_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20968), .Q(conf5_9_), .QN(n18063) );
  SDFFARX1 rf_conf6_reg_9_ ( .D(n1280), .SI(conf6_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20965), .Q(conf6_9_), .QN(n18155) );
  SDFFARX1 rf_conf7_reg_9_ ( .D(n1230), .SI(conf7_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20962), .Q(conf7_9_), .QN(n17964) );
  SDFFARX1 rf_conf8_reg_9_ ( .D(n1180), .SI(conf8_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20959), .Q(conf8_9_), .QN(n17933) );
  SDFFARX1 rf_conf9_reg_9_ ( .D(n1130), .SI(conf9_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20956), .Q(conf9_9_), .QN(n18153) );
  SDFFARX1 rf_conf10_reg_9_ ( .D(n1080), .SI(conf10_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20952), .Q(conf10_9_), .QN(n17957) );
  SDFFARX1 rf_conf11_reg_9_ ( .D(n1030), .SI(conf11_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20949), .Q(conf11_9_), .QN(n18061) );
  SDFFARX1 rf_conf12_reg_9_ ( .D(n980), .SI(conf12_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20946), .Q(conf12_9_), .QN(n17958) );
  SDFFARX1 rf_conf13_reg_9_ ( .D(n930), .SI(conf13_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20943), .Q(conf13_9_), .QN(n18062) );
  SDFFARX1 rf_conf14_reg_9_ ( .D(n880), .SI(conf14_10_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20940), .Q(conf14_9_), .QN(n18156) );
  SDFFARX1 rf_conf0_reg_8_ ( .D(n1579), .SI(conf0_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20984), .Q(conf0_8_), .QN(n18085) );
  SDFFARX1 rf_conf1_reg_8_ ( .D(n1529), .SI(conf1_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20981), .Q(conf1_8_), .QN(n17938) );
  SDFFARX1 rf_conf2_reg_8_ ( .D(n1479), .SI(conf2_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20978), .Q(conf2_8_), .QN(n17946) );
  SDFFARX1 rf_conf3_reg_8_ ( .D(n1429), .SI(conf3_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20975), .Q(conf3_8_), .QN(n18151) );
  SDFFARX1 rf_conf4_reg_8_ ( .D(n1379), .SI(conf4_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20971), .Q(conf4_8_), .QN(n18066) );
  SDFFARX1 rf_conf5_reg_8_ ( .D(n1329), .SI(conf5_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20968), .Q(conf5_8_), .QN(n17935) );
  SDFFARX1 rf_conf6_reg_8_ ( .D(n1279), .SI(conf6_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20965), .Q(conf6_8_), .QN(n17947) );
  SDFFARX1 rf_conf7_reg_8_ ( .D(n1229), .SI(conf7_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20962), .Q(conf7_8_), .QN(n18152) );
  SDFFARX1 rf_conf8_reg_8_ ( .D(n1179), .SI(conf8_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20959), .Q(conf8_8_), .QN(n18065) );
  SDFFARX1 rf_conf9_reg_8_ ( .D(n1129), .SI(conf9_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20955), .Q(conf9_8_), .QN(n17940) );
  SDFFARX1 rf_conf10_reg_8_ ( .D(n1079), .SI(conf10_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20952), .Q(conf10_8_), .QN(n18084) );
  SDFFARX1 rf_conf11_reg_8_ ( .D(n1029), .SI(conf11_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20949), .Q(conf11_8_), .QN(n17937) );
  SDFFARX1 rf_conf12_reg_8_ ( .D(n979), .SI(conf12_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20946), .Q(conf12_8_), .QN(n18083) );
  SDFFARX1 rf_conf13_reg_8_ ( .D(n929), .SI(conf13_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20943), .Q(conf13_8_), .QN(n17936) );
  SDFFARX1 rf_conf14_reg_8_ ( .D(n879), .SI(conf14_9_), .SE(test_se), .CLK(
        clk_i), .RSTB(n20939), .Q(conf14_8_), .QN(n17948) );
  SDFFARX1 m5_s6_cyc_o_reg ( .D(n17674), .SI(m5s5_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20917), .Q(m5s6_cyc), .QN(n18304) );
  SDFFARX1 m5_s13_cyc_o_reg ( .D(n17681), .SI(m5s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20918), .Q(test_so30), .QN(n18308) );
  SDFFARX1 m5_s11_cyc_o_reg ( .D(n17679), .SI(m5s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20918), .Q(m5s11_cyc), .QN(n18312) );
  SDFFARX1 m5_s9_cyc_o_reg ( .D(n17677), .SI(m5s8_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20917), .Q(m5s9_cyc), .QN(n18316) );
  SDFFARX1 m5_s14_cyc_o_reg ( .D(n17682), .SI(test_si31), .SE(test_se), .CLK(
        clk_i), .RSTB(n20918), .Q(m5s14_cyc), .QN(n18305) );
  SDFFARX1 m5_s12_cyc_o_reg ( .D(n17680), .SI(m5s11_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20918), .Q(m5s12_cyc), .QN(n18309) );
  SDFFARX1 m5_s10_cyc_o_reg ( .D(n17678), .SI(m5s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20917), .Q(m5s10_cyc), .QN(n18313) );
  SDFFARX1 m5_s8_cyc_o_reg ( .D(n17676), .SI(test_si30), .SE(test_se), .CLK(
        clk_i), .RSTB(n20917), .Q(m5s8_cyc), .QN(n18317) );
  SDFFARX1 m5_s5_cyc_o_reg ( .D(n17673), .SI(m5s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20916), .Q(m5s5_cyc), .QN(n18306) );
  SDFFARX1 m5_s3_cyc_o_reg ( .D(n17671), .SI(m5s2_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20916), .Q(m5s3_cyc), .QN(n18310) );
  SDFFARX1 m5_s1_cyc_o_reg ( .D(n17669), .SI(m5s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20916), .Q(test_so28), .QN(n18314) );
  SDFFARX1 m5_s7_cyc_o_reg ( .D(n17675), .SI(m5s6_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20917), .Q(test_so29), .QN(n18303) );
  SDFFARX1 m5_s4_cyc_o_reg ( .D(n17672), .SI(m5s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20916), .Q(m5s4_cyc), .QN(n18307) );
  SDFFARX1 m5_s2_cyc_o_reg ( .D(n17670), .SI(test_si29), .SE(test_se), .CLK(
        clk_i), .RSTB(n20916), .Q(m5s2_cyc), .QN(n18311) );
  SDFFARX1 m5_s0_cyc_o_reg ( .D(n17668), .SI(m4s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20915), .Q(m5s0_cyc), .QN(n18315) );
  SDFFARX1 m5_s15_cyc_o_reg ( .D(n17683), .SI(m5s14_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20918), .Q(m5s15_cyc), .QN(n18302) );
  SDFFARX1 m4_s13_cyc_o_reg ( .D(n17697), .SI(m4s12_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20921), .Q(m4s13_cyc), .QN() );
  SDFFARX1 m4_s12_cyc_o_reg ( .D(n17696), .SI(test_si28), .SE(test_se), .CLK(
        clk_i), .RSTB(n20921), .Q(m4s12_cyc), .QN() );
  SDFFARX1 m4_s11_cyc_o_reg ( .D(n17695), .SI(m4s10_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20921), .Q(test_so27), .QN() );
  SDFFARX1 m4_s10_cyc_o_reg ( .D(n17694), .SI(m4s9_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20921), .Q(m4s10_cyc), .QN() );
  SDFFARX1 m4_s8_cyc_o_reg ( .D(n17692), .SI(m4s7_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20920), .Q(m4s8_cyc), .QN() );
  SDFFARX1 m4_s5_cyc_o_reg ( .D(n17689), .SI(m4s4_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20920), .Q(test_so26), .QN() );
  SDFFARX1 m4_s4_cyc_o_reg ( .D(n17688), .SI(m4s3_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20919), .Q(m4s4_cyc), .QN() );
  SDFFARX1 m4_s1_cyc_o_reg ( .D(n17685), .SI(m4s0_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20919), .Q(m4s1_cyc), .QN() );
  SDFFARX1 m4_s0_cyc_o_reg ( .D(n17684), .SI(m3s15_cyc), .SE(test_se), .CLK(
        clk_i), .RSTB(n20919), .Q(m4s0_cyc), .QN() );
  INVX0 U18428 ( .IN(n18260), .QN(n13358) );
  INVX0 U18429 ( .IN(n18259), .QN(n11192) );
  INVX0 U18430 ( .IN(n18258), .QN(n12122) );
  INVX0 U18431 ( .IN(n18261), .QN(n9644) );
  INVX0 U18432 ( .IN(n13830), .QN(n3321) );
  INVX0 U18433 ( .IN(n13767), .QN(n3319) );
  LSDNENX1 U18434 ( .D(n18247), .ENB(n18333), .Q(n13670) );
  INVX0 U18435 ( .IN(n13704), .QN(n3317) );
  LSDNENX1 U18436 ( .D(n13358), .ENB(n18332), .Q(n13325) );
  INVX0 U18437 ( .IN(n13521), .QN(n3329) );
  INVX0 U18438 ( .IN(n13458), .QN(n3327) );
  INVX0 U18439 ( .IN(n13395), .QN(n3325) );
  LSDNENX1 U18440 ( .D(n11192), .ENB(n18331), .Q(n11159) );
  INVX0 U18441 ( .IN(n11355), .QN(n3265) );
  INVX0 U18442 ( .IN(n11292), .QN(n3263) );
  INVX0 U18443 ( .IN(n11229), .QN(n3261) );
  INVX0 U18444 ( .IN(n13212), .QN(n3337) );
  INVX0 U18445 ( .IN(n13149), .QN(n3335) );
  LSDNENX1 U18446 ( .D(n18256), .ENB(n18330), .Q(n13052) );
  INVX0 U18447 ( .IN(n13086), .QN(n3333) );
  INVX0 U18448 ( .IN(n12903), .QN(n3345) );
  INVX0 U18449 ( .IN(n12840), .QN(n3343) );
  LSDNENX1 U18450 ( .D(n18252), .ENB(n18329), .Q(n12743) );
  INVX0 U18451 ( .IN(n12777), .QN(n3341) );
  INVX0 U18452 ( .IN(n11046), .QN(n3273) );
  INVX0 U18453 ( .IN(n10983), .QN(n3271) );
  LSDNENX1 U18454 ( .D(n18255), .ENB(n18328), .Q(n10886) );
  INVX0 U18455 ( .IN(n10920), .QN(n3269) );
  INVX0 U18456 ( .IN(n10736), .QN(n3281) );
  INVX0 U18457 ( .IN(n10673), .QN(n3279) );
  LSDNENX1 U18458 ( .D(n18264), .ENB(m4s12_cyc), .Q(n10690) );
  LSDNENX1 U18459 ( .D(n18251), .ENB(n18327), .Q(n10576) );
  INVX0 U18460 ( .IN(n10610), .QN(n3277) );
  INVX0 U18461 ( .IN(n12594), .QN(n3353) );
  INVX0 U18462 ( .IN(n12531), .QN(n3351) );
  LSDNENX1 U18463 ( .D(n18248), .ENB(n18326), .Q(n12434) );
  INVX0 U18464 ( .IN(n12468), .QN(n3349) );
  LSDNENX1 U18465 ( .D(n12122), .ENB(n18325), .Q(n12089) );
  INVX0 U18466 ( .IN(n12285), .QN(n3361) );
  INVX0 U18467 ( .IN(n12222), .QN(n3359) );
  INVX0 U18468 ( .IN(n12159), .QN(n3357) );
  INVX0 U18469 ( .IN(n10427), .QN(n3289) );
  INVX0 U18470 ( .IN(n10364), .QN(n3287) );
  LSDNENX1 U18471 ( .D(n18254), .ENB(n18324), .Q(n10267) );
  INVX0 U18472 ( .IN(n10301), .QN(n3285) );
  INVX0 U18473 ( .IN(n10117), .QN(n3297) );
  INVX0 U18474 ( .IN(n10054), .QN(n3295) );
  LSDNENX1 U18475 ( .D(n18263), .ENB(m4s10_cyc), .Q(n10071) );
  LSDNENX1 U18476 ( .D(n18250), .ENB(n18323), .Q(n9957) );
  INVX0 U18477 ( .IN(n9991), .QN(n3293) );
  INVX0 U18478 ( .IN(n11975), .QN(n3369) );
  INVX0 U18479 ( .IN(n11912), .QN(n3367) );
  LSDNENX1 U18480 ( .D(n18253), .ENB(n18322), .Q(n11815) );
  INVX0 U18481 ( .IN(n11849), .QN(n3365) );
  INVX0 U18482 ( .IN(n11665), .QN(n3377) );
  INVX0 U18483 ( .IN(n11602), .QN(n3375) );
  LSDNENX1 U18484 ( .D(n18262), .ENB(m4s0_cyc), .Q(n11619) );
  LSDNENX1 U18485 ( .D(n18249), .ENB(n18321), .Q(n11505) );
  INVX0 U18486 ( .IN(n11539), .QN(n3373) );
  LSDNENX1 U18487 ( .D(n9644), .ENB(n18320), .Q(n9611) );
  INVX0 U18488 ( .IN(n9807), .QN(n3305) );
  INVX0 U18489 ( .IN(n9744), .QN(n3303) );
  INVX0 U18490 ( .IN(n9681), .QN(n3301) );
  INVX0 U18491 ( .IN(n9496), .QN(n3313) );
  INVX0 U18492 ( .IN(n9433), .QN(n3311) );
  LSDNENX1 U18493 ( .D(n18257), .ENB(n18319), .Q(n9336) );
  INVX0 U18494 ( .IN(n9370), .QN(n3309) );
  INVX0 U18495 ( .IN(n14031), .QN(n3253) );
  AND2X1 U18496 ( .IN1(n13851), .IN2(n13852), .Q(n13831) );
  NAND2X0 U18497 ( .IN1(n13634), .IN2(n18221), .QN(n13852) );
  INVX0 U18498 ( .IN(n13804), .QN(n2973) );
  AND2X1 U18499 ( .IN1(n13721), .IN2(n13722), .Q(n13705) );
  NAND2X0 U18500 ( .IN1(n13670), .IN2(n18222), .QN(n13722) );
  INVX0 U18501 ( .IN(n13679), .QN(n2965) );
  INVX0 U18502 ( .IN(n13495), .QN(n2989) );
  AND2X1 U18503 ( .IN1(n13412), .IN2(n13413), .Q(n13396) );
  NAND2X0 U18504 ( .IN1(n13361), .IN2(n18226), .QN(n13413) );
  INVX0 U18505 ( .IN(n13370), .QN(n2981) );
  INVX0 U18506 ( .IN(n11329), .QN(n2861) );
  AND2X1 U18507 ( .IN1(n11246), .IN2(n11247), .Q(n11230) );
  NAND2X0 U18508 ( .IN1(n11195), .IN2(n18225), .QN(n11247) );
  INVX0 U18509 ( .IN(n11204), .QN(n2853) );
  NAND2X0 U18510 ( .IN1(n13016), .IN2(n18239), .QN(n13234) );
  INVX0 U18511 ( .IN(n13186), .QN(n3005) );
  NAND2X0 U18512 ( .IN1(n13052), .IN2(n18242), .QN(n13104) );
  INVX0 U18513 ( .IN(n13061), .QN(n2997) );
  NAND2X0 U18514 ( .IN1(n12707), .IN2(n18234), .QN(n12925) );
  INVX0 U18515 ( .IN(n12877), .QN(n3021) );
  NAND2X0 U18516 ( .IN1(n12743), .IN2(n18246), .QN(n12795) );
  INVX0 U18517 ( .IN(n12752), .QN(n3013) );
  NAND2X0 U18518 ( .IN1(n10850), .IN2(n18240), .QN(n11068) );
  INVX0 U18519 ( .IN(n11020), .QN(n2877) );
  NAND2X0 U18520 ( .IN1(n10886), .IN2(n18243), .QN(n10938) );
  INVX0 U18521 ( .IN(n10895), .QN(n2869) );
  NAND2X0 U18522 ( .IN1(n10540), .IN2(n18231), .QN(n10758) );
  INVX0 U18523 ( .IN(n10710), .QN(n2893) );
  NAND2X0 U18524 ( .IN1(n10576), .IN2(n18235), .QN(n10628) );
  INVX0 U18525 ( .IN(n10585), .QN(n2885) );
  AND2X1 U18526 ( .IN1(n12615), .IN2(n12616), .Q(n12595) );
  NAND2X0 U18527 ( .IN1(n12398), .IN2(n18223), .QN(n12616) );
  INVX0 U18528 ( .IN(n12568), .QN(n3037) );
  AND2X1 U18529 ( .IN1(n12485), .IN2(n12486), .Q(n12469) );
  NAND2X0 U18530 ( .IN1(n12434), .IN2(n18228), .QN(n12486) );
  INVX0 U18531 ( .IN(n12443), .QN(n3029) );
  INVX0 U18532 ( .IN(n12259), .QN(n3053) );
  AND2X1 U18533 ( .IN1(n12176), .IN2(n12177), .Q(n12160) );
  NAND2X0 U18534 ( .IN1(n12125), .IN2(n18224), .QN(n12177) );
  INVX0 U18535 ( .IN(n12134), .QN(n3045) );
  NAND2X0 U18536 ( .IN1(n10231), .IN2(n18229), .QN(n10449) );
  INVX0 U18537 ( .IN(n10401), .QN(n2909) );
  NAND2X0 U18538 ( .IN1(n10267), .IN2(n18244), .QN(n10319) );
  INVX0 U18539 ( .IN(n10276), .QN(n2901) );
  NAND2X0 U18540 ( .IN1(n9921), .IN2(n18232), .QN(n10139) );
  INVX0 U18541 ( .IN(n10091), .QN(n2925) );
  NAND2X0 U18542 ( .IN1(n9957), .IN2(n18236), .QN(n10009) );
  INVX0 U18543 ( .IN(n9966), .QN(n2917) );
  NAND2X0 U18544 ( .IN1(n11779), .IN2(n18230), .QN(n11997) );
  INVX0 U18545 ( .IN(n11949), .QN(n3069) );
  NAND2X0 U18546 ( .IN1(n11815), .IN2(n18245), .QN(n11867) );
  INVX0 U18547 ( .IN(n11824), .QN(n3061) );
  NAND2X0 U18548 ( .IN1(n11469), .IN2(n18233), .QN(n11687) );
  INVX0 U18549 ( .IN(n11639), .QN(n3085) );
  NAND2X0 U18550 ( .IN1(n11505), .IN2(n18237), .QN(n11557) );
  INVX0 U18551 ( .IN(n11514), .QN(n3077) );
  INVX0 U18552 ( .IN(n9781), .QN(n2941) );
  AND2X1 U18553 ( .IN1(n9698), .IN2(n9699), .Q(n9682) );
  NAND2X0 U18554 ( .IN1(n9647), .IN2(n18227), .QN(n9699) );
  INVX0 U18555 ( .IN(n9656), .QN(n2933) );
  NAND2X0 U18556 ( .IN1(n9300), .IN2(n18238), .QN(n9518) );
  INVX0 U18557 ( .IN(n9470), .QN(n2957) );
  NAND2X0 U18558 ( .IN1(n9336), .IN2(n18241), .QN(n9388) );
  INVX0 U18559 ( .IN(n9345), .QN(n2949) );
  AND4X1 U18560 ( .IN1(s15_addr_o[25]), .IN2(s15_addr_o[26]), .IN3(
        s15_addr_o[24]), .IN4(n17086), .Q(n17780) );
  AND2X1 U18561 ( .IN1(n14822), .IN2(n14831), .Q(n17781) );
  AND2X1 U18562 ( .IN1(n15475), .IN2(n15478), .Q(n17782) );
  AND2X1 U18563 ( .IN1(n16085), .IN2(n16088), .Q(n17783) );
  AND2X1 U18564 ( .IN1(n16695), .IN2(n16698), .Q(n17784) );
  AND2X1 U18565 ( .IN1(n15170), .IN2(n15173), .Q(n17785) );
  AND2X1 U18566 ( .IN1(n16390), .IN2(n16393), .Q(n17786) );
  AND2X1 U18567 ( .IN1(n17007), .IN2(n17024), .Q(n17787) );
  AND2X1 U18568 ( .IN1(n15780), .IN2(n15783), .Q(n17788) );
  AND2X1 U18569 ( .IN1(n15781), .IN2(n15780), .Q(n17789) );
  AND3X1 U18570 ( .IN1(n3985), .IN2(n14870), .IN3(n3980), .Q(n17790) );
  AND3X1 U18571 ( .IN1(n3580), .IN2(n14860), .IN3(n3575), .Q(n17791) );
  AND3X1 U18572 ( .IN1(n3535), .IN2(n14873), .IN3(n3530), .Q(n17792) );
  AND2X1 U18573 ( .IN1(n14847), .IN2(n14826), .Q(n17793) );
  AND2X1 U18574 ( .IN1(n14847), .IN2(n14821), .Q(n17794) );
  AND2X1 U18575 ( .IN1(n14840), .IN2(n14826), .Q(n17795) );
  AND2X1 U18576 ( .IN1(n14840), .IN2(n14821), .Q(n17796) );
  AND2X1 U18577 ( .IN1(n15482), .IN2(n15476), .Q(n17797) );
  AND2X1 U18578 ( .IN1(n15482), .IN2(n15474), .Q(n17798) );
  AND2X1 U18579 ( .IN1(n15481), .IN2(n15476), .Q(n17799) );
  AND2X1 U18580 ( .IN1(n15481), .IN2(n15474), .Q(n17800) );
  AND2X1 U18581 ( .IN1(n16092), .IN2(n16086), .Q(n17801) );
  AND2X1 U18582 ( .IN1(n16092), .IN2(n16084), .Q(n17802) );
  AND2X1 U18583 ( .IN1(n16091), .IN2(n16086), .Q(n17803) );
  AND2X1 U18584 ( .IN1(n16091), .IN2(n16084), .Q(n17804) );
  AND2X1 U18585 ( .IN1(n16702), .IN2(n16696), .Q(n17805) );
  AND2X1 U18586 ( .IN1(n16702), .IN2(n16694), .Q(n17806) );
  AND2X1 U18587 ( .IN1(n16701), .IN2(n16696), .Q(n17807) );
  AND2X1 U18588 ( .IN1(n16701), .IN2(n16694), .Q(n17808) );
  AND2X1 U18589 ( .IN1(n14840), .IN2(n14835), .Q(n17809) );
  AND2X1 U18590 ( .IN1(n14840), .IN2(n14831), .Q(n17810) );
  AND2X1 U18591 ( .IN1(n15481), .IN2(n15479), .Q(n17811) );
  AND2X1 U18592 ( .IN1(n15481), .IN2(n15478), .Q(n17812) );
  AND2X1 U18593 ( .IN1(n16091), .IN2(n16089), .Q(n17813) );
  AND2X1 U18594 ( .IN1(n16091), .IN2(n16088), .Q(n17814) );
  AND2X1 U18595 ( .IN1(n16701), .IN2(n16699), .Q(n17815) );
  AND2X1 U18596 ( .IN1(n16701), .IN2(n16698), .Q(n17816) );
  AND2X1 U18597 ( .IN1(n14822), .IN2(n14835), .Q(n17817) );
  AND2X1 U18598 ( .IN1(n16085), .IN2(n16089), .Q(n17818) );
  AND2X1 U18599 ( .IN1(n16695), .IN2(n16699), .Q(n17819) );
  AND2X1 U18600 ( .IN1(n14847), .IN2(n14831), .Q(n17820) );
  AND2X1 U18601 ( .IN1(n15482), .IN2(n15478), .Q(n17821) );
  AND2X1 U18602 ( .IN1(n16092), .IN2(n16088), .Q(n17822) );
  AND2X1 U18603 ( .IN1(n16702), .IN2(n16698), .Q(n17823) );
  AND2X1 U18604 ( .IN1(n14826), .IN2(n14830), .Q(n17824) );
  AND2X1 U18605 ( .IN1(n16086), .IN2(n16087), .Q(n17825) );
  AND2X1 U18606 ( .IN1(n16696), .IN2(n16697), .Q(n17826) );
  AND2X1 U18607 ( .IN1(n15475), .IN2(n15479), .Q(n17827) );
  AND2X1 U18608 ( .IN1(n15476), .IN2(n15475), .Q(n17828) );
  AND2X1 U18609 ( .IN1(n15476), .IN2(n15477), .Q(n17829) );
  AND2X1 U18610 ( .IN1(n14835), .IN2(n14830), .Q(n17830) );
  AND2X1 U18611 ( .IN1(n15479), .IN2(n15477), .Q(n17831) );
  AND2X1 U18612 ( .IN1(n16089), .IN2(n16087), .Q(n17832) );
  AND2X1 U18613 ( .IN1(n16699), .IN2(n16697), .Q(n17833) );
  AND2X1 U18614 ( .IN1(n15177), .IN2(n15169), .Q(n17834) );
  AND2X1 U18615 ( .IN1(n15176), .IN2(n15171), .Q(n17835) );
  AND2X1 U18616 ( .IN1(n15176), .IN2(n15169), .Q(n17836) );
  AND2X1 U18617 ( .IN1(n15787), .IN2(n15779), .Q(n17837) );
  AND2X1 U18618 ( .IN1(n15786), .IN2(n15781), .Q(n17838) );
  AND2X1 U18619 ( .IN1(n15786), .IN2(n15779), .Q(n17839) );
  AND2X1 U18620 ( .IN1(n16397), .IN2(n16389), .Q(n17840) );
  AND2X1 U18621 ( .IN1(n16396), .IN2(n16391), .Q(n17841) );
  AND2X1 U18622 ( .IN1(n16396), .IN2(n16389), .Q(n17842) );
  AND2X1 U18623 ( .IN1(n17056), .IN2(n17006), .Q(n17843) );
  AND2X1 U18624 ( .IN1(n17041), .IN2(n17015), .Q(n17844) );
  AND2X1 U18625 ( .IN1(n17041), .IN2(n17006), .Q(n17845) );
  AND2X1 U18626 ( .IN1(n15176), .IN2(n15173), .Q(n17846) );
  AND2X1 U18627 ( .IN1(n15786), .IN2(n15783), .Q(n17847) );
  AND2X1 U18628 ( .IN1(n16396), .IN2(n16393), .Q(n17848) );
  AND2X1 U18629 ( .IN1(n17041), .IN2(n17024), .Q(n17849) );
  AND2X1 U18630 ( .IN1(n15177), .IN2(n15173), .Q(n17850) );
  AND2X1 U18631 ( .IN1(n15787), .IN2(n15783), .Q(n17851) );
  AND2X1 U18632 ( .IN1(n16397), .IN2(n16393), .Q(n17852) );
  AND2X1 U18633 ( .IN1(n17056), .IN2(n17024), .Q(n17853) );
  AND2X1 U18634 ( .IN1(n15170), .IN2(n15174), .Q(n17854) );
  AND2X1 U18635 ( .IN1(n15780), .IN2(n15784), .Q(n17855) );
  AND2X1 U18636 ( .IN1(n16390), .IN2(n16394), .Q(n17856) );
  AND2X1 U18637 ( .IN1(n17007), .IN2(n17032), .Q(n17857) );
  AND2X1 U18638 ( .IN1(n15171), .IN2(n15170), .Q(n17858) );
  AND2X1 U18639 ( .IN1(n15171), .IN2(n15172), .Q(n17859) );
  AND2X1 U18640 ( .IN1(n15781), .IN2(n15782), .Q(n17860) );
  AND2X1 U18641 ( .IN1(n16391), .IN2(n16390), .Q(n17861) );
  AND2X1 U18642 ( .IN1(n16391), .IN2(n16392), .Q(n17862) );
  AND2X1 U18643 ( .IN1(n17015), .IN2(n17007), .Q(n17863) );
  AND2X1 U18644 ( .IN1(n17015), .IN2(n17023), .Q(n17864) );
  AND2X1 U18645 ( .IN1(n15174), .IN2(n15172), .Q(n17865) );
  AND2X1 U18646 ( .IN1(n15784), .IN2(n15782), .Q(n17866) );
  AND2X1 U18647 ( .IN1(n16394), .IN2(n16392), .Q(n17867) );
  AND2X1 U18648 ( .IN1(n17032), .IN2(n17023), .Q(n17868) );
  AND2X1 U18649 ( .IN1(n14821), .IN2(n14822), .Q(n17869) );
  AND2X1 U18650 ( .IN1(n16084), .IN2(n16085), .Q(n17870) );
  AND2X1 U18651 ( .IN1(n16694), .IN2(n16695), .Q(n17871) );
  AND2X1 U18652 ( .IN1(n15474), .IN2(n15475), .Q(n17872) );
  AND2X1 U18653 ( .IN1(n14830), .IN2(n14831), .Q(n17873) );
  AND2X1 U18654 ( .IN1(n15477), .IN2(n15478), .Q(n17874) );
  AND2X1 U18655 ( .IN1(n16087), .IN2(n16088), .Q(n17875) );
  AND2X1 U18656 ( .IN1(n16697), .IN2(n16698), .Q(n17876) );
  AND2X1 U18657 ( .IN1(n15172), .IN2(n15173), .Q(n17877) );
  AND2X1 U18658 ( .IN1(n15782), .IN2(n15783), .Q(n17878) );
  AND2X1 U18659 ( .IN1(n16392), .IN2(n16393), .Q(n17879) );
  AND2X1 U18660 ( .IN1(n17023), .IN2(n17024), .Q(n17880) );
  AND3X1 U18661 ( .IN1(n3850), .IN2(n14824), .IN3(n3845), .Q(n17881) );
  AND2X1 U18662 ( .IN1(n14826), .IN2(n14822), .Q(n17882) );
  AND2X1 U18663 ( .IN1(n16086), .IN2(n16085), .Q(n17883) );
  AND2X1 U18664 ( .IN1(n16696), .IN2(n16695), .Q(n17884) );
  AND3X1 U18665 ( .IN1(n4160), .IN2(n4165), .IN3(n4166), .Q(n17885) );
  AND3X1 U18666 ( .IN1(n4115), .IN2(n4120), .IN3(n4121), .Q(n17886) );
  AND3X1 U18667 ( .IN1(n4070), .IN2(n4075), .IN3(n4076), .Q(n17887) );
  AND3X1 U18668 ( .IN1(n4025), .IN2(n4030), .IN3(n4031), .Q(n17888) );
  AND3X1 U18669 ( .IN1(n3980), .IN2(n3985), .IN3(n3986), .Q(n17889) );
  AND3X1 U18670 ( .IN1(n3890), .IN2(n3895), .IN3(n3896), .Q(n17890) );
  AND3X1 U18671 ( .IN1(n3845), .IN2(n3850), .IN3(n3851), .Q(n17891) );
  AND3X1 U18672 ( .IN1(n3800), .IN2(n3805), .IN3(n3806), .Q(n17892) );
  AND3X1 U18673 ( .IN1(n3755), .IN2(n3760), .IN3(n3761), .Q(n17893) );
  AND3X1 U18674 ( .IN1(n3710), .IN2(n3715), .IN3(n3716), .Q(n17894) );
  AND3X1 U18675 ( .IN1(n3665), .IN2(n3670), .IN3(n3671), .Q(n17895) );
  AND3X1 U18676 ( .IN1(n3620), .IN2(n3625), .IN3(n3626), .Q(n17896) );
  AND3X1 U18677 ( .IN1(n3575), .IN2(n3580), .IN3(n3581), .Q(n17897) );
  AND3X1 U18678 ( .IN1(n3530), .IN2(n3535), .IN3(n3536), .Q(n17898) );
  AND3X1 U18679 ( .IN1(n4165), .IN2(n14856), .IN3(n4166), .Q(n17899) );
  AND3X1 U18680 ( .IN1(n4120), .IN2(n14853), .IN3(n4121), .Q(n17900) );
  AND3X1 U18681 ( .IN1(n4120), .IN2(n14854), .IN3(n4115), .Q(n17901) );
  AND3X1 U18682 ( .IN1(n4075), .IN2(n14866), .IN3(n4076), .Q(n17902) );
  AND3X1 U18683 ( .IN1(n4075), .IN2(n14867), .IN3(n4070), .Q(n17903) );
  AND3X1 U18684 ( .IN1(n4030), .IN2(n14863), .IN3(n4031), .Q(n17904) );
  AND3X1 U18685 ( .IN1(n4030), .IN2(n14864), .IN3(n4025), .Q(n17905) );
  AND3X1 U18686 ( .IN1(n3985), .IN2(n14869), .IN3(n3986), .Q(n17906) );
  AND3X1 U18687 ( .IN1(n3895), .IN2(n14833), .IN3(n3890), .Q(n17907) );
  AND3X1 U18688 ( .IN1(n3895), .IN2(n14832), .IN3(n3896), .Q(n17908) );
  AND3X1 U18689 ( .IN1(n3850), .IN2(n14823), .IN3(n3851), .Q(n17909) );
  AND3X1 U18690 ( .IN1(n3805), .IN2(n14818), .IN3(n3806), .Q(n17910) );
  AND3X1 U18691 ( .IN1(n3760), .IN2(n14841), .IN3(n3761), .Q(n17911) );
  AND3X1 U18692 ( .IN1(n3760), .IN2(n14842), .IN3(n3755), .Q(n17912) );
  AND3X1 U18693 ( .IN1(n3715), .IN2(n14837), .IN3(n3716), .Q(n17913) );
  AND3X1 U18694 ( .IN1(n3715), .IN2(n14838), .IN3(n3710), .Q(n17914) );
  AND3X1 U18695 ( .IN1(n3670), .IN2(n14844), .IN3(n3671), .Q(n17915) );
  AND3X1 U18696 ( .IN1(n3625), .IN2(n14848), .IN3(n3626), .Q(n17916) );
  AND3X1 U18697 ( .IN1(n3580), .IN2(n14859), .IN3(n3581), .Q(n17917) );
  AND3X1 U18698 ( .IN1(n3535), .IN2(n14872), .IN3(n3536), .Q(n17918) );
  AND3X1 U18699 ( .IN1(n14869), .IN2(n14870), .IN3(n3985), .Q(n17919) );
  AND3X1 U18700 ( .IN1(n14832), .IN2(n14833), .IN3(n3895), .Q(n17920) );
  AND3X1 U18701 ( .IN1(n14844), .IN2(n14845), .IN3(n3670), .Q(n17921) );
  AND3X1 U18702 ( .IN1(n14848), .IN2(n14849), .IN3(n3625), .Q(n17922) );
  AND3X1 U18703 ( .IN1(n14859), .IN2(n14860), .IN3(n3580), .Q(n17923) );
  AND3X1 U18704 ( .IN1(n14872), .IN2(n14873), .IN3(n3535), .Q(n17924) );
  AND3X1 U18705 ( .IN1(n14856), .IN2(n14857), .IN3(n4165), .Q(n17925) );
  AND3X1 U18706 ( .IN1(n14853), .IN2(n14854), .IN3(n4120), .Q(n17926) );
  AND3X1 U18707 ( .IN1(n14866), .IN2(n14867), .IN3(n4075), .Q(n17927) );
  AND3X1 U18708 ( .IN1(n14863), .IN2(n14864), .IN3(n4030), .Q(n17928) );
  AND3X1 U18709 ( .IN1(n14823), .IN2(n14824), .IN3(n3850), .Q(n17929) );
  AND3X1 U18710 ( .IN1(n14818), .IN2(n14819), .IN3(n3805), .Q(n17930) );
  AND3X1 U18711 ( .IN1(n14841), .IN2(n14842), .IN3(n3760), .Q(n17931) );
  AND3X1 U18712 ( .IN1(n14837), .IN2(n14838), .IN3(n3715), .Q(n17932) );
  OR2X1 U18713 ( .IN1(n14282), .IN2(n18302), .Q(n18157) );
  OR2X1 U18714 ( .IN1(n14300), .IN2(n18302), .Q(n18158) );
  OR2X1 U18715 ( .IN1(n13355), .IN2(n18304), .Q(n18159) );
  OR2X1 U18716 ( .IN1(n11189), .IN2(n18305), .Q(n18160) );
  OR2X1 U18717 ( .IN1(n12119), .IN2(n18311), .Q(n18161) );
  OR2X1 U18718 ( .IN1(n9641), .IN2(n18316), .Q(n18162) );
  OR2X1 U18719 ( .IN1(n13664), .IN2(n18303), .Q(n18163) );
  OR2X1 U18720 ( .IN1(n13665), .IN2(n18303), .Q(n18164) );
  OR2X1 U18721 ( .IN1(n13356), .IN2(n18304), .Q(n18165) );
  OR2X1 U18722 ( .IN1(n11190), .IN2(n18305), .Q(n18166) );
  OR2X1 U18723 ( .IN1(n13046), .IN2(n18306), .Q(n18167) );
  OR2X1 U18724 ( .IN1(n13047), .IN2(n18306), .Q(n18168) );
  OR2X1 U18725 ( .IN1(n12737), .IN2(n18307), .Q(n18169) );
  OR2X1 U18726 ( .IN1(n12738), .IN2(n18307), .Q(n18170) );
  OR2X1 U18727 ( .IN1(n10880), .IN2(n18308), .Q(n18171) );
  OR2X1 U18728 ( .IN1(n10881), .IN2(n18308), .Q(n18172) );
  OR2X1 U18729 ( .IN1(n10570), .IN2(n18309), .Q(n18173) );
  OR2X1 U18730 ( .IN1(n10571), .IN2(n18309), .Q(n18174) );
  OR2X1 U18731 ( .IN1(n12428), .IN2(n18310), .Q(n18175) );
  OR2X1 U18732 ( .IN1(n12429), .IN2(n18310), .Q(n18176) );
  OR2X1 U18733 ( .IN1(n12120), .IN2(n18311), .Q(n18177) );
  OR2X1 U18734 ( .IN1(n10261), .IN2(n18312), .Q(n18178) );
  OR2X1 U18735 ( .IN1(n10262), .IN2(n18312), .Q(n18179) );
  OR2X1 U18736 ( .IN1(n9951), .IN2(n18313), .Q(n18180) );
  OR2X1 U18737 ( .IN1(n9952), .IN2(n18313), .Q(n18181) );
  OR2X1 U18738 ( .IN1(n11809), .IN2(n18314), .Q(n18182) );
  OR2X1 U18739 ( .IN1(n11810), .IN2(n18314), .Q(n18183) );
  OR2X1 U18740 ( .IN1(n11499), .IN2(n18315), .Q(n18184) );
  OR2X1 U18741 ( .IN1(n11500), .IN2(n18315), .Q(n18185) );
  OR2X1 U18742 ( .IN1(n9642), .IN2(n18316), .Q(n18186) );
  OR2X1 U18743 ( .IN1(n9330), .IN2(n18317), .Q(n18187) );
  OR2X1 U18744 ( .IN1(n9331), .IN2(n18317), .Q(n18188) );
  AND2X1 U18745 ( .IN1(n18163), .IN2(n3863), .Q(n18221) );
  AND2X1 U18746 ( .IN1(n18164), .IN2(n3871), .Q(n18222) );
  AND2X1 U18747 ( .IN1(n18175), .IN2(n3683), .Q(n18223) );
  AND2X1 U18748 ( .IN1(n18177), .IN2(n3646), .Q(n18224) );
  AND2X1 U18749 ( .IN1(n18166), .IN2(n4186), .Q(n18225) );
  AND2X1 U18750 ( .IN1(n18165), .IN2(n3826), .Q(n18226) );
  AND2X1 U18751 ( .IN1(n18186), .IN2(n3961), .Q(n18227) );
  AND2X1 U18752 ( .IN1(n18176), .IN2(n3691), .Q(n18228) );
  AND2X1 U18753 ( .IN1(n18178), .IN2(n4043), .Q(n18229) );
  AND2X1 U18754 ( .IN1(n18182), .IN2(n3593), .Q(n18230) );
  AND2X1 U18755 ( .IN1(n18173), .IN2(n4088), .Q(n18231) );
  AND2X1 U18756 ( .IN1(n18180), .IN2(n3998), .Q(n18232) );
  AND2X1 U18757 ( .IN1(n18184), .IN2(n3548), .Q(n18233) );
  AND2X1 U18758 ( .IN1(n18169), .IN2(n3728), .Q(n18234) );
  AND2X1 U18759 ( .IN1(n18174), .IN2(n4096), .Q(n18235) );
  AND2X1 U18760 ( .IN1(n18181), .IN2(n4006), .Q(n18236) );
  AND2X1 U18761 ( .IN1(n18185), .IN2(n3556), .Q(n18237) );
  AND2X1 U18762 ( .IN1(n18187), .IN2(n3908), .Q(n18238) );
  AND2X1 U18763 ( .IN1(n18167), .IN2(n3773), .Q(n18239) );
  AND2X1 U18764 ( .IN1(n18171), .IN2(n4133), .Q(n18240) );
  AND2X1 U18765 ( .IN1(n18188), .IN2(n3916), .Q(n18241) );
  AND2X1 U18766 ( .IN1(n18168), .IN2(n3781), .Q(n18242) );
  AND2X1 U18767 ( .IN1(n18172), .IN2(n4141), .Q(n18243) );
  AND2X1 U18768 ( .IN1(n18179), .IN2(n4051), .Q(n18244) );
  AND2X1 U18769 ( .IN1(n18183), .IN2(n3601), .Q(n18245) );
  AND2X1 U18770 ( .IN1(n18170), .IN2(n3736), .Q(n18246) );
  LSDNENX1 U18771 ( .D(n13667), .ENB(n18333), .Q(n13634) );
  NAND2X1 U18772 ( .IN1(conf7_8_), .IN2(n17964), .QN(n13667) );
  NBUFFX2 U18773 ( .IN(n13668), .Q(n18247) );
  LSDNENX1 U18774 ( .D(n12431), .ENB(n18326), .Q(n12398) );
  NAND2X1 U18775 ( .IN1(conf3_8_), .IN2(n17945), .QN(n12431) );
  LSDNENX1 U18776 ( .D(n12123), .ENB(n18325), .Q(n12125) );
  NAND2X1 U18777 ( .IN1(conf2_9_), .IN2(n17946), .QN(n12123) );
  LSDNENX1 U18778 ( .D(n11193), .ENB(n18331), .Q(n11195) );
  NAND2X1 U18779 ( .IN1(conf14_9_), .IN2(n17948), .QN(n11193) );
  LSDNENX1 U18780 ( .D(n13359), .ENB(n18332), .Q(n13361) );
  NAND2X1 U18781 ( .IN1(conf6_9_), .IN2(n17947), .QN(n13359) );
  LSDNENX1 U18782 ( .D(n9645), .ENB(n18320), .Q(n9647) );
  NAND2X1 U18783 ( .IN1(conf9_9_), .IN2(n17940), .QN(n9645) );
  NBUFFX2 U18784 ( .IN(n12432), .Q(n18248) );
  LSDNENX1 U18785 ( .D(n11502), .ENB(n18321), .Q(n11469) );
  NAND2X1 U18786 ( .IN1(conf0_8_), .IN2(n17959), .QN(n11502) );
  LSDNENX1 U18787 ( .D(n9954), .ENB(n18323), .Q(n9921) );
  NAND2X1 U18788 ( .IN1(conf10_8_), .IN2(n17957), .QN(n9954) );
  LSDNENX1 U18789 ( .D(n10573), .ENB(n18327), .Q(n10540) );
  NAND2X1 U18790 ( .IN1(conf12_8_), .IN2(n17958), .QN(n10573) );
  LSDNENX1 U18791 ( .D(n12740), .ENB(n18329), .Q(n12707) );
  NAND2X1 U18792 ( .IN1(conf4_8_), .IN2(n17934), .QN(n12740) );
  LSDNENX1 U18793 ( .D(n11812), .ENB(n18322), .Q(n11779) );
  NAND2X1 U18794 ( .IN1(conf1_8_), .IN2(n18064), .QN(n11812) );
  LSDNENX1 U18795 ( .D(n10264), .ENB(n18324), .Q(n10231) );
  NAND2X1 U18796 ( .IN1(conf11_8_), .IN2(n18061), .QN(n10264) );
  LSDNENX1 U18797 ( .D(n10883), .ENB(n18328), .Q(n10850) );
  NAND2X1 U18798 ( .IN1(conf13_8_), .IN2(n18062), .QN(n10883) );
  LSDNENX1 U18799 ( .D(n13049), .ENB(n18330), .Q(n13016) );
  NAND2X1 U18800 ( .IN1(conf5_8_), .IN2(n18063), .QN(n13049) );
  LSDNENX1 U18801 ( .D(n9333), .ENB(n18319), .Q(n9300) );
  NAND2X1 U18802 ( .IN1(conf8_8_), .IN2(n17933), .QN(n9333) );
  NBUFFX2 U18803 ( .IN(n11503), .Q(n18249) );
  NBUFFX2 U18804 ( .IN(n9955), .Q(n18250) );
  NBUFFX2 U18805 ( .IN(n10574), .Q(n18251) );
  NBUFFX2 U18806 ( .IN(n12741), .Q(n18252) );
  NBUFFX2 U18807 ( .IN(n11813), .Q(n18253) );
  NBUFFX2 U18808 ( .IN(n10265), .Q(n18254) );
  NBUFFX2 U18809 ( .IN(n10884), .Q(n18255) );
  NBUFFX2 U18810 ( .IN(n13050), .Q(n18256) );
  NBUFFX2 U18811 ( .IN(n9334), .Q(n18257) );
  ISOLANDX1 U18812 ( .D(conf2_8_), .ISO(conf2_9_), .Q(n18258) );
  ISOLANDX1 U18813 ( .D(conf14_8_), .ISO(conf14_9_), .Q(n18259) );
  ISOLANDX1 U18814 ( .D(conf6_8_), .ISO(conf6_9_), .Q(n18260) );
  ISOLANDX1 U18815 ( .D(conf9_8_), .ISO(conf9_9_), .Q(n18261) );
  AND2X1 U18816 ( .IN1(n10448), .IN2(n10449), .Q(n10428) );
  AND2X1 U18817 ( .IN1(n11996), .IN2(n11997), .Q(n11976) );
  AND2X1 U18818 ( .IN1(n10757), .IN2(n10758), .Q(n10737) );
  AND2X1 U18819 ( .IN1(n10138), .IN2(n10139), .Q(n10118) );
  AND2X1 U18820 ( .IN1(n11686), .IN2(n11687), .Q(n11666) );
  AND2X1 U18821 ( .IN1(n12924), .IN2(n12925), .Q(n12904) );
  AND2X1 U18822 ( .IN1(n10627), .IN2(n10628), .Q(n10611) );
  AND2X1 U18823 ( .IN1(n10008), .IN2(n10009), .Q(n9992) );
  AND2X1 U18824 ( .IN1(n11556), .IN2(n11557), .Q(n11540) );
  AND2X1 U18825 ( .IN1(n9517), .IN2(n9518), .Q(n9497) );
  AND2X1 U18826 ( .IN1(n13233), .IN2(n13234), .Q(n13213) );
  AND2X1 U18827 ( .IN1(n11067), .IN2(n11068), .Q(n11047) );
  AND2X1 U18828 ( .IN1(n9387), .IN2(n9388), .Q(n9371) );
  AND2X1 U18829 ( .IN1(n13103), .IN2(n13104), .Q(n13087) );
  AND2X1 U18830 ( .IN1(n10937), .IN2(n10938), .Q(n10921) );
  AND2X1 U18831 ( .IN1(n10318), .IN2(n10319), .Q(n10302) );
  AND2X1 U18832 ( .IN1(n11866), .IN2(n11867), .Q(n11850) );
  AND2X1 U18833 ( .IN1(n12794), .IN2(n12795), .Q(n12778) );
  INVX0 U18834 ( .IN(n14001), .QN(n2837) );
  LSDNENX1 U18835 ( .D(n12118), .ENB(m5s2_cyc), .Q(n12235) );
  NAND2X1 U18836 ( .IN1(n18077), .IN2(n17943), .QN(n12118) );
  LSDNENX1 U18837 ( .D(n11188), .ENB(m5s14_cyc), .Q(n11305) );
  NAND2X1 U18838 ( .IN1(n18076), .IN2(n17942), .QN(n11188) );
  LSDNENX1 U18839 ( .D(n13354), .ENB(m5s6_cyc), .Q(n13471) );
  NAND2X1 U18840 ( .IN1(n18075), .IN2(n17941), .QN(n13354) );
  LSDNENX1 U18841 ( .D(n9640), .ENB(m5s9_cyc), .Q(n9757) );
  NAND2X1 U18842 ( .IN1(n17952), .IN2(n18068), .QN(n9640) );
  LSDNENX1 U18843 ( .D(n12427), .ENB(m5s3_cyc), .Q(n12544) );
  NAND2X1 U18844 ( .IN1(n17951), .IN2(n18067), .QN(n12427) );
  LSDNENX1 U18845 ( .D(n13663), .ENB(test_so29), .Q(n13780) );
  NAND2X1 U18846 ( .IN1(n17950), .IN2(n18069), .QN(n13663) );
  LSDNENX1 U18847 ( .D(n14071), .ENB(m5s15_cyc), .Q(n14044) );
  NAND2X1 U18848 ( .IN1(n17949), .IN2(n18070), .QN(n14071) );
  LSDNENX1 U18849 ( .D(n11498), .ENB(m5s0_cyc), .Q(n11615) );
  NAND2X1 U18850 ( .IN1(n18082), .IN2(n17956), .QN(n11498) );
  LSDNENX1 U18851 ( .D(n9950), .ENB(m5s10_cyc), .Q(n10067) );
  NAND2X1 U18852 ( .IN1(n18081), .IN2(n17955), .QN(n9950) );
  LSDNENX1 U18853 ( .D(n10569), .ENB(m5s12_cyc), .Q(n10686) );
  NAND2X1 U18854 ( .IN1(n18080), .IN2(n17954), .QN(n10569) );
  LSDNENX1 U18855 ( .D(n12736), .ENB(m5s4_cyc), .Q(n12853) );
  NAND2X1 U18856 ( .IN1(n18079), .IN2(n17953), .QN(n12736) );
  LSDNENX1 U18857 ( .D(n11808), .ENB(test_so28), .Q(n11925) );
  NAND2X1 U18858 ( .IN1(n17963), .IN2(n18074), .QN(n11808) );
  LSDNENX1 U18859 ( .D(n10260), .ENB(m5s11_cyc), .Q(n10377) );
  NAND2X1 U18860 ( .IN1(n17962), .IN2(n18073), .QN(n10260) );
  LSDNENX1 U18861 ( .D(n10879), .ENB(test_so30), .Q(n10996) );
  NAND2X1 U18862 ( .IN1(n17961), .IN2(n18072), .QN(n10879) );
  LSDNENX1 U18863 ( .D(n13045), .ENB(m5s5_cyc), .Q(n13162) );
  NAND2X1 U18864 ( .IN1(n17960), .IN2(n18071), .QN(n13045) );
  LSDNENX1 U18865 ( .D(n9329), .ENB(m5s8_cyc), .Q(n9446) );
  NAND2X1 U18866 ( .IN1(n18078), .IN2(n17944), .QN(n9329) );
  INVX0 U18867 ( .IN(n13250), .QN(n3009) );
  INVX0 U18868 ( .IN(n12941), .QN(n3025) );
  INVX0 U18869 ( .IN(n11084), .QN(n2881) );
  INVX0 U18870 ( .IN(n10774), .QN(n2897) );
  INVX0 U18871 ( .IN(n10465), .QN(n2913) );
  INVX0 U18872 ( .IN(n10155), .QN(n2929) );
  INVX0 U18873 ( .IN(n12013), .QN(n3073) );
  INVX0 U18874 ( .IN(n11703), .QN(n3089) );
  INVX0 U18875 ( .IN(n9534), .QN(n2961) );
  INVX0 U18876 ( .IN(n13280), .QN(n3340) );
  INVX0 U18877 ( .IN(n12971), .QN(n3348) );
  INVX0 U18878 ( .IN(n11114), .QN(n3276) );
  INVX0 U18879 ( .IN(n10804), .QN(n3284) );
  INVX0 U18880 ( .IN(n10495), .QN(n3292) );
  INVX0 U18881 ( .IN(n10185), .QN(n3300) );
  INVX0 U18882 ( .IN(n12043), .QN(n3372) );
  INVX0 U18883 ( .IN(n11733), .QN(n3380) );
  INVX0 U18884 ( .IN(n9564), .QN(n3316) );
  INVX0 U18885 ( .IN(n13295), .QN(n3392) );
  INVX0 U18886 ( .IN(n12986), .QN(n3393) );
  INVX0 U18887 ( .IN(n11129), .QN(n3384) );
  INVX0 U18888 ( .IN(n10819), .QN(n3385) );
  INVX0 U18889 ( .IN(n10510), .QN(n3386) );
  INVX0 U18890 ( .IN(n10200), .QN(n3387) );
  INVX0 U18891 ( .IN(n12058), .QN(n3396) );
  INVX0 U18892 ( .IN(n11748), .QN(n3397) );
  INVX0 U18893 ( .IN(n9579), .QN(n3389) );
  LSDNENX1 U18894 ( .D(n18279), .ENB(m4s8_cyc), .Q(n9450) );
  LSDNENX1 U18895 ( .D(n18278), .ENB(test_so26), .Q(n13166) );
  LSDNENX1 U18896 ( .D(n18277), .ENB(m4s13_cyc), .Q(n11000) );
  LSDNENX1 U18897 ( .D(n18276), .ENB(test_so27), .Q(n10381) );
  LSDNENX1 U18898 ( .D(n18275), .ENB(m4s1_cyc), .Q(n11929) );
  LSDNENX1 U18899 ( .D(n18274), .ENB(m4s4_cyc), .Q(n12857) );
  NOR2X0 U18900 ( .IN1(n14430), .IN2(n14431), .QN(n17774) );
  NOR2X0 U18901 ( .IN1(n14440), .IN2(n14441), .QN(n17775) );
  NOR2X0 U18902 ( .IN1(n14350), .IN2(n14351), .QN(n17766) );
  NOR2X0 U18903 ( .IN1(n14360), .IN2(n14361), .QN(n17767) );
  NOR2X0 U18904 ( .IN1(n14370), .IN2(n14371), .QN(n17768) );
  NOR2X0 U18905 ( .IN1(n14380), .IN2(n14381), .QN(n17769) );
  NOR2X0 U18906 ( .IN1(n14470), .IN2(n14471), .QN(n17778) );
  NOR2X0 U18907 ( .IN1(n14480), .IN2(n14481), .QN(n17779) );
  NOR2X0 U18908 ( .IN1(n14400), .IN2(n14401), .QN(n17771) );
  NBUFFX2 U18909 ( .IN(n11501), .Q(n18262) );
  NBUFFX2 U18910 ( .IN(n9953), .Q(n18263) );
  NBUFFX2 U18911 ( .IN(n10572), .Q(n18264) );
  INVX0 U18912 ( .IN(n13935), .QN(n2843) );
  INVX0 U18913 ( .IN(n13963), .QN(n3257) );
  NAND4X0 U18914 ( .IN1(n9466), .IN2(n9467), .IN3(n9468), .IN4(n9469), .QN(
        n9403) );
  NAND4X0 U18915 ( .IN1(n13182), .IN2(n13183), .IN3(n13184), .IN4(n13185), 
        .QN(n13119) );
  NAND4X0 U18916 ( .IN1(n11016), .IN2(n11017), .IN3(n11018), .IN4(n11019), 
        .QN(n10953) );
  NAND4X0 U18917 ( .IN1(n10397), .IN2(n10398), .IN3(n10399), .IN4(n10400), 
        .QN(n10334) );
  NAND4X0 U18918 ( .IN1(n11945), .IN2(n11946), .IN3(n11947), .IN4(n11948), 
        .QN(n11882) );
  NAND4X0 U18919 ( .IN1(n12873), .IN2(n12874), .IN3(n12875), .IN4(n12876), 
        .QN(n12810) );
  NAND4X0 U18920 ( .IN1(n10706), .IN2(n10707), .IN3(n10708), .IN4(n10709), 
        .QN(n10643) );
  NAND4X0 U18921 ( .IN1(n10087), .IN2(n10088), .IN3(n10089), .IN4(n10090), 
        .QN(n10024) );
  NAND4X0 U18922 ( .IN1(n11635), .IN2(n11636), .IN3(n11637), .IN4(n11638), 
        .QN(n11572) );
  NAND4X0 U18923 ( .IN1(n13800), .IN2(n13801), .IN3(n13802), .IN4(n13803), 
        .QN(n13737) );
  NAND4X0 U18924 ( .IN1(n12564), .IN2(n12565), .IN3(n12566), .IN4(n12567), 
        .QN(n12501) );
  NAND4X0 U18925 ( .IN1(n9777), .IN2(n9778), .IN3(n9779), .IN4(n9780), .QN(
        n9714) );
  NAND4X0 U18926 ( .IN1(n13491), .IN2(n13492), .IN3(n13493), .IN4(n13494), 
        .QN(n13428) );
  NAND4X0 U18927 ( .IN1(n11325), .IN2(n11326), .IN3(n11327), .IN4(n11328), 
        .QN(n11262) );
  NAND4X0 U18928 ( .IN1(n12255), .IN2(n12256), .IN3(n12257), .IN4(n12258), 
        .QN(n12192) );
  NBUFFX2 U18929 ( .IN(m4s12_cyc), .Q(n18327) );
  NBUFFX2 U18930 ( .IN(m4s10_cyc), .Q(n18323) );
  NBUFFX2 U18931 ( .IN(m4s4_cyc), .Q(n18329) );
  NBUFFX2 U18932 ( .IN(m4s0_cyc), .Q(n18321) );
  NBUFFX2 U18933 ( .IN(m4s13_cyc), .Q(n18328) );
  NBUFFX2 U18934 ( .IN(test_so27), .Q(n18324) );
  NBUFFX2 U18935 ( .IN(test_so26), .Q(n18330) );
  NBUFFX2 U18936 ( .IN(m4s1_cyc), .Q(n18322) );
  NBUFFX2 U18937 ( .IN(m4s8_cyc), .Q(n18319) );
  LSDNENX1 U18938 ( .D(n14277), .ENB(m4s15_cyc), .Q(n13944) );
  OR2X1 U18939 ( .IN1(n13357), .IN2(n18282), .Q(n13475) );
  OR2X1 U18940 ( .IN1(n11191), .IN2(n18281), .Q(n11309) );
  OR2X1 U18941 ( .IN1(n12430), .IN2(n18284), .Q(n12548) );
  OR2X1 U18942 ( .IN1(n12121), .IN2(n18280), .Q(n12239) );
  OR2X1 U18943 ( .IN1(n9643), .IN2(n18283), .Q(n9761) );
  NBUFFX2 U18944 ( .IN(n12739), .Q(n18274) );
  NBUFFX2 U18945 ( .IN(n11811), .Q(n18275) );
  NBUFFX2 U18946 ( .IN(n10263), .Q(n18276) );
  NBUFFX2 U18947 ( .IN(n10882), .Q(n18277) );
  NBUFFX2 U18948 ( .IN(n13048), .Q(n18278) );
  NBUFFX2 U18949 ( .IN(n9332), .Q(n18279) );
  NAND2X1 U18950 ( .IN1(conf15_8_), .IN2(n17939), .QN(n14277) );
  OR2X1 U18951 ( .IN1(n13666), .IN2(n18285), .Q(n13784) );
  INVX0 U18952 ( .IN(n19634), .QN(n19621) );
  INVX0 U18953 ( .IN(n19634), .QN(n19622) );
  INVX0 U18954 ( .IN(n19635), .QN(n19623) );
  INVX0 U18955 ( .IN(n19635), .QN(n19624) );
  INVX0 U18956 ( .IN(n19635), .QN(n19625) );
  INVX0 U18957 ( .IN(n19635), .QN(n19626) );
  INVX0 U18958 ( .IN(n19635), .QN(n19627) );
  INVX0 U18959 ( .IN(n19635), .QN(n19628) );
  INVX0 U18960 ( .IN(n19635), .QN(n19629) );
  INVX0 U18961 ( .IN(n19635), .QN(n19630) );
  INVX0 U18962 ( .IN(n19501), .QN(n19485) );
  INVX0 U18963 ( .IN(n19502), .QN(n19486) );
  INVX0 U18964 ( .IN(n19501), .QN(n19487) );
  INVX0 U18965 ( .IN(n19501), .QN(n19488) );
  INVX0 U18966 ( .IN(n17885), .QN(n19489) );
  INVX0 U18967 ( .IN(n17885), .QN(n19490) );
  INVX0 U18968 ( .IN(n19502), .QN(n19491) );
  INVX0 U18969 ( .IN(n19503), .QN(n19498) );
  INVX0 U18970 ( .IN(n19502), .QN(n19492) );
  INVX0 U18971 ( .IN(n19501), .QN(n19493) );
  INVX0 U18972 ( .IN(n19503), .QN(n19494) );
  INVX0 U18973 ( .IN(n19503), .QN(n19495) );
  INVX0 U18974 ( .IN(n19503), .QN(n19496) );
  INVX0 U18975 ( .IN(n19369), .QN(n19353) );
  INVX0 U18976 ( .IN(n19370), .QN(n19354) );
  INVX0 U18977 ( .IN(n19369), .QN(n19355) );
  INVX0 U18978 ( .IN(n19369), .QN(n19356) );
  INVX0 U18979 ( .IN(n17886), .QN(n19357) );
  INVX0 U18980 ( .IN(n17886), .QN(n19358) );
  INVX0 U18981 ( .IN(n19370), .QN(n19359) );
  INVX0 U18982 ( .IN(n19371), .QN(n19366) );
  INVX0 U18983 ( .IN(n19370), .QN(n19360) );
  INVX0 U18984 ( .IN(n19369), .QN(n19361) );
  INVX0 U18985 ( .IN(n19371), .QN(n19362) );
  INVX0 U18986 ( .IN(n19371), .QN(n19363) );
  INVX0 U18987 ( .IN(n19371), .QN(n19364) );
  INVX0 U18988 ( .IN(n19237), .QN(n19221) );
  INVX0 U18989 ( .IN(n19238), .QN(n19222) );
  INVX0 U18990 ( .IN(n19237), .QN(n19223) );
  INVX0 U18991 ( .IN(n19237), .QN(n19224) );
  INVX0 U18992 ( .IN(n17887), .QN(n19225) );
  INVX0 U18993 ( .IN(n17887), .QN(n19226) );
  INVX0 U18994 ( .IN(n19238), .QN(n19227) );
  INVX0 U18995 ( .IN(n19239), .QN(n19234) );
  INVX0 U18996 ( .IN(n19238), .QN(n19228) );
  INVX0 U18997 ( .IN(n19237), .QN(n19229) );
  INVX0 U18998 ( .IN(n19239), .QN(n19230) );
  INVX0 U18999 ( .IN(n19239), .QN(n19231) );
  INVX0 U19000 ( .IN(n19239), .QN(n19232) );
  INVX0 U19001 ( .IN(n19105), .QN(n19089) );
  INVX0 U19002 ( .IN(n19106), .QN(n19090) );
  INVX0 U19003 ( .IN(n19105), .QN(n19091) );
  INVX0 U19004 ( .IN(n19105), .QN(n19092) );
  INVX0 U19005 ( .IN(n17888), .QN(n19093) );
  INVX0 U19006 ( .IN(n17888), .QN(n19094) );
  INVX0 U19007 ( .IN(n19106), .QN(n19095) );
  INVX0 U19008 ( .IN(n19107), .QN(n19102) );
  INVX0 U19009 ( .IN(n19106), .QN(n19096) );
  INVX0 U19010 ( .IN(n19105), .QN(n19097) );
  INVX0 U19011 ( .IN(n19107), .QN(n19098) );
  INVX0 U19012 ( .IN(n19107), .QN(n19099) );
  INVX0 U19013 ( .IN(n19107), .QN(n19100) );
  INVX0 U19014 ( .IN(n18974), .QN(n18963) );
  INVX0 U19015 ( .IN(n18973), .QN(n18957) );
  INVX0 U19016 ( .IN(n18975), .QN(n18958) );
  INVX0 U19017 ( .IN(n18973), .QN(n18959) );
  INVX0 U19018 ( .IN(n18973), .QN(n18960) );
  INVX0 U19019 ( .IN(n18974), .QN(n18961) );
  INVX0 U19020 ( .IN(n18974), .QN(n18962) );
  INVX0 U19021 ( .IN(n18975), .QN(n18964) );
  INVX0 U19022 ( .IN(n17889), .QN(n18969) );
  INVX0 U19023 ( .IN(n18975), .QN(n18965) );
  INVX0 U19024 ( .IN(n17889), .QN(n18966) );
  INVX0 U19025 ( .IN(n18973), .QN(n18967) );
  INVX0 U19026 ( .IN(n18972), .QN(n18968) );
  INVX0 U19027 ( .IN(n20688), .QN(n20677) );
  INVX0 U19028 ( .IN(n20687), .QN(n20671) );
  INVX0 U19029 ( .IN(n20689), .QN(n20672) );
  INVX0 U19030 ( .IN(n20687), .QN(n20673) );
  INVX0 U19031 ( .IN(n20687), .QN(n20674) );
  INVX0 U19032 ( .IN(n20688), .QN(n20675) );
  INVX0 U19033 ( .IN(n20688), .QN(n20676) );
  INVX0 U19034 ( .IN(n20689), .QN(n20678) );
  INVX0 U19035 ( .IN(n17890), .QN(n20683) );
  INVX0 U19036 ( .IN(n20689), .QN(n20679) );
  INVX0 U19037 ( .IN(n17890), .QN(n20680) );
  INVX0 U19038 ( .IN(n20687), .QN(n20681) );
  INVX0 U19039 ( .IN(n20686), .QN(n20682) );
  INVX0 U19040 ( .IN(n20556), .QN(n20544) );
  INVX0 U19041 ( .IN(n20555), .QN(n20539) );
  INVX0 U19042 ( .IN(n20557), .QN(n20540) );
  INVX0 U19043 ( .IN(n20555), .QN(n20541) );
  INVX0 U19044 ( .IN(n20555), .QN(n20542) );
  INVX0 U19045 ( .IN(n20556), .QN(n20543) );
  INVX0 U19046 ( .IN(n20557), .QN(n20545) );
  INVX0 U19047 ( .IN(n20558), .QN(n20551) );
  INVX0 U19048 ( .IN(n20554), .QN(n20552) );
  INVX0 U19049 ( .IN(n20557), .QN(n20546) );
  INVX0 U19050 ( .IN(n20555), .QN(n20547) );
  INVX0 U19051 ( .IN(n20556), .QN(n20548) );
  INVX0 U19052 ( .IN(n20558), .QN(n20549) );
  INVX0 U19053 ( .IN(n20558), .QN(n20550) );
  INVX0 U19054 ( .IN(n20424), .QN(n20412) );
  INVX0 U19055 ( .IN(n20423), .QN(n20407) );
  INVX0 U19056 ( .IN(n20425), .QN(n20408) );
  INVX0 U19057 ( .IN(n20423), .QN(n20409) );
  INVX0 U19058 ( .IN(n20423), .QN(n20410) );
  INVX0 U19059 ( .IN(n20424), .QN(n20411) );
  INVX0 U19060 ( .IN(n20425), .QN(n20413) );
  INVX0 U19061 ( .IN(n20426), .QN(n20419) );
  INVX0 U19062 ( .IN(n20422), .QN(n20420) );
  INVX0 U19063 ( .IN(n20425), .QN(n20414) );
  INVX0 U19064 ( .IN(n20423), .QN(n20415) );
  INVX0 U19065 ( .IN(n20424), .QN(n20416) );
  INVX0 U19066 ( .IN(n20426), .QN(n20417) );
  INVX0 U19067 ( .IN(n20426), .QN(n20418) );
  INVX0 U19068 ( .IN(n20292), .QN(n20280) );
  INVX0 U19069 ( .IN(n20291), .QN(n20275) );
  INVX0 U19070 ( .IN(n20293), .QN(n20276) );
  INVX0 U19071 ( .IN(n20291), .QN(n20277) );
  INVX0 U19072 ( .IN(n20291), .QN(n20278) );
  INVX0 U19073 ( .IN(n20292), .QN(n20279) );
  INVX0 U19074 ( .IN(n20293), .QN(n20281) );
  INVX0 U19075 ( .IN(n20294), .QN(n20287) );
  INVX0 U19076 ( .IN(n20290), .QN(n20288) );
  INVX0 U19077 ( .IN(n20293), .QN(n20282) );
  INVX0 U19078 ( .IN(n20291), .QN(n20283) );
  INVX0 U19079 ( .IN(n20292), .QN(n20284) );
  INVX0 U19080 ( .IN(n20294), .QN(n20285) );
  INVX0 U19081 ( .IN(n20294), .QN(n20286) );
  INVX0 U19082 ( .IN(n20159), .QN(n20143) );
  INVX0 U19083 ( .IN(n20160), .QN(n20144) );
  INVX0 U19084 ( .IN(n20159), .QN(n20145) );
  INVX0 U19085 ( .IN(n20159), .QN(n20146) );
  INVX0 U19086 ( .IN(n17894), .QN(n20147) );
  INVX0 U19087 ( .IN(n17894), .QN(n20148) );
  INVX0 U19088 ( .IN(n20160), .QN(n20149) );
  INVX0 U19089 ( .IN(n20161), .QN(n20156) );
  INVX0 U19090 ( .IN(n20160), .QN(n20150) );
  INVX0 U19091 ( .IN(n20159), .QN(n20151) );
  INVX0 U19092 ( .IN(n20161), .QN(n20152) );
  INVX0 U19093 ( .IN(n20161), .QN(n20153) );
  INVX0 U19094 ( .IN(n20161), .QN(n20154) );
  INVX0 U19095 ( .IN(n20029), .QN(n20018) );
  INVX0 U19096 ( .IN(n20028), .QN(n20012) );
  INVX0 U19097 ( .IN(n20030), .QN(n20013) );
  INVX0 U19098 ( .IN(n20028), .QN(n20014) );
  INVX0 U19099 ( .IN(n20028), .QN(n20015) );
  INVX0 U19100 ( .IN(n20029), .QN(n20016) );
  INVX0 U19101 ( .IN(n20029), .QN(n20017) );
  INVX0 U19102 ( .IN(n20030), .QN(n20019) );
  INVX0 U19103 ( .IN(n17895), .QN(n20024) );
  INVX0 U19104 ( .IN(n20030), .QN(n20020) );
  INVX0 U19105 ( .IN(n17895), .QN(n20021) );
  INVX0 U19106 ( .IN(n20028), .QN(n20022) );
  INVX0 U19107 ( .IN(n20027), .QN(n20023) );
  INVX0 U19108 ( .IN(n19898), .QN(n19887) );
  INVX0 U19109 ( .IN(n19897), .QN(n19881) );
  INVX0 U19110 ( .IN(n19899), .QN(n19882) );
  INVX0 U19111 ( .IN(n19897), .QN(n19883) );
  INVX0 U19112 ( .IN(n19897), .QN(n19884) );
  INVX0 U19113 ( .IN(n19898), .QN(n19885) );
  INVX0 U19114 ( .IN(n19898), .QN(n19886) );
  INVX0 U19115 ( .IN(n19899), .QN(n19888) );
  INVX0 U19116 ( .IN(n17896), .QN(n19893) );
  INVX0 U19117 ( .IN(n19899), .QN(n19889) );
  INVX0 U19118 ( .IN(n17896), .QN(n19890) );
  INVX0 U19119 ( .IN(n19897), .QN(n19891) );
  INVX0 U19120 ( .IN(n19896), .QN(n19892) );
  INVX0 U19121 ( .IN(n19766), .QN(n19755) );
  INVX0 U19122 ( .IN(n19765), .QN(n19749) );
  INVX0 U19123 ( .IN(n19767), .QN(n19750) );
  INVX0 U19124 ( .IN(n19765), .QN(n19751) );
  INVX0 U19125 ( .IN(n19765), .QN(n19752) );
  INVX0 U19126 ( .IN(n19766), .QN(n19753) );
  INVX0 U19127 ( .IN(n19766), .QN(n19754) );
  INVX0 U19128 ( .IN(n19767), .QN(n19756) );
  INVX0 U19129 ( .IN(n17897), .QN(n19761) );
  INVX0 U19130 ( .IN(n19767), .QN(n19757) );
  INVX0 U19131 ( .IN(n17897), .QN(n19758) );
  INVX0 U19132 ( .IN(n19765), .QN(n19759) );
  INVX0 U19133 ( .IN(n19764), .QN(n19760) );
  INVX0 U19134 ( .IN(n18842), .QN(n18831) );
  INVX0 U19135 ( .IN(n18841), .QN(n18825) );
  INVX0 U19136 ( .IN(n18843), .QN(n18826) );
  INVX0 U19137 ( .IN(n18841), .QN(n18827) );
  INVX0 U19138 ( .IN(n18841), .QN(n18828) );
  INVX0 U19139 ( .IN(n18842), .QN(n18829) );
  INVX0 U19140 ( .IN(n18842), .QN(n18830) );
  INVX0 U19141 ( .IN(n18843), .QN(n18832) );
  INVX0 U19142 ( .IN(n17898), .QN(n18837) );
  INVX0 U19143 ( .IN(n18843), .QN(n18833) );
  INVX0 U19144 ( .IN(n17898), .QN(n18834) );
  INVX0 U19145 ( .IN(n18841), .QN(n18835) );
  INVX0 U19146 ( .IN(n18840), .QN(n18836) );
  INVX0 U19147 ( .IN(n20990), .QN(n20874) );
  INVX0 U19148 ( .IN(n20991), .QN(n20875) );
  INVX0 U19149 ( .IN(n20992), .QN(n20876) );
  INVX0 U19150 ( .IN(n20993), .QN(n20877) );
  INVX0 U19151 ( .IN(n20994), .QN(n20878) );
  INVX0 U19152 ( .IN(n20995), .QN(n20879) );
  INVX0 U19153 ( .IN(n20996), .QN(n20880) );
  INVX0 U19154 ( .IN(n20997), .QN(n20881) );
  INVX0 U19155 ( .IN(n20998), .QN(n20882) );
  INVX0 U19156 ( .IN(n20999), .QN(n20883) );
  INVX0 U19157 ( .IN(n21000), .QN(n20884) );
  INVX0 U19158 ( .IN(n21001), .QN(n20885) );
  INVX0 U19159 ( .IN(n21002), .QN(n20886) );
  INVX0 U19160 ( .IN(n21003), .QN(n20887) );
  INVX0 U19161 ( .IN(n21004), .QN(n20888) );
  INVX0 U19162 ( .IN(n21005), .QN(n20889) );
  INVX0 U19163 ( .IN(n21006), .QN(n20890) );
  INVX0 U19164 ( .IN(n21007), .QN(n20891) );
  INVX0 U19165 ( .IN(n21008), .QN(n20892) );
  INVX0 U19166 ( .IN(n21009), .QN(n20893) );
  INVX0 U19167 ( .IN(n21010), .QN(n20894) );
  INVX0 U19168 ( .IN(n21011), .QN(n20895) );
  INVX0 U19169 ( .IN(n21012), .QN(n20896) );
  INVX0 U19170 ( .IN(n21013), .QN(n20897) );
  INVX0 U19171 ( .IN(n21014), .QN(n20898) );
  INVX0 U19172 ( .IN(n21015), .QN(n20899) );
  INVX0 U19173 ( .IN(n21016), .QN(n20900) );
  INVX0 U19174 ( .IN(n21017), .QN(n20901) );
  INVX0 U19175 ( .IN(n21018), .QN(n20902) );
  INVX0 U19176 ( .IN(n21018), .QN(n20903) );
  INVX0 U19177 ( .IN(n21018), .QN(n20904) );
  INVX0 U19178 ( .IN(n21019), .QN(n20905) );
  INVX0 U19179 ( .IN(n21019), .QN(n20906) );
  INVX0 U19180 ( .IN(n21019), .QN(n20907) );
  INVX0 U19181 ( .IN(n21020), .QN(n20908) );
  INVX0 U19182 ( .IN(n21020), .QN(n20909) );
  INVX0 U19183 ( .IN(n21020), .QN(n20910) );
  INVX0 U19184 ( .IN(n21021), .QN(n20911) );
  INVX0 U19185 ( .IN(n21021), .QN(n20912) );
  INVX0 U19186 ( .IN(n21022), .QN(n20913) );
  INVX0 U19187 ( .IN(n21022), .QN(n20914) );
  INVX0 U19188 ( .IN(n21024), .QN(n20919) );
  INVX0 U19189 ( .IN(n21024), .QN(n20920) );
  INVX0 U19190 ( .IN(n21024), .QN(n20921) );
  INVX0 U19191 ( .IN(n21025), .QN(n20922) );
  INVX0 U19192 ( .IN(n21025), .QN(n20923) );
  INVX0 U19193 ( .IN(n21025), .QN(n20924) );
  INVX0 U19194 ( .IN(n21026), .QN(n20925) );
  INVX0 U19195 ( .IN(n21026), .QN(n20926) );
  INVX0 U19196 ( .IN(n21026), .QN(n20927) );
  INVX0 U19197 ( .IN(n21077), .QN(n20928) );
  INVX0 U19198 ( .IN(n21038), .QN(n20929) );
  INVX0 U19199 ( .IN(n21027), .QN(n20930) );
  INVX0 U19200 ( .IN(n21027), .QN(n20931) );
  INVX0 U19201 ( .IN(n21027), .QN(n20932) );
  INVX0 U19202 ( .IN(n21027), .QN(n20933) );
  INVX0 U19203 ( .IN(n21028), .QN(n20934) );
  INVX0 U19204 ( .IN(n21022), .QN(n20915) );
  INVX0 U19205 ( .IN(n21023), .QN(n20916) );
  INVX0 U19206 ( .IN(n21023), .QN(n20918) );
  INVX0 U19207 ( .IN(n21023), .QN(n20917) );
  INVX0 U19208 ( .IN(n21028), .QN(n20935) );
  INVX0 U19209 ( .IN(n21028), .QN(n20936) );
  INVX0 U19210 ( .IN(n21029), .QN(n20937) );
  INVX0 U19211 ( .IN(n21029), .QN(n20938) );
  INVX0 U19212 ( .IN(n21029), .QN(n20939) );
  INVX0 U19213 ( .IN(n21030), .QN(n20940) );
  INVX0 U19214 ( .IN(n21030), .QN(n20941) );
  INVX0 U19215 ( .IN(n21030), .QN(n20942) );
  INVX0 U19216 ( .IN(n21031), .QN(n20943) );
  INVX0 U19217 ( .IN(n21031), .QN(n20944) );
  INVX0 U19218 ( .IN(n21031), .QN(n20945) );
  INVX0 U19219 ( .IN(n21032), .QN(n20946) );
  INVX0 U19220 ( .IN(n21032), .QN(n20947) );
  INVX0 U19221 ( .IN(n21032), .QN(n20948) );
  INVX0 U19222 ( .IN(n21033), .QN(n20949) );
  INVX0 U19223 ( .IN(n21033), .QN(n20950) );
  INVX0 U19224 ( .IN(n21033), .QN(n20951) );
  INVX0 U19225 ( .IN(n21034), .QN(n20952) );
  INVX0 U19226 ( .IN(n21034), .QN(n20953) );
  INVX0 U19227 ( .IN(n21034), .QN(n20954) );
  INVX0 U19228 ( .IN(n21035), .QN(n20955) );
  INVX0 U19229 ( .IN(n21035), .QN(n20956) );
  INVX0 U19230 ( .IN(n21035), .QN(n20957) );
  INVX0 U19231 ( .IN(n21036), .QN(n20958) );
  INVX0 U19232 ( .IN(n21036), .QN(n20959) );
  INVX0 U19233 ( .IN(n21036), .QN(n20960) );
  INVX0 U19234 ( .IN(n21037), .QN(n20961) );
  INVX0 U19235 ( .IN(n21037), .QN(n20962) );
  INVX0 U19236 ( .IN(n21037), .QN(n20963) );
  INVX0 U19237 ( .IN(n21038), .QN(n20964) );
  INVX0 U19238 ( .IN(n21038), .QN(n20965) );
  INVX0 U19239 ( .IN(n21038), .QN(n20966) );
  INVX0 U19240 ( .IN(n21039), .QN(n20967) );
  INVX0 U19241 ( .IN(n21039), .QN(n20968) );
  INVX0 U19242 ( .IN(n21039), .QN(n20969) );
  INVX0 U19243 ( .IN(n21040), .QN(n20970) );
  INVX0 U19244 ( .IN(n21040), .QN(n20971) );
  INVX0 U19245 ( .IN(n21040), .QN(n20972) );
  INVX0 U19246 ( .IN(n21041), .QN(n20973) );
  INVX0 U19247 ( .IN(n21041), .QN(n20974) );
  INVX0 U19248 ( .IN(n21041), .QN(n20975) );
  INVX0 U19249 ( .IN(n21042), .QN(n20976) );
  INVX0 U19250 ( .IN(n21042), .QN(n20977) );
  INVX0 U19251 ( .IN(n21042), .QN(n20978) );
  INVX0 U19252 ( .IN(n21043), .QN(n20979) );
  INVX0 U19253 ( .IN(n21043), .QN(n20980) );
  INVX0 U19254 ( .IN(n21043), .QN(n20981) );
  INVX0 U19255 ( .IN(n21044), .QN(n20982) );
  INVX0 U19256 ( .IN(n21044), .QN(n20983) );
  INVX0 U19257 ( .IN(n21044), .QN(n20984) );
  INVX0 U19258 ( .IN(n17780), .QN(n18816) );
  INVX0 U19259 ( .IN(n19633), .QN(n19619) );
  INVX0 U19260 ( .IN(n19633), .QN(n19620) );
  INVX0 U19261 ( .IN(n19614), .QN(n19634) );
  INVX0 U19262 ( .IN(n19733), .QN(n19720) );
  INVX0 U19263 ( .IN(n19700), .QN(n19687) );
  INVX0 U19264 ( .IN(n19667), .QN(n19654) );
  INVX0 U19265 ( .IN(n21060), .QN(n21001) );
  INVX0 U19266 ( .IN(n21060), .QN(n21000) );
  INVX0 U19267 ( .IN(n21065), .QN(n20990) );
  INVX0 U19268 ( .IN(n21062), .QN(n20996) );
  INVX0 U19269 ( .IN(n21061), .QN(n20998) );
  INVX0 U19270 ( .IN(n21064), .QN(n20992) );
  INVX0 U19271 ( .IN(n21065), .QN(n20991) );
  INVX0 U19272 ( .IN(n21062), .QN(n20997) );
  INVX0 U19273 ( .IN(n21064), .QN(n20993) );
  INVX0 U19274 ( .IN(n21063), .QN(n20995) );
  INVX0 U19275 ( .IN(n21063), .QN(n20994) );
  INVX0 U19276 ( .IN(n21061), .QN(n20999) );
  INVX0 U19277 ( .IN(n19622), .QN(n19635) );
  INVX0 U19278 ( .IN(n19481), .QN(n19501) );
  INVX0 U19279 ( .IN(n19481), .QN(n19502) );
  INVX0 U19280 ( .IN(n19481), .QN(n19503) );
  INVX0 U19281 ( .IN(n19349), .QN(n19369) );
  INVX0 U19282 ( .IN(n19349), .QN(n19370) );
  INVX0 U19283 ( .IN(n19349), .QN(n19371) );
  INVX0 U19284 ( .IN(n19217), .QN(n19237) );
  INVX0 U19285 ( .IN(n19217), .QN(n19238) );
  INVX0 U19286 ( .IN(n19217), .QN(n19239) );
  INVX0 U19287 ( .IN(n19085), .QN(n19105) );
  INVX0 U19288 ( .IN(n19085), .QN(n19106) );
  INVX0 U19289 ( .IN(n19085), .QN(n19107) );
  INVX0 U19290 ( .IN(n18953), .QN(n18973) );
  INVX0 U19291 ( .IN(n18953), .QN(n18974) );
  INVX0 U19292 ( .IN(n18953), .QN(n18975) );
  INVX0 U19293 ( .IN(n20667), .QN(n20687) );
  INVX0 U19294 ( .IN(n20667), .QN(n20688) );
  INVX0 U19295 ( .IN(n20667), .QN(n20689) );
  INVX0 U19296 ( .IN(n20535), .QN(n20555) );
  INVX0 U19297 ( .IN(n20535), .QN(n20556) );
  INVX0 U19298 ( .IN(n20535), .QN(n20557) );
  INVX0 U19299 ( .IN(n20535), .QN(n20558) );
  INVX0 U19300 ( .IN(n20403), .QN(n20423) );
  INVX0 U19301 ( .IN(n20403), .QN(n20424) );
  INVX0 U19302 ( .IN(n20403), .QN(n20425) );
  INVX0 U19303 ( .IN(n20403), .QN(n20426) );
  INVX0 U19304 ( .IN(n20271), .QN(n20291) );
  INVX0 U19305 ( .IN(n20271), .QN(n20292) );
  INVX0 U19306 ( .IN(n20271), .QN(n20293) );
  INVX0 U19307 ( .IN(n20271), .QN(n20294) );
  INVX0 U19308 ( .IN(n20139), .QN(n20159) );
  INVX0 U19309 ( .IN(n20139), .QN(n20160) );
  INVX0 U19310 ( .IN(n20139), .QN(n20161) );
  INVX0 U19311 ( .IN(n20008), .QN(n20028) );
  INVX0 U19312 ( .IN(n20008), .QN(n20029) );
  INVX0 U19313 ( .IN(n20008), .QN(n20030) );
  INVX0 U19314 ( .IN(n19877), .QN(n19897) );
  INVX0 U19315 ( .IN(n19877), .QN(n19898) );
  INVX0 U19316 ( .IN(n19877), .QN(n19899) );
  INVX0 U19317 ( .IN(n19745), .QN(n19765) );
  INVX0 U19318 ( .IN(n19745), .QN(n19766) );
  INVX0 U19319 ( .IN(n19745), .QN(n19767) );
  INVX0 U19320 ( .IN(n18821), .QN(n18841) );
  INVX0 U19321 ( .IN(n18821), .QN(n18842) );
  INVX0 U19322 ( .IN(n18821), .QN(n18843) );
  INVX0 U19323 ( .IN(n19733), .QN(n19722) );
  INVX0 U19324 ( .IN(n19700), .QN(n19689) );
  INVX0 U19325 ( .IN(n19667), .QN(n19656) );
  INVX0 U19326 ( .IN(n19734), .QN(n19723) );
  INVX0 U19327 ( .IN(n19701), .QN(n19690) );
  INVX0 U19328 ( .IN(n19668), .QN(n19657) );
  INVX0 U19329 ( .IN(n19632), .QN(n19631) );
  INVX0 U19330 ( .IN(n19734), .QN(n19728) );
  INVX0 U19331 ( .IN(n19701), .QN(n19694) );
  INVX0 U19332 ( .IN(n19668), .QN(n19661) );
  INVX0 U19333 ( .IN(n19734), .QN(n19724) );
  INVX0 U19334 ( .IN(n19701), .QN(n19691) );
  INVX0 U19335 ( .IN(n19668), .QN(n19658) );
  INVX0 U19336 ( .IN(n19734), .QN(n19725) );
  INVX0 U19337 ( .IN(n19701), .QN(n19692) );
  INVX0 U19338 ( .IN(n19668), .QN(n19659) );
  INVX0 U19339 ( .IN(n19734), .QN(n19726) );
  INVX0 U19340 ( .IN(n19701), .QN(n19693) );
  INVX0 U19341 ( .IN(n19668), .QN(n19660) );
  INVX0 U19342 ( .IN(n19734), .QN(n19727) );
  INVX0 U19343 ( .IN(n19734), .QN(n19729) );
  INVX0 U19344 ( .IN(n19701), .QN(n19695) );
  INVX0 U19345 ( .IN(n19668), .QN(n19662) );
  INVX0 U19346 ( .IN(n19701), .QN(n19696) );
  INVX0 U19347 ( .IN(n19668), .QN(n19663) );
  INVX0 U19348 ( .IN(n19504), .QN(n19499) );
  INVX0 U19349 ( .IN(n19568), .QN(n19556) );
  INVX0 U19350 ( .IN(n19500), .QN(n19482) );
  INVX0 U19351 ( .IN(n19500), .QN(n19483) );
  INVX0 U19352 ( .IN(n19500), .QN(n19484) );
  INVX0 U19353 ( .IN(n19600), .QN(n19584) );
  INVX0 U19354 ( .IN(n19568), .QN(n19551) );
  INVX0 U19355 ( .IN(n19534), .QN(n19518) );
  INVX0 U19356 ( .IN(n19601), .QN(n19585) );
  INVX0 U19357 ( .IN(n19569), .QN(n19552) );
  INVX0 U19358 ( .IN(n19535), .QN(n19519) );
  INVX0 U19359 ( .IN(n19600), .QN(n19586) );
  INVX0 U19360 ( .IN(n19568), .QN(n19553) );
  INVX0 U19361 ( .IN(n19534), .QN(n19520) );
  INVX0 U19362 ( .IN(n19600), .QN(n19587) );
  INVX0 U19363 ( .IN(n19568), .QN(n19554) );
  INVX0 U19364 ( .IN(n19534), .QN(n19521) );
  INVX0 U19365 ( .IN(n19600), .QN(n19588) );
  INVX0 U19366 ( .IN(n19568), .QN(n19555) );
  INVX0 U19367 ( .IN(n17899), .QN(n19522) );
  INVX0 U19368 ( .IN(n17899), .QN(n19523) );
  INVX0 U19369 ( .IN(n19601), .QN(n19589) );
  INVX0 U19370 ( .IN(n19569), .QN(n19557) );
  INVX0 U19371 ( .IN(n19535), .QN(n19524) );
  INVX0 U19372 ( .IN(n19603), .QN(n19595) );
  INVX0 U19373 ( .IN(n19569), .QN(n19563) );
  INVX0 U19374 ( .IN(n19504), .QN(n19497) );
  INVX0 U19375 ( .IN(n19602), .QN(n19597) );
  INVX0 U19376 ( .IN(n19569), .QN(n19565) );
  INVX0 U19377 ( .IN(n19536), .QN(n19531) );
  INVX0 U19378 ( .IN(n19601), .QN(n19590) );
  INVX0 U19379 ( .IN(n19569), .QN(n19558) );
  INVX0 U19380 ( .IN(n19535), .QN(n19525) );
  INVX0 U19381 ( .IN(n17925), .QN(n19591) );
  INVX0 U19382 ( .IN(n19569), .QN(n19559) );
  INVX0 U19383 ( .IN(n19534), .QN(n19526) );
  INVX0 U19384 ( .IN(n19602), .QN(n19592) );
  INVX0 U19385 ( .IN(n19570), .QN(n19560) );
  INVX0 U19386 ( .IN(n19536), .QN(n19527) );
  INVX0 U19387 ( .IN(n19602), .QN(n19593) );
  INVX0 U19388 ( .IN(n19570), .QN(n19561) );
  INVX0 U19389 ( .IN(n19536), .QN(n19528) );
  INVX0 U19390 ( .IN(n19602), .QN(n19594) );
  INVX0 U19391 ( .IN(n19570), .QN(n19562) );
  INVX0 U19392 ( .IN(n19536), .QN(n19529) );
  INVX0 U19393 ( .IN(n19372), .QN(n19367) );
  INVX0 U19394 ( .IN(n17926), .QN(n19455) );
  INVX0 U19395 ( .IN(n19368), .QN(n19350) );
  INVX0 U19396 ( .IN(n19368), .QN(n19351) );
  INVX0 U19397 ( .IN(n19368), .QN(n19352) );
  INVX0 U19398 ( .IN(n19469), .QN(n19452) );
  INVX0 U19399 ( .IN(n19435), .QN(n19419) );
  INVX0 U19400 ( .IN(n19402), .QN(n19386) );
  INVX0 U19401 ( .IN(n19468), .QN(n19453) );
  INVX0 U19402 ( .IN(n19436), .QN(n19420) );
  INVX0 U19403 ( .IN(n19403), .QN(n19387) );
  INVX0 U19404 ( .IN(n19468), .QN(n19454) );
  INVX0 U19405 ( .IN(n19435), .QN(n19421) );
  INVX0 U19406 ( .IN(n19402), .QN(n19388) );
  INVX0 U19407 ( .IN(n19435), .QN(n19422) );
  INVX0 U19408 ( .IN(n19402), .QN(n19389) );
  INVX0 U19409 ( .IN(n17901), .QN(n19423) );
  INVX0 U19410 ( .IN(n17900), .QN(n19390) );
  INVX0 U19411 ( .IN(n17901), .QN(n19424) );
  INVX0 U19412 ( .IN(n17900), .QN(n19391) );
  INVX0 U19413 ( .IN(n19468), .QN(n19456) );
  INVX0 U19414 ( .IN(n19436), .QN(n19425) );
  INVX0 U19415 ( .IN(n19403), .QN(n19392) );
  INVX0 U19416 ( .IN(n19470), .QN(n19464) );
  INVX0 U19417 ( .IN(n19372), .QN(n19365) );
  INVX0 U19418 ( .IN(n19467), .QN(n19465) );
  INVX0 U19419 ( .IN(n19437), .QN(n19432) );
  INVX0 U19420 ( .IN(n19404), .QN(n19399) );
  INVX0 U19421 ( .IN(n19468), .QN(n19457) );
  INVX0 U19422 ( .IN(n19436), .QN(n19426) );
  INVX0 U19423 ( .IN(n19403), .QN(n19393) );
  INVX0 U19424 ( .IN(n19469), .QN(n19458) );
  INVX0 U19425 ( .IN(n19469), .QN(n19459) );
  INVX0 U19426 ( .IN(n19435), .QN(n19427) );
  INVX0 U19427 ( .IN(n19402), .QN(n19394) );
  INVX0 U19428 ( .IN(n19469), .QN(n19460) );
  INVX0 U19429 ( .IN(n19470), .QN(n19461) );
  INVX0 U19430 ( .IN(n19437), .QN(n19428) );
  INVX0 U19431 ( .IN(n19404), .QN(n19395) );
  INVX0 U19432 ( .IN(n19470), .QN(n19462) );
  INVX0 U19433 ( .IN(n19437), .QN(n19429) );
  INVX0 U19434 ( .IN(n19404), .QN(n19396) );
  INVX0 U19435 ( .IN(n19470), .QN(n19463) );
  INVX0 U19436 ( .IN(n19437), .QN(n19430) );
  INVX0 U19437 ( .IN(n19404), .QN(n19397) );
  INVX0 U19438 ( .IN(n19240), .QN(n19235) );
  INVX0 U19439 ( .IN(n17927), .QN(n19323) );
  INVX0 U19440 ( .IN(n19236), .QN(n19218) );
  INVX0 U19441 ( .IN(n19236), .QN(n19219) );
  INVX0 U19442 ( .IN(n19236), .QN(n19220) );
  INVX0 U19443 ( .IN(n19337), .QN(n19320) );
  INVX0 U19444 ( .IN(n19303), .QN(n19287) );
  INVX0 U19445 ( .IN(n19270), .QN(n19254) );
  INVX0 U19446 ( .IN(n19336), .QN(n19321) );
  INVX0 U19447 ( .IN(n19304), .QN(n19288) );
  INVX0 U19448 ( .IN(n19271), .QN(n19255) );
  INVX0 U19449 ( .IN(n19336), .QN(n19322) );
  INVX0 U19450 ( .IN(n19303), .QN(n19289) );
  INVX0 U19451 ( .IN(n19270), .QN(n19256) );
  INVX0 U19452 ( .IN(n19303), .QN(n19290) );
  INVX0 U19453 ( .IN(n19270), .QN(n19257) );
  INVX0 U19454 ( .IN(n17903), .QN(n19291) );
  INVX0 U19455 ( .IN(n17902), .QN(n19258) );
  INVX0 U19456 ( .IN(n17903), .QN(n19292) );
  INVX0 U19457 ( .IN(n17902), .QN(n19259) );
  INVX0 U19458 ( .IN(n19336), .QN(n19324) );
  INVX0 U19459 ( .IN(n19304), .QN(n19293) );
  INVX0 U19460 ( .IN(n19271), .QN(n19260) );
  INVX0 U19461 ( .IN(n19338), .QN(n19332) );
  INVX0 U19462 ( .IN(n19240), .QN(n19233) );
  INVX0 U19463 ( .IN(n19335), .QN(n19333) );
  INVX0 U19464 ( .IN(n19305), .QN(n19300) );
  INVX0 U19465 ( .IN(n19272), .QN(n19267) );
  INVX0 U19466 ( .IN(n19336), .QN(n19325) );
  INVX0 U19467 ( .IN(n19304), .QN(n19294) );
  INVX0 U19468 ( .IN(n19271), .QN(n19261) );
  INVX0 U19469 ( .IN(n19337), .QN(n19326) );
  INVX0 U19470 ( .IN(n19337), .QN(n19327) );
  INVX0 U19471 ( .IN(n19303), .QN(n19295) );
  INVX0 U19472 ( .IN(n19270), .QN(n19262) );
  INVX0 U19473 ( .IN(n19337), .QN(n19328) );
  INVX0 U19474 ( .IN(n19338), .QN(n19329) );
  INVX0 U19475 ( .IN(n19305), .QN(n19296) );
  INVX0 U19476 ( .IN(n19272), .QN(n19263) );
  INVX0 U19477 ( .IN(n19338), .QN(n19330) );
  INVX0 U19478 ( .IN(n19305), .QN(n19297) );
  INVX0 U19479 ( .IN(n19272), .QN(n19264) );
  INVX0 U19480 ( .IN(n19338), .QN(n19331) );
  INVX0 U19481 ( .IN(n19305), .QN(n19298) );
  INVX0 U19482 ( .IN(n19272), .QN(n19265) );
  INVX0 U19483 ( .IN(n19108), .QN(n19103) );
  INVX0 U19484 ( .IN(n17928), .QN(n19191) );
  INVX0 U19485 ( .IN(n19172), .QN(n19161) );
  INVX0 U19486 ( .IN(n19104), .QN(n19086) );
  INVX0 U19487 ( .IN(n19104), .QN(n19087) );
  INVX0 U19488 ( .IN(n19104), .QN(n19088) );
  INVX0 U19489 ( .IN(n19205), .QN(n19188) );
  INVX0 U19490 ( .IN(n19171), .QN(n19155) );
  INVX0 U19491 ( .IN(n19138), .QN(n19122) );
  INVX0 U19492 ( .IN(n19204), .QN(n19189) );
  INVX0 U19493 ( .IN(n19173), .QN(n19156) );
  INVX0 U19494 ( .IN(n19139), .QN(n19123) );
  INVX0 U19495 ( .IN(n19204), .QN(n19190) );
  INVX0 U19496 ( .IN(n19171), .QN(n19157) );
  INVX0 U19497 ( .IN(n19138), .QN(n19124) );
  INVX0 U19498 ( .IN(n19171), .QN(n19158) );
  INVX0 U19499 ( .IN(n19138), .QN(n19125) );
  INVX0 U19500 ( .IN(n19172), .QN(n19159) );
  INVX0 U19501 ( .IN(n17904), .QN(n19126) );
  INVX0 U19502 ( .IN(n19172), .QN(n19160) );
  INVX0 U19503 ( .IN(n17904), .QN(n19127) );
  INVX0 U19504 ( .IN(n19204), .QN(n19192) );
  INVX0 U19505 ( .IN(n19173), .QN(n19162) );
  INVX0 U19506 ( .IN(n19139), .QN(n19128) );
  INVX0 U19507 ( .IN(n19206), .QN(n19200) );
  INVX0 U19508 ( .IN(n17905), .QN(n19167) );
  INVX0 U19509 ( .IN(n19108), .QN(n19101) );
  INVX0 U19510 ( .IN(n19203), .QN(n19201) );
  INVX0 U19511 ( .IN(n19140), .QN(n19135) );
  INVX0 U19512 ( .IN(n19204), .QN(n19193) );
  INVX0 U19513 ( .IN(n19139), .QN(n19129) );
  INVX0 U19514 ( .IN(n19205), .QN(n19194) );
  INVX0 U19515 ( .IN(n19171), .QN(n19163) );
  INVX0 U19516 ( .IN(n19205), .QN(n19195) );
  INVX0 U19517 ( .IN(n19172), .QN(n19164) );
  INVX0 U19518 ( .IN(n19138), .QN(n19130) );
  INVX0 U19519 ( .IN(n19205), .QN(n19196) );
  INVX0 U19520 ( .IN(n19206), .QN(n19197) );
  INVX0 U19521 ( .IN(n19170), .QN(n19165) );
  INVX0 U19522 ( .IN(n19140), .QN(n19131) );
  INVX0 U19523 ( .IN(n19206), .QN(n19198) );
  INVX0 U19524 ( .IN(n19174), .QN(n19166) );
  INVX0 U19525 ( .IN(n19140), .QN(n19132) );
  INVX0 U19526 ( .IN(n19206), .QN(n19199) );
  INVX0 U19527 ( .IN(n19140), .QN(n19133) );
  INVX0 U19528 ( .IN(n18976), .QN(n18971) );
  INVX0 U19529 ( .IN(n17919), .QN(n19059) );
  INVX0 U19530 ( .IN(n19039), .QN(n19027) );
  INVX0 U19531 ( .IN(n19007), .QN(n18996) );
  INVX0 U19532 ( .IN(n18972), .QN(n18954) );
  INVX0 U19533 ( .IN(n18972), .QN(n18955) );
  INVX0 U19534 ( .IN(n18972), .QN(n18956) );
  INVX0 U19535 ( .IN(n19073), .QN(n19056) );
  INVX0 U19536 ( .IN(n19038), .QN(n19021) );
  INVX0 U19537 ( .IN(n19006), .QN(n18990) );
  INVX0 U19538 ( .IN(n19072), .QN(n19057) );
  INVX0 U19539 ( .IN(n19040), .QN(n19022) );
  INVX0 U19540 ( .IN(n19008), .QN(n18991) );
  INVX0 U19541 ( .IN(n19072), .QN(n19058) );
  INVX0 U19542 ( .IN(n19038), .QN(n19023) );
  INVX0 U19543 ( .IN(n19006), .QN(n18992) );
  INVX0 U19544 ( .IN(n19038), .QN(n19024) );
  INVX0 U19545 ( .IN(n19006), .QN(n18993) );
  INVX0 U19546 ( .IN(n19039), .QN(n19025) );
  INVX0 U19547 ( .IN(n19007), .QN(n18994) );
  INVX0 U19548 ( .IN(n19039), .QN(n19026) );
  INVX0 U19549 ( .IN(n19007), .QN(n18995) );
  INVX0 U19550 ( .IN(n19072), .QN(n19060) );
  INVX0 U19551 ( .IN(n19040), .QN(n19028) );
  INVX0 U19552 ( .IN(n19008), .QN(n18997) );
  INVX0 U19553 ( .IN(n19074), .QN(n19068) );
  INVX0 U19554 ( .IN(n19042), .QN(n19035) );
  INVX0 U19555 ( .IN(n17906), .QN(n19004) );
  INVX0 U19556 ( .IN(n18976), .QN(n18970) );
  INVX0 U19557 ( .IN(n19071), .QN(n19069) );
  INVX0 U19558 ( .IN(n19042), .QN(n19037) );
  INVX0 U19559 ( .IN(n19072), .QN(n19061) );
  INVX0 U19560 ( .IN(n19008), .QN(n18998) );
  INVX0 U19561 ( .IN(n19073), .QN(n19062) );
  INVX0 U19562 ( .IN(n19038), .QN(n19029) );
  INVX0 U19563 ( .IN(n19009), .QN(n18999) );
  INVX0 U19564 ( .IN(n19073), .QN(n19063) );
  INVX0 U19565 ( .IN(n19039), .QN(n19030) );
  INVX0 U19566 ( .IN(n19009), .QN(n19000) );
  INVX0 U19567 ( .IN(n19073), .QN(n19064) );
  INVX0 U19568 ( .IN(n19009), .QN(n19001) );
  INVX0 U19569 ( .IN(n19074), .QN(n19065) );
  INVX0 U19570 ( .IN(n19041), .QN(n19031) );
  INVX0 U19571 ( .IN(n17906), .QN(n19002) );
  INVX0 U19572 ( .IN(n19074), .QN(n19066) );
  INVX0 U19573 ( .IN(n19041), .QN(n19032) );
  INVX0 U19574 ( .IN(n19005), .QN(n19003) );
  INVX0 U19575 ( .IN(n19074), .QN(n19067) );
  INVX0 U19576 ( .IN(n19041), .QN(n19033) );
  INVX0 U19577 ( .IN(n19042), .QN(n19034) );
  INVX0 U19578 ( .IN(n20690), .QN(n20685) );
  INVX0 U19579 ( .IN(n17920), .QN(n20773) );
  INVX0 U19580 ( .IN(n20754), .QN(n20743) );
  INVX0 U19581 ( .IN(n20721), .QN(n20710) );
  INVX0 U19582 ( .IN(n20686), .QN(n20668) );
  INVX0 U19583 ( .IN(n20686), .QN(n20669) );
  INVX0 U19584 ( .IN(n20686), .QN(n20670) );
  INVX0 U19585 ( .IN(n20787), .QN(n20770) );
  INVX0 U19586 ( .IN(n20753), .QN(n20737) );
  INVX0 U19587 ( .IN(n20720), .QN(n20704) );
  INVX0 U19588 ( .IN(n20786), .QN(n20771) );
  INVX0 U19589 ( .IN(n20755), .QN(n20738) );
  INVX0 U19590 ( .IN(n20722), .QN(n20705) );
  INVX0 U19591 ( .IN(n20786), .QN(n20772) );
  INVX0 U19592 ( .IN(n20753), .QN(n20739) );
  INVX0 U19593 ( .IN(n20720), .QN(n20706) );
  INVX0 U19594 ( .IN(n20753), .QN(n20740) );
  INVX0 U19595 ( .IN(n20720), .QN(n20707) );
  INVX0 U19596 ( .IN(n20754), .QN(n20741) );
  INVX0 U19597 ( .IN(n20721), .QN(n20708) );
  INVX0 U19598 ( .IN(n20754), .QN(n20742) );
  INVX0 U19599 ( .IN(n20721), .QN(n20709) );
  INVX0 U19600 ( .IN(n20786), .QN(n20774) );
  INVX0 U19601 ( .IN(n20755), .QN(n20744) );
  INVX0 U19602 ( .IN(n20722), .QN(n20711) );
  INVX0 U19603 ( .IN(n20788), .QN(n20782) );
  INVX0 U19604 ( .IN(n17907), .QN(n20749) );
  INVX0 U19605 ( .IN(n17908), .QN(n20718) );
  INVX0 U19606 ( .IN(n20690), .QN(n20684) );
  INVX0 U19607 ( .IN(n20785), .QN(n20783) );
  INVX0 U19608 ( .IN(n20786), .QN(n20775) );
  INVX0 U19609 ( .IN(n20722), .QN(n20712) );
  INVX0 U19610 ( .IN(n20787), .QN(n20776) );
  INVX0 U19611 ( .IN(n20753), .QN(n20745) );
  INVX0 U19612 ( .IN(n20723), .QN(n20713) );
  INVX0 U19613 ( .IN(n20787), .QN(n20777) );
  INVX0 U19614 ( .IN(n20754), .QN(n20746) );
  INVX0 U19615 ( .IN(n20723), .QN(n20714) );
  INVX0 U19616 ( .IN(n20787), .QN(n20778) );
  INVX0 U19617 ( .IN(n20723), .QN(n20715) );
  INVX0 U19618 ( .IN(n20788), .QN(n20779) );
  INVX0 U19619 ( .IN(n20752), .QN(n20747) );
  INVX0 U19620 ( .IN(n17908), .QN(n20716) );
  INVX0 U19621 ( .IN(n20788), .QN(n20780) );
  INVX0 U19622 ( .IN(n20756), .QN(n20748) );
  INVX0 U19623 ( .IN(n20719), .QN(n20717) );
  INVX0 U19624 ( .IN(n20788), .QN(n20781) );
  INVX0 U19625 ( .IN(n17891), .QN(n20553) );
  INVX0 U19626 ( .IN(n20623), .QN(n20611) );
  INVX0 U19627 ( .IN(n20554), .QN(n20536) );
  INVX0 U19628 ( .IN(n20554), .QN(n20537) );
  INVX0 U19629 ( .IN(n20554), .QN(n20538) );
  INVX0 U19630 ( .IN(n20654), .QN(n20638) );
  INVX0 U19631 ( .IN(n20622), .QN(n20605) );
  INVX0 U19632 ( .IN(n20588), .QN(n20572) );
  INVX0 U19633 ( .IN(n20655), .QN(n20639) );
  INVX0 U19634 ( .IN(n20623), .QN(n20606) );
  INVX0 U19635 ( .IN(n20589), .QN(n20573) );
  INVX0 U19636 ( .IN(n20654), .QN(n20640) );
  INVX0 U19637 ( .IN(n20622), .QN(n20607) );
  INVX0 U19638 ( .IN(n20588), .QN(n20574) );
  INVX0 U19639 ( .IN(n20654), .QN(n20641) );
  INVX0 U19640 ( .IN(n20622), .QN(n20608) );
  INVX0 U19641 ( .IN(n20588), .QN(n20575) );
  INVX0 U19642 ( .IN(n20654), .QN(n20642) );
  INVX0 U19643 ( .IN(n20623), .QN(n20609) );
  INVX0 U19644 ( .IN(n17909), .QN(n20576) );
  INVX0 U19645 ( .IN(n20623), .QN(n20610) );
  INVX0 U19646 ( .IN(n17909), .QN(n20577) );
  INVX0 U19647 ( .IN(n20655), .QN(n20643) );
  INVX0 U19648 ( .IN(n17881), .QN(n20612) );
  INVX0 U19649 ( .IN(n20589), .QN(n20578) );
  INVX0 U19650 ( .IN(n20656), .QN(n20649) );
  INVX0 U19651 ( .IN(n20653), .QN(n20651) );
  INVX0 U19652 ( .IN(n20624), .QN(n20619) );
  INVX0 U19653 ( .IN(n20590), .QN(n20585) );
  INVX0 U19654 ( .IN(n20655), .QN(n20644) );
  INVX0 U19655 ( .IN(n20589), .QN(n20579) );
  INVX0 U19656 ( .IN(n20655), .QN(n20645) );
  INVX0 U19657 ( .IN(n20622), .QN(n20613) );
  INVX0 U19658 ( .IN(n20623), .QN(n20614) );
  INVX0 U19659 ( .IN(n20588), .QN(n20580) );
  INVX0 U19660 ( .IN(n20656), .QN(n20646) );
  INVX0 U19661 ( .IN(n20624), .QN(n20615) );
  INVX0 U19662 ( .IN(n20590), .QN(n20581) );
  INVX0 U19663 ( .IN(n20656), .QN(n20647) );
  INVX0 U19664 ( .IN(n20624), .QN(n20616) );
  INVX0 U19665 ( .IN(n20590), .QN(n20582) );
  INVX0 U19666 ( .IN(n20656), .QN(n20648) );
  INVX0 U19667 ( .IN(n20624), .QN(n20617) );
  INVX0 U19668 ( .IN(n20590), .QN(n20583) );
  INVX0 U19669 ( .IN(n17892), .QN(n20421) );
  INVX0 U19670 ( .IN(n20491), .QN(n20478) );
  INVX0 U19671 ( .IN(n20422), .QN(n20404) );
  INVX0 U19672 ( .IN(n20422), .QN(n20405) );
  INVX0 U19673 ( .IN(n20422), .QN(n20406) );
  INVX0 U19674 ( .IN(n20522), .QN(n20506) );
  INVX0 U19675 ( .IN(n20490), .QN(n20473) );
  INVX0 U19676 ( .IN(n20456), .QN(n20440) );
  INVX0 U19677 ( .IN(n20523), .QN(n20507) );
  INVX0 U19678 ( .IN(n20491), .QN(n20474) );
  INVX0 U19679 ( .IN(n20457), .QN(n20441) );
  INVX0 U19680 ( .IN(n20522), .QN(n20508) );
  INVX0 U19681 ( .IN(n20490), .QN(n20475) );
  INVX0 U19682 ( .IN(n20456), .QN(n20442) );
  INVX0 U19683 ( .IN(n20522), .QN(n20509) );
  INVX0 U19684 ( .IN(n20490), .QN(n20476) );
  INVX0 U19685 ( .IN(n20456), .QN(n20443) );
  INVX0 U19686 ( .IN(n20522), .QN(n20510) );
  INVX0 U19687 ( .IN(n20492), .QN(n20477) );
  INVX0 U19688 ( .IN(n17910), .QN(n20444) );
  INVX0 U19689 ( .IN(n17910), .QN(n20445) );
  INVX0 U19690 ( .IN(n20523), .QN(n20511) );
  INVX0 U19691 ( .IN(n20491), .QN(n20479) );
  INVX0 U19692 ( .IN(n20457), .QN(n20446) );
  INVX0 U19693 ( .IN(n20524), .QN(n20517) );
  INVX0 U19694 ( .IN(n20489), .QN(n20486) );
  INVX0 U19695 ( .IN(n20521), .QN(n20519) );
  INVX0 U19696 ( .IN(n20458), .QN(n20453) );
  INVX0 U19697 ( .IN(n20523), .QN(n20512) );
  INVX0 U19698 ( .IN(n20491), .QN(n20480) );
  INVX0 U19699 ( .IN(n20457), .QN(n20447) );
  INVX0 U19700 ( .IN(n20523), .QN(n20513) );
  INVX0 U19701 ( .IN(n20491), .QN(n20481) );
  INVX0 U19702 ( .IN(n20490), .QN(n20482) );
  INVX0 U19703 ( .IN(n20456), .QN(n20448) );
  INVX0 U19704 ( .IN(n20524), .QN(n20514) );
  INVX0 U19705 ( .IN(n20492), .QN(n20483) );
  INVX0 U19706 ( .IN(n20458), .QN(n20449) );
  INVX0 U19707 ( .IN(n20524), .QN(n20515) );
  INVX0 U19708 ( .IN(n20492), .QN(n20484) );
  INVX0 U19709 ( .IN(n20458), .QN(n20450) );
  INVX0 U19710 ( .IN(n20524), .QN(n20516) );
  INVX0 U19711 ( .IN(n20492), .QN(n20485) );
  INVX0 U19712 ( .IN(n20458), .QN(n20451) );
  INVX0 U19713 ( .IN(n17893), .QN(n20289) );
  INVX0 U19714 ( .IN(n20290), .QN(n20272) );
  INVX0 U19715 ( .IN(n20290), .QN(n20273) );
  INVX0 U19716 ( .IN(n20290), .QN(n20274) );
  INVX0 U19717 ( .IN(n20390), .QN(n20374) );
  INVX0 U19718 ( .IN(n20357), .QN(n20341) );
  INVX0 U19719 ( .IN(n20324), .QN(n20308) );
  INVX0 U19720 ( .IN(n20391), .QN(n20375) );
  INVX0 U19721 ( .IN(n20358), .QN(n20342) );
  INVX0 U19722 ( .IN(n20325), .QN(n20309) );
  INVX0 U19723 ( .IN(n20390), .QN(n20376) );
  INVX0 U19724 ( .IN(n20357), .QN(n20343) );
  INVX0 U19725 ( .IN(n20324), .QN(n20310) );
  INVX0 U19726 ( .IN(n20390), .QN(n20377) );
  INVX0 U19727 ( .IN(n20357), .QN(n20344) );
  INVX0 U19728 ( .IN(n20324), .QN(n20311) );
  INVX0 U19729 ( .IN(n20390), .QN(n20378) );
  INVX0 U19730 ( .IN(n17912), .QN(n20345) );
  INVX0 U19731 ( .IN(n17911), .QN(n20312) );
  INVX0 U19732 ( .IN(n17912), .QN(n20346) );
  INVX0 U19733 ( .IN(n17911), .QN(n20313) );
  INVX0 U19734 ( .IN(n20391), .QN(n20379) );
  INVX0 U19735 ( .IN(n20358), .QN(n20347) );
  INVX0 U19736 ( .IN(n20325), .QN(n20314) );
  INVX0 U19737 ( .IN(n20392), .QN(n20385) );
  INVX0 U19738 ( .IN(n20389), .QN(n20387) );
  INVX0 U19739 ( .IN(n20359), .QN(n20354) );
  INVX0 U19740 ( .IN(n20326), .QN(n20321) );
  INVX0 U19741 ( .IN(n20391), .QN(n20380) );
  INVX0 U19742 ( .IN(n20358), .QN(n20348) );
  INVX0 U19743 ( .IN(n20325), .QN(n20315) );
  INVX0 U19744 ( .IN(n20391), .QN(n20381) );
  INVX0 U19745 ( .IN(n20357), .QN(n20349) );
  INVX0 U19746 ( .IN(n20324), .QN(n20316) );
  INVX0 U19747 ( .IN(n20392), .QN(n20382) );
  INVX0 U19748 ( .IN(n20359), .QN(n20350) );
  INVX0 U19749 ( .IN(n20326), .QN(n20317) );
  INVX0 U19750 ( .IN(n20392), .QN(n20383) );
  INVX0 U19751 ( .IN(n20359), .QN(n20351) );
  INVX0 U19752 ( .IN(n20326), .QN(n20318) );
  INVX0 U19753 ( .IN(n20392), .QN(n20384) );
  INVX0 U19754 ( .IN(n20359), .QN(n20352) );
  INVX0 U19755 ( .IN(n20326), .QN(n20319) );
  INVX0 U19756 ( .IN(n20162), .QN(n20157) );
  INVX0 U19757 ( .IN(n20158), .QN(n20140) );
  INVX0 U19758 ( .IN(n20158), .QN(n20141) );
  INVX0 U19759 ( .IN(n20158), .QN(n20142) );
  INVX0 U19760 ( .IN(n20258), .QN(n20242) );
  INVX0 U19761 ( .IN(n20225), .QN(n20209) );
  INVX0 U19762 ( .IN(n20192), .QN(n20176) );
  INVX0 U19763 ( .IN(n20259), .QN(n20243) );
  INVX0 U19764 ( .IN(n20226), .QN(n20210) );
  INVX0 U19765 ( .IN(n20193), .QN(n20177) );
  INVX0 U19766 ( .IN(n20258), .QN(n20244) );
  INVX0 U19767 ( .IN(n20225), .QN(n20211) );
  INVX0 U19768 ( .IN(n20192), .QN(n20178) );
  INVX0 U19769 ( .IN(n20258), .QN(n20245) );
  INVX0 U19770 ( .IN(n20225), .QN(n20212) );
  INVX0 U19771 ( .IN(n20192), .QN(n20179) );
  INVX0 U19772 ( .IN(n20258), .QN(n20246) );
  INVX0 U19773 ( .IN(n17914), .QN(n20213) );
  INVX0 U19774 ( .IN(n17913), .QN(n20180) );
  INVX0 U19775 ( .IN(n17914), .QN(n20214) );
  INVX0 U19776 ( .IN(n17913), .QN(n20181) );
  INVX0 U19777 ( .IN(n20259), .QN(n20247) );
  INVX0 U19778 ( .IN(n20226), .QN(n20215) );
  INVX0 U19779 ( .IN(n20193), .QN(n20182) );
  INVX0 U19780 ( .IN(n20261), .QN(n20253) );
  INVX0 U19781 ( .IN(n20162), .QN(n20155) );
  INVX0 U19782 ( .IN(n20260), .QN(n20255) );
  INVX0 U19783 ( .IN(n20227), .QN(n20222) );
  INVX0 U19784 ( .IN(n20194), .QN(n20189) );
  INVX0 U19785 ( .IN(n20259), .QN(n20248) );
  INVX0 U19786 ( .IN(n20226), .QN(n20216) );
  INVX0 U19787 ( .IN(n20193), .QN(n20183) );
  INVX0 U19788 ( .IN(n17932), .QN(n20249) );
  INVX0 U19789 ( .IN(n20225), .QN(n20217) );
  INVX0 U19790 ( .IN(n20192), .QN(n20184) );
  INVX0 U19791 ( .IN(n20260), .QN(n20250) );
  INVX0 U19792 ( .IN(n20227), .QN(n20218) );
  INVX0 U19793 ( .IN(n20194), .QN(n20185) );
  INVX0 U19794 ( .IN(n20260), .QN(n20251) );
  INVX0 U19795 ( .IN(n20227), .QN(n20219) );
  INVX0 U19796 ( .IN(n20194), .QN(n20186) );
  INVX0 U19797 ( .IN(n20260), .QN(n20252) );
  INVX0 U19798 ( .IN(n20227), .QN(n20220) );
  INVX0 U19799 ( .IN(n20194), .QN(n20187) );
  INVX0 U19800 ( .IN(n20031), .QN(n20026) );
  INVX0 U19801 ( .IN(n17921), .QN(n20113) );
  INVX0 U19802 ( .IN(n20074), .QN(n20082) );
  INVX0 U19803 ( .IN(n20062), .QN(n20051) );
  INVX0 U19804 ( .IN(n20027), .QN(n20009) );
  INVX0 U19805 ( .IN(n20027), .QN(n20010) );
  INVX0 U19806 ( .IN(n20027), .QN(n20011) );
  INVX0 U19807 ( .IN(n20127), .QN(n20110) );
  INVX0 U19808 ( .IN(n20094), .QN(n20078) );
  INVX0 U19809 ( .IN(n20061), .QN(n20045) );
  INVX0 U19810 ( .IN(n20126), .QN(n20111) );
  INVX0 U19811 ( .IN(n20096), .QN(n20079) );
  INVX0 U19812 ( .IN(n20063), .QN(n20046) );
  INVX0 U19813 ( .IN(n20126), .QN(n20112) );
  INVX0 U19814 ( .IN(n20094), .QN(n20080) );
  INVX0 U19815 ( .IN(n20061), .QN(n20047) );
  INVX0 U19816 ( .IN(n20094), .QN(n20081) );
  INVX0 U19817 ( .IN(n20061), .QN(n20048) );
  INVX0 U19818 ( .IN(n20062), .QN(n20049) );
  INVX0 U19819 ( .IN(n20062), .QN(n20050) );
  INVX0 U19820 ( .IN(n20126), .QN(n20114) );
  INVX0 U19821 ( .IN(n20093), .QN(n20083) );
  INVX0 U19822 ( .IN(n20063), .QN(n20052) );
  INVX0 U19823 ( .IN(n20128), .QN(n20122) );
  INVX0 U19824 ( .IN(n20096), .QN(n20090) );
  INVX0 U19825 ( .IN(n17915), .QN(n20059) );
  INVX0 U19826 ( .IN(n20031), .QN(n20025) );
  INVX0 U19827 ( .IN(n20125), .QN(n20123) );
  INVX0 U19828 ( .IN(n20096), .QN(n20092) );
  INVX0 U19829 ( .IN(n20126), .QN(n20115) );
  INVX0 U19830 ( .IN(n20063), .QN(n20053) );
  INVX0 U19831 ( .IN(n20127), .QN(n20116) );
  INVX0 U19832 ( .IN(n20096), .QN(n20084) );
  INVX0 U19833 ( .IN(n20064), .QN(n20054) );
  INVX0 U19834 ( .IN(n20127), .QN(n20117) );
  INVX0 U19835 ( .IN(n20096), .QN(n20085) );
  INVX0 U19836 ( .IN(n20064), .QN(n20055) );
  INVX0 U19837 ( .IN(n20127), .QN(n20118) );
  INVX0 U19838 ( .IN(n20064), .QN(n20056) );
  INVX0 U19839 ( .IN(n20128), .QN(n20119) );
  INVX0 U19840 ( .IN(n20095), .QN(n20086) );
  INVX0 U19841 ( .IN(n17915), .QN(n20057) );
  INVX0 U19842 ( .IN(n20128), .QN(n20120) );
  INVX0 U19843 ( .IN(n20095), .QN(n20087) );
  INVX0 U19844 ( .IN(n20060), .QN(n20058) );
  INVX0 U19845 ( .IN(n20128), .QN(n20121) );
  INVX0 U19846 ( .IN(n20095), .QN(n20088) );
  INVX0 U19847 ( .IN(n20096), .QN(n20089) );
  INVX0 U19848 ( .IN(n19900), .QN(n19895) );
  INVX0 U19849 ( .IN(n17922), .QN(n19982) );
  INVX0 U19850 ( .IN(n19962), .QN(n19951) );
  INVX0 U19851 ( .IN(n19931), .QN(n19920) );
  INVX0 U19852 ( .IN(n19896), .QN(n19878) );
  INVX0 U19853 ( .IN(n19896), .QN(n19879) );
  INVX0 U19854 ( .IN(n19896), .QN(n19880) );
  INVX0 U19855 ( .IN(n19996), .QN(n19979) );
  INVX0 U19856 ( .IN(n19963), .QN(n19947) );
  INVX0 U19857 ( .IN(n19930), .QN(n19914) );
  INVX0 U19858 ( .IN(n19995), .QN(n19980) );
  INVX0 U19859 ( .IN(n19964), .QN(n19948) );
  INVX0 U19860 ( .IN(n19932), .QN(n19915) );
  INVX0 U19861 ( .IN(n19995), .QN(n19981) );
  INVX0 U19862 ( .IN(n19963), .QN(n19949) );
  INVX0 U19863 ( .IN(n19930), .QN(n19916) );
  INVX0 U19864 ( .IN(n19963), .QN(n19950) );
  INVX0 U19865 ( .IN(n19930), .QN(n19917) );
  INVX0 U19866 ( .IN(n19931), .QN(n19918) );
  INVX0 U19867 ( .IN(n19931), .QN(n19919) );
  INVX0 U19868 ( .IN(n19995), .QN(n19983) );
  INVX0 U19869 ( .IN(n19964), .QN(n19952) );
  INVX0 U19870 ( .IN(n19932), .QN(n19921) );
  INVX0 U19871 ( .IN(n19997), .QN(n19991) );
  INVX0 U19872 ( .IN(n19962), .QN(n19958) );
  INVX0 U19873 ( .IN(n17916), .QN(n19928) );
  INVX0 U19874 ( .IN(n19900), .QN(n19894) );
  INVX0 U19875 ( .IN(n19994), .QN(n19992) );
  INVX0 U19876 ( .IN(n19963), .QN(n19960) );
  INVX0 U19877 ( .IN(n19995), .QN(n19984) );
  INVX0 U19878 ( .IN(n19964), .QN(n19953) );
  INVX0 U19879 ( .IN(n19932), .QN(n19922) );
  INVX0 U19880 ( .IN(n19996), .QN(n19985) );
  INVX0 U19881 ( .IN(n19965), .QN(n19954) );
  INVX0 U19882 ( .IN(n19933), .QN(n19923) );
  INVX0 U19883 ( .IN(n19996), .QN(n19986) );
  INVX0 U19884 ( .IN(n19965), .QN(n19955) );
  INVX0 U19885 ( .IN(n19933), .QN(n19924) );
  INVX0 U19886 ( .IN(n19996), .QN(n19987) );
  INVX0 U19887 ( .IN(n19965), .QN(n19956) );
  INVX0 U19888 ( .IN(n19933), .QN(n19925) );
  INVX0 U19889 ( .IN(n19997), .QN(n19988) );
  INVX0 U19890 ( .IN(n19964), .QN(n19957) );
  INVX0 U19891 ( .IN(n17916), .QN(n19926) );
  INVX0 U19892 ( .IN(n19997), .QN(n19989) );
  INVX0 U19893 ( .IN(n19929), .QN(n19927) );
  INVX0 U19894 ( .IN(n19997), .QN(n19990) );
  INVX0 U19895 ( .IN(n19768), .QN(n19763) );
  INVX0 U19896 ( .IN(n17923), .QN(n19851) );
  INVX0 U19897 ( .IN(n19831), .QN(n19819) );
  INVX0 U19898 ( .IN(n19799), .QN(n19788) );
  INVX0 U19899 ( .IN(n19764), .QN(n19746) );
  INVX0 U19900 ( .IN(n19764), .QN(n19747) );
  INVX0 U19901 ( .IN(n19764), .QN(n19748) );
  INVX0 U19902 ( .IN(n19865), .QN(n19848) );
  INVX0 U19903 ( .IN(n19830), .QN(n19813) );
  INVX0 U19904 ( .IN(n19798), .QN(n19782) );
  INVX0 U19905 ( .IN(n19864), .QN(n19849) );
  INVX0 U19906 ( .IN(n19832), .QN(n19814) );
  INVX0 U19907 ( .IN(n19800), .QN(n19783) );
  INVX0 U19908 ( .IN(n19864), .QN(n19850) );
  INVX0 U19909 ( .IN(n19830), .QN(n19815) );
  INVX0 U19910 ( .IN(n19798), .QN(n19784) );
  INVX0 U19911 ( .IN(n19830), .QN(n19816) );
  INVX0 U19912 ( .IN(n19798), .QN(n19785) );
  INVX0 U19913 ( .IN(n19831), .QN(n19817) );
  INVX0 U19914 ( .IN(n19799), .QN(n19786) );
  INVX0 U19915 ( .IN(n19831), .QN(n19818) );
  INVX0 U19916 ( .IN(n19799), .QN(n19787) );
  INVX0 U19917 ( .IN(n19864), .QN(n19852) );
  INVX0 U19918 ( .IN(n19832), .QN(n19820) );
  INVX0 U19919 ( .IN(n19800), .QN(n19789) );
  INVX0 U19920 ( .IN(n19866), .QN(n19860) );
  INVX0 U19921 ( .IN(n19834), .QN(n19827) );
  INVX0 U19922 ( .IN(n17917), .QN(n19796) );
  INVX0 U19923 ( .IN(n19768), .QN(n19762) );
  INVX0 U19924 ( .IN(n19863), .QN(n19861) );
  INVX0 U19925 ( .IN(n19834), .QN(n19829) );
  INVX0 U19926 ( .IN(n19864), .QN(n19853) );
  INVX0 U19927 ( .IN(n19800), .QN(n19790) );
  INVX0 U19928 ( .IN(n19865), .QN(n19854) );
  INVX0 U19929 ( .IN(n19830), .QN(n19821) );
  INVX0 U19930 ( .IN(n19801), .QN(n19791) );
  INVX0 U19931 ( .IN(n19865), .QN(n19855) );
  INVX0 U19932 ( .IN(n19831), .QN(n19822) );
  INVX0 U19933 ( .IN(n19801), .QN(n19792) );
  INVX0 U19934 ( .IN(n19865), .QN(n19856) );
  INVX0 U19935 ( .IN(n19801), .QN(n19793) );
  INVX0 U19936 ( .IN(n19866), .QN(n19857) );
  INVX0 U19937 ( .IN(n19833), .QN(n19823) );
  INVX0 U19938 ( .IN(n17917), .QN(n19794) );
  INVX0 U19939 ( .IN(n19866), .QN(n19858) );
  INVX0 U19940 ( .IN(n19833), .QN(n19824) );
  INVX0 U19941 ( .IN(n19797), .QN(n19795) );
  INVX0 U19942 ( .IN(n19866), .QN(n19859) );
  INVX0 U19943 ( .IN(n19833), .QN(n19825) );
  INVX0 U19944 ( .IN(n19834), .QN(n19826) );
  INVX0 U19945 ( .IN(n18844), .QN(n18839) );
  INVX0 U19946 ( .IN(n17924), .QN(n18927) );
  INVX0 U19947 ( .IN(n18907), .QN(n18895) );
  INVX0 U19948 ( .IN(n18875), .QN(n18864) );
  INVX0 U19949 ( .IN(n18840), .QN(n18822) );
  INVX0 U19950 ( .IN(n18840), .QN(n18823) );
  INVX0 U19951 ( .IN(n18840), .QN(n18824) );
  INVX0 U19952 ( .IN(n18941), .QN(n18924) );
  INVX0 U19953 ( .IN(n18906), .QN(n18889) );
  INVX0 U19954 ( .IN(n18874), .QN(n18858) );
  INVX0 U19955 ( .IN(n18940), .QN(n18925) );
  INVX0 U19956 ( .IN(n18908), .QN(n18890) );
  INVX0 U19957 ( .IN(n18876), .QN(n18859) );
  INVX0 U19958 ( .IN(n18940), .QN(n18926) );
  INVX0 U19959 ( .IN(n18906), .QN(n18891) );
  INVX0 U19960 ( .IN(n18874), .QN(n18860) );
  INVX0 U19961 ( .IN(n18906), .QN(n18892) );
  INVX0 U19962 ( .IN(n18874), .QN(n18861) );
  INVX0 U19963 ( .IN(n18907), .QN(n18893) );
  INVX0 U19964 ( .IN(n18875), .QN(n18862) );
  INVX0 U19965 ( .IN(n18907), .QN(n18894) );
  INVX0 U19966 ( .IN(n18875), .QN(n18863) );
  INVX0 U19967 ( .IN(n18940), .QN(n18928) );
  INVX0 U19968 ( .IN(n18908), .QN(n18896) );
  INVX0 U19969 ( .IN(n18876), .QN(n18865) );
  INVX0 U19970 ( .IN(n18942), .QN(n18936) );
  INVX0 U19971 ( .IN(n18910), .QN(n18903) );
  INVX0 U19972 ( .IN(n17918), .QN(n18872) );
  INVX0 U19973 ( .IN(n18844), .QN(n18838) );
  INVX0 U19974 ( .IN(n18939), .QN(n18937) );
  INVX0 U19975 ( .IN(n18910), .QN(n18905) );
  INVX0 U19976 ( .IN(n18940), .QN(n18929) );
  INVX0 U19977 ( .IN(n18876), .QN(n18866) );
  INVX0 U19978 ( .IN(n18941), .QN(n18930) );
  INVX0 U19979 ( .IN(n18906), .QN(n18897) );
  INVX0 U19980 ( .IN(n18877), .QN(n18867) );
  INVX0 U19981 ( .IN(n18941), .QN(n18931) );
  INVX0 U19982 ( .IN(n18907), .QN(n18898) );
  INVX0 U19983 ( .IN(n18877), .QN(n18868) );
  INVX0 U19984 ( .IN(n18941), .QN(n18932) );
  INVX0 U19985 ( .IN(n18877), .QN(n18869) );
  INVX0 U19986 ( .IN(n18942), .QN(n18933) );
  INVX0 U19987 ( .IN(n18909), .QN(n18899) );
  INVX0 U19988 ( .IN(n17918), .QN(n18870) );
  INVX0 U19989 ( .IN(n18942), .QN(n18934) );
  INVX0 U19990 ( .IN(n18909), .QN(n18900) );
  INVX0 U19991 ( .IN(n18873), .QN(n18871) );
  INVX0 U19992 ( .IN(n18942), .QN(n18935) );
  INVX0 U19993 ( .IN(n18909), .QN(n18901) );
  INVX0 U19994 ( .IN(n18910), .QN(n18902) );
  INVX0 U19995 ( .IN(n21052), .QN(n21016) );
  INVX0 U19996 ( .IN(n21053), .QN(n21015) );
  INVX0 U19997 ( .IN(n21056), .QN(n21008) );
  INVX0 U19998 ( .IN(n21053), .QN(n21014) );
  INVX0 U19999 ( .IN(n21054), .QN(n21013) );
  INVX0 U20000 ( .IN(n21057), .QN(n21007) );
  INVX0 U20001 ( .IN(n21057), .QN(n21006) );
  INVX0 U20002 ( .IN(n21054), .QN(n21012) );
  INVX0 U20003 ( .IN(n21055), .QN(n21011) );
  INVX0 U20004 ( .IN(n21058), .QN(n21005) );
  INVX0 U20005 ( .IN(n21058), .QN(n21004) );
  INVX0 U20006 ( .IN(n21055), .QN(n21010) );
  INVX0 U20007 ( .IN(n21056), .QN(n21009) );
  INVX0 U20008 ( .IN(n21059), .QN(n21003) );
  INVX0 U20009 ( .IN(n21059), .QN(n21002) );
  INVX0 U20010 ( .IN(n21052), .QN(n21017) );
  INVX0 U20011 ( .IN(n20987), .QN(n20871) );
  INVX0 U20012 ( .IN(n20988), .QN(n20872) );
  INVX0 U20013 ( .IN(n20989), .QN(n20873) );
  INVX0 U20014 ( .IN(n20986), .QN(n20985) );
  INVX0 U20015 ( .IN(n21046), .QN(n21023) );
  INVX0 U20016 ( .IN(n21051), .QN(n21018) );
  INVX0 U20017 ( .IN(n21051), .QN(n21019) );
  INVX0 U20018 ( .IN(n21049), .QN(n21020) );
  INVX0 U20019 ( .IN(n21048), .QN(n21022) );
  INVX0 U20020 ( .IN(n21050), .QN(n21024) );
  INVX0 U20021 ( .IN(n21047), .QN(n21025) );
  INVX0 U20022 ( .IN(n21050), .QN(n21026) );
  INVX0 U20023 ( .IN(n21051), .QN(n21027) );
  INVX0 U20024 ( .IN(n21078), .QN(n21028) );
  INVX0 U20025 ( .IN(n21049), .QN(n21029) );
  INVX0 U20026 ( .IN(n21049), .QN(n21030) );
  INVX0 U20027 ( .IN(n21048), .QN(n21031) );
  INVX0 U20028 ( .IN(n21048), .QN(n21032) );
  INVX0 U20029 ( .IN(n21047), .QN(n21033) );
  INVX0 U20030 ( .IN(n21047), .QN(n21034) );
  INVX0 U20031 ( .IN(n21046), .QN(n21035) );
  INVX0 U20032 ( .IN(n21046), .QN(n21036) );
  INVX0 U20033 ( .IN(n21049), .QN(n21037) );
  INVX0 U20034 ( .IN(n21051), .QN(n21038) );
  INVX0 U20035 ( .IN(n21078), .QN(n21039) );
  INVX0 U20036 ( .IN(n21045), .QN(n21040) );
  INVX0 U20037 ( .IN(n21045), .QN(n21041) );
  INVX0 U20038 ( .IN(n21045), .QN(n21042) );
  INVX0 U20039 ( .IN(n21078), .QN(n21043) );
  INVX0 U20040 ( .IN(n21045), .QN(n21044) );
  INVX0 U20041 ( .IN(n21048), .QN(n21021) );
  INVX0 U20042 ( .IN(n17780), .QN(n18818) );
  INVX0 U20043 ( .IN(n17780), .QN(n18819) );
  INVX0 U20044 ( .IN(n17780), .QN(n18817) );
  INVX0 U20045 ( .IN(n19613), .QN(n19633) );
  INVX0 U20046 ( .IN(n19613), .QN(n19632) );
  INVX0 U20047 ( .IN(n19732), .QN(n19718) );
  INVX0 U20048 ( .IN(n19699), .QN(n19685) );
  INVX0 U20049 ( .IN(n19666), .QN(n19652) );
  INVX0 U20050 ( .IN(n19732), .QN(n19719) );
  INVX0 U20051 ( .IN(n19699), .QN(n19686) );
  INVX0 U20052 ( .IN(n19666), .QN(n19653) );
  INVX0 U20053 ( .IN(n19615), .QN(n19636) );
  INVX0 U20054 ( .IN(n19616), .QN(n19615) );
  NAND2X0 U20055 ( .IN1(n17785), .IN2(n19731), .QN(n14881) );
  NAND2X0 U20056 ( .IN1(n17788), .IN2(n19698), .QN(n15491) );
  NAND2X0 U20057 ( .IN1(n17786), .IN2(n19665), .QN(n16101) );
  NAND2X0 U20058 ( .IN1(n17787), .IN2(n19632), .QN(n16711) );
  INVX0 U20059 ( .IN(n19680), .QN(n19700) );
  INVX0 U20060 ( .IN(n19647), .QN(n19667) );
  INVX0 U20061 ( .IN(n19713), .QN(n19733) );
  INVX0 U20062 ( .IN(n19617), .QN(n19614) );
  INVX0 U20063 ( .IN(n18295), .QN(n18395) );
  INVX0 U20064 ( .IN(n18286), .QN(n18423) );
  INVX0 U20065 ( .IN(n18289), .QN(n18399) );
  INVX0 U20066 ( .IN(n18287), .QN(n18427) );
  INVX0 U20067 ( .IN(n18290), .QN(n18375) );
  INVX0 U20068 ( .IN(n18298), .QN(n18335) );
  INVX0 U20069 ( .IN(n18292), .QN(n18415) );
  INVX0 U20070 ( .IN(n18294), .QN(n18379) );
  INVX0 U20071 ( .IN(n18299), .QN(n18403) );
  INVX0 U20072 ( .IN(n18293), .QN(n18419) );
  INVX0 U20073 ( .IN(n18288), .QN(n18383) );
  INVX0 U20074 ( .IN(n18300), .QN(n18407) );
  INVX0 U20075 ( .IN(n18301), .QN(n18411) );
  INVX0 U20076 ( .IN(n18297), .QN(n18386) );
  INVX0 U20077 ( .IN(n18291), .QN(n18390) );
  INVX0 U20078 ( .IN(n18295), .QN(n18394) );
  INVX0 U20079 ( .IN(n18289), .QN(n18398) );
  INVX0 U20080 ( .IN(n18286), .QN(n18422) );
  INVX0 U20081 ( .IN(n18296), .QN(n18370) );
  INVX0 U20082 ( .IN(n18287), .QN(n18426) );
  INVX0 U20083 ( .IN(n18290), .QN(n18374) );
  INVX0 U20084 ( .IN(n18292), .QN(n18414) );
  INVX0 U20085 ( .IN(n18294), .QN(n18378) );
  INVX0 U20086 ( .IN(n18298), .QN(n18334) );
  INVX0 U20087 ( .IN(n18293), .QN(n18418) );
  INVX0 U20088 ( .IN(n18288), .QN(n18382) );
  INVX0 U20089 ( .IN(n18299), .QN(n18402) );
  INVX0 U20090 ( .IN(n18300), .QN(n18406) );
  INVX0 U20091 ( .IN(n18301), .QN(n18410) );
  INVX0 U20092 ( .IN(n17781), .QN(n18809) );
  INVX0 U20093 ( .IN(n17785), .QN(n18761) );
  INVX0 U20094 ( .IN(n17782), .QN(n18713) );
  INVX0 U20095 ( .IN(n17788), .QN(n18665) );
  INVX0 U20096 ( .IN(n17783), .QN(n18617) );
  INVX0 U20097 ( .IN(n17786), .QN(n18569) );
  INVX0 U20098 ( .IN(n17784), .QN(n18521) );
  INVX0 U20099 ( .IN(n17787), .QN(n18473) );
  INVX0 U20100 ( .IN(n17781), .QN(n18810) );
  INVX0 U20101 ( .IN(n17781), .QN(n18811) );
  INVX0 U20102 ( .IN(n17785), .QN(n18762) );
  INVX0 U20103 ( .IN(n17785), .QN(n18763) );
  INVX0 U20104 ( .IN(n17782), .QN(n18714) );
  INVX0 U20105 ( .IN(n17782), .QN(n18715) );
  INVX0 U20106 ( .IN(n17788), .QN(n18666) );
  INVX0 U20107 ( .IN(n17788), .QN(n18667) );
  INVX0 U20108 ( .IN(n17783), .QN(n18618) );
  INVX0 U20109 ( .IN(n17783), .QN(n18619) );
  INVX0 U20110 ( .IN(n17786), .QN(n18570) );
  INVX0 U20111 ( .IN(n17786), .QN(n18571) );
  INVX0 U20112 ( .IN(n17784), .QN(n18522) );
  INVX0 U20113 ( .IN(n17784), .QN(n18523) );
  INVX0 U20114 ( .IN(n17787), .QN(n18474) );
  INVX0 U20115 ( .IN(n17787), .QN(n18475) );
  INVX0 U20116 ( .IN(n20807), .QN(n20803) );
  INVX0 U20117 ( .IN(n20807), .QN(n20799) );
  INVX0 U20118 ( .IN(n20807), .QN(n20800) );
  INVX0 U20119 ( .IN(n20807), .QN(n20801) );
  INVX0 U20120 ( .IN(n20807), .QN(n20802) );
  INVX0 U20121 ( .IN(n20807), .QN(n20806) );
  INVX0 U20122 ( .IN(n20807), .QN(n20804) );
  INVX0 U20123 ( .IN(n20807), .QN(n20805) );
  INVX0 U20124 ( .IN(n21067), .QN(n20987) );
  INVX0 U20125 ( .IN(n21066), .QN(n20989) );
  INVX0 U20126 ( .IN(n21066), .QN(n20988) );
  INVX0 U20127 ( .IN(n21067), .QN(n20986) );
  INVX0 U20128 ( .IN(n19730), .QN(n19734) );
  INVX0 U20129 ( .IN(n19697), .QN(n19701) );
  INVX0 U20130 ( .IN(n19664), .QN(n19668) );
  INVX0 U20131 ( .IN(n19481), .QN(n19500) );
  INVX0 U20132 ( .IN(n19591), .QN(n19600) );
  INVX0 U20133 ( .IN(n19547), .QN(n19568) );
  INVX0 U20134 ( .IN(n19514), .QN(n19534) );
  INVX0 U20135 ( .IN(n19580), .QN(n19601) );
  INVX0 U20136 ( .IN(n19547), .QN(n19569) );
  INVX0 U20137 ( .IN(n19514), .QN(n19535) );
  INVX0 U20138 ( .IN(n19580), .QN(n19602) );
  INVX0 U20139 ( .IN(n7358), .QN(n19570) );
  INVX0 U20140 ( .IN(n19514), .QN(n19536) );
  INVX0 U20141 ( .IN(n19349), .QN(n19368) );
  INVX0 U20142 ( .IN(n19415), .QN(n19435) );
  INVX0 U20143 ( .IN(n19382), .QN(n19402) );
  INVX0 U20144 ( .IN(n19448), .QN(n19468) );
  INVX0 U20145 ( .IN(n19415), .QN(n19436) );
  INVX0 U20146 ( .IN(n19382), .QN(n19403) );
  INVX0 U20147 ( .IN(n19448), .QN(n19469) );
  INVX0 U20148 ( .IN(n19448), .QN(n19470) );
  INVX0 U20149 ( .IN(n19415), .QN(n19437) );
  INVX0 U20150 ( .IN(n19382), .QN(n19404) );
  INVX0 U20151 ( .IN(n19217), .QN(n19236) );
  INVX0 U20152 ( .IN(n19283), .QN(n19303) );
  INVX0 U20153 ( .IN(n19250), .QN(n19270) );
  INVX0 U20154 ( .IN(n19316), .QN(n19336) );
  INVX0 U20155 ( .IN(n19283), .QN(n19304) );
  INVX0 U20156 ( .IN(n19250), .QN(n19271) );
  INVX0 U20157 ( .IN(n19316), .QN(n19337) );
  INVX0 U20158 ( .IN(n19316), .QN(n19338) );
  INVX0 U20159 ( .IN(n19283), .QN(n19305) );
  INVX0 U20160 ( .IN(n19250), .QN(n19272) );
  INVX0 U20161 ( .IN(n19085), .QN(n19104) );
  INVX0 U20162 ( .IN(n19151), .QN(n19171) );
  INVX0 U20163 ( .IN(n19118), .QN(n19138) );
  INVX0 U20164 ( .IN(n19151), .QN(n19172) );
  INVX0 U20165 ( .IN(n19184), .QN(n19204) );
  INVX0 U20166 ( .IN(n19151), .QN(n19173) );
  INVX0 U20167 ( .IN(n19118), .QN(n19139) );
  INVX0 U20168 ( .IN(n19184), .QN(n19205) );
  INVX0 U20169 ( .IN(n19184), .QN(n19206) );
  INVX0 U20170 ( .IN(n19118), .QN(n19140) );
  INVX0 U20171 ( .IN(n18953), .QN(n18972) );
  INVX0 U20172 ( .IN(n19019), .QN(n19038) );
  INVX0 U20173 ( .IN(n18986), .QN(n19006) );
  INVX0 U20174 ( .IN(n19019), .QN(n19039) );
  INVX0 U20175 ( .IN(n18986), .QN(n19007) );
  INVX0 U20176 ( .IN(n19052), .QN(n19072) );
  INVX0 U20177 ( .IN(n19019), .QN(n19040) );
  INVX0 U20178 ( .IN(n18986), .QN(n19008) );
  INVX0 U20179 ( .IN(n19052), .QN(n19073) );
  INVX0 U20180 ( .IN(n18986), .QN(n19009) );
  INVX0 U20181 ( .IN(n19052), .QN(n19074) );
  INVX0 U20182 ( .IN(n19019), .QN(n19041) );
  INVX0 U20183 ( .IN(n19019), .QN(n19042) );
  INVX0 U20184 ( .IN(n20667), .QN(n20686) );
  INVX0 U20185 ( .IN(n20733), .QN(n20753) );
  INVX0 U20186 ( .IN(n20700), .QN(n20720) );
  INVX0 U20187 ( .IN(n20733), .QN(n20754) );
  INVX0 U20188 ( .IN(n20700), .QN(n20721) );
  INVX0 U20189 ( .IN(n20766), .QN(n20786) );
  INVX0 U20190 ( .IN(n20733), .QN(n20755) );
  INVX0 U20191 ( .IN(n20700), .QN(n20722) );
  INVX0 U20192 ( .IN(n20766), .QN(n20787) );
  INVX0 U20193 ( .IN(n20700), .QN(n20723) );
  INVX0 U20194 ( .IN(n20766), .QN(n20788) );
  INVX0 U20195 ( .IN(n20553), .QN(n20554) );
  INVX0 U20196 ( .IN(n20634), .QN(n20654) );
  INVX0 U20197 ( .IN(n20601), .QN(n20622) );
  INVX0 U20198 ( .IN(n20568), .QN(n20588) );
  INVX0 U20199 ( .IN(n20601), .QN(n20623) );
  INVX0 U20200 ( .IN(n20634), .QN(n20655) );
  INVX0 U20201 ( .IN(n20568), .QN(n20589) );
  INVX0 U20202 ( .IN(n20634), .QN(n20656) );
  INVX0 U20203 ( .IN(n20601), .QN(n20624) );
  INVX0 U20204 ( .IN(n20568), .QN(n20590) );
  INVX0 U20205 ( .IN(n20421), .QN(n20422) );
  INVX0 U20206 ( .IN(n20502), .QN(n20522) );
  INVX0 U20207 ( .IN(n20469), .QN(n20490) );
  INVX0 U20208 ( .IN(n20436), .QN(n20456) );
  INVX0 U20209 ( .IN(n20502), .QN(n20523) );
  INVX0 U20210 ( .IN(n20469), .QN(n20491) );
  INVX0 U20211 ( .IN(n20436), .QN(n20457) );
  INVX0 U20212 ( .IN(n20502), .QN(n20524) );
  INVX0 U20213 ( .IN(n20469), .QN(n20492) );
  INVX0 U20214 ( .IN(n20436), .QN(n20458) );
  INVX0 U20215 ( .IN(n20289), .QN(n20290) );
  INVX0 U20216 ( .IN(n20370), .QN(n20390) );
  INVX0 U20217 ( .IN(n20337), .QN(n20357) );
  INVX0 U20218 ( .IN(n20304), .QN(n20324) );
  INVX0 U20219 ( .IN(n20370), .QN(n20391) );
  INVX0 U20220 ( .IN(n20337), .QN(n20358) );
  INVX0 U20221 ( .IN(n20304), .QN(n20325) );
  INVX0 U20222 ( .IN(n20370), .QN(n20392) );
  INVX0 U20223 ( .IN(n20337), .QN(n20359) );
  INVX0 U20224 ( .IN(n20304), .QN(n20326) );
  INVX0 U20225 ( .IN(n20139), .QN(n20158) );
  INVX0 U20226 ( .IN(n20249), .QN(n20258) );
  INVX0 U20227 ( .IN(n20205), .QN(n20225) );
  INVX0 U20228 ( .IN(n20172), .QN(n20192) );
  INVX0 U20229 ( .IN(n20238), .QN(n20259) );
  INVX0 U20230 ( .IN(n20205), .QN(n20226) );
  INVX0 U20231 ( .IN(n20172), .QN(n20193) );
  INVX0 U20232 ( .IN(n20238), .QN(n20260) );
  INVX0 U20233 ( .IN(n20205), .QN(n20227) );
  INVX0 U20234 ( .IN(n20172), .QN(n20194) );
  INVX0 U20235 ( .IN(n20008), .QN(n20027) );
  INVX0 U20236 ( .IN(n6286), .QN(n20094) );
  INVX0 U20237 ( .IN(n20041), .QN(n20061) );
  INVX0 U20238 ( .IN(n20041), .QN(n20062) );
  INVX0 U20239 ( .IN(n20106), .QN(n20126) );
  INVX0 U20240 ( .IN(n20041), .QN(n20063) );
  INVX0 U20241 ( .IN(n20106), .QN(n20127) );
  INVX0 U20242 ( .IN(n20041), .QN(n20064) );
  INVX0 U20243 ( .IN(n20106), .QN(n20128) );
  INVX0 U20244 ( .IN(n6286), .QN(n20095) );
  INVX0 U20245 ( .IN(n6286), .QN(n20096) );
  INVX0 U20246 ( .IN(n19877), .QN(n19896) );
  INVX0 U20247 ( .IN(n19943), .QN(n19963) );
  INVX0 U20248 ( .IN(n19910), .QN(n19930) );
  INVX0 U20249 ( .IN(n19910), .QN(n19931) );
  INVX0 U20250 ( .IN(n19975), .QN(n19995) );
  INVX0 U20251 ( .IN(n19943), .QN(n19964) );
  INVX0 U20252 ( .IN(n19910), .QN(n19932) );
  INVX0 U20253 ( .IN(n19975), .QN(n19996) );
  INVX0 U20254 ( .IN(n19943), .QN(n19965) );
  INVX0 U20255 ( .IN(n19910), .QN(n19933) );
  INVX0 U20256 ( .IN(n19975), .QN(n19997) );
  INVX0 U20257 ( .IN(n19745), .QN(n19764) );
  INVX0 U20258 ( .IN(n19811), .QN(n19830) );
  INVX0 U20259 ( .IN(n19778), .QN(n19798) );
  INVX0 U20260 ( .IN(n19811), .QN(n19831) );
  INVX0 U20261 ( .IN(n19778), .QN(n19799) );
  INVX0 U20262 ( .IN(n19844), .QN(n19864) );
  INVX0 U20263 ( .IN(n19811), .QN(n19832) );
  INVX0 U20264 ( .IN(n19778), .QN(n19800) );
  INVX0 U20265 ( .IN(n19844), .QN(n19865) );
  INVX0 U20266 ( .IN(n19778), .QN(n19801) );
  INVX0 U20267 ( .IN(n19844), .QN(n19866) );
  INVX0 U20268 ( .IN(n19811), .QN(n19833) );
  INVX0 U20269 ( .IN(n19811), .QN(n19834) );
  INVX0 U20270 ( .IN(n18821), .QN(n18840) );
  INVX0 U20271 ( .IN(n18887), .QN(n18906) );
  INVX0 U20272 ( .IN(n18854), .QN(n18874) );
  INVX0 U20273 ( .IN(n18887), .QN(n18907) );
  INVX0 U20274 ( .IN(n18854), .QN(n18875) );
  INVX0 U20275 ( .IN(n18920), .QN(n18940) );
  INVX0 U20276 ( .IN(n18887), .QN(n18908) );
  INVX0 U20277 ( .IN(n18854), .QN(n18876) );
  INVX0 U20278 ( .IN(n18920), .QN(n18941) );
  INVX0 U20279 ( .IN(n18854), .QN(n18877) );
  INVX0 U20280 ( .IN(n18920), .QN(n18942) );
  INVX0 U20281 ( .IN(n18887), .QN(n18909) );
  INVX0 U20282 ( .IN(n18887), .QN(n18910) );
  INVX0 U20283 ( .IN(n19732), .QN(n19721) );
  INVX0 U20284 ( .IN(n19699), .QN(n19688) );
  INVX0 U20285 ( .IN(n19666), .QN(n19655) );
  INVX0 U20286 ( .IN(n19731), .QN(n19730) );
  INVX0 U20287 ( .IN(n19698), .QN(n19697) );
  INVX0 U20288 ( .IN(n19665), .QN(n19664) );
  INVX0 U20289 ( .IN(n19603), .QN(n19598) );
  INVX0 U20290 ( .IN(n19567), .QN(n19566) );
  INVX0 U20291 ( .IN(n19537), .QN(n19532) );
  INVX0 U20292 ( .IN(n19599), .QN(n19581) );
  INVX0 U20293 ( .IN(n19567), .QN(n19548) );
  INVX0 U20294 ( .IN(n19533), .QN(n19515) );
  INVX0 U20295 ( .IN(n19599), .QN(n19582) );
  INVX0 U20296 ( .IN(n19567), .QN(n19549) );
  INVX0 U20297 ( .IN(n19533), .QN(n19516) );
  INVX0 U20298 ( .IN(n19599), .QN(n19583) );
  INVX0 U20299 ( .IN(n19567), .QN(n19550) );
  INVX0 U20300 ( .IN(n19533), .QN(n19517) );
  INVX0 U20301 ( .IN(n19603), .QN(n19596) );
  INVX0 U20302 ( .IN(n19570), .QN(n19564) );
  INVX0 U20303 ( .IN(n19537), .QN(n19530) );
  INVX0 U20304 ( .IN(n19471), .QN(n19466) );
  INVX0 U20305 ( .IN(n19438), .QN(n19433) );
  INVX0 U20306 ( .IN(n19405), .QN(n19400) );
  INVX0 U20307 ( .IN(n19467), .QN(n19449) );
  INVX0 U20308 ( .IN(n19434), .QN(n19416) );
  INVX0 U20309 ( .IN(n19401), .QN(n19383) );
  INVX0 U20310 ( .IN(n19467), .QN(n19450) );
  INVX0 U20311 ( .IN(n19434), .QN(n19417) );
  INVX0 U20312 ( .IN(n19401), .QN(n19384) );
  INVX0 U20313 ( .IN(n19467), .QN(n19451) );
  INVX0 U20314 ( .IN(n19434), .QN(n19418) );
  INVX0 U20315 ( .IN(n19401), .QN(n19385) );
  INVX0 U20316 ( .IN(n19438), .QN(n19431) );
  INVX0 U20317 ( .IN(n19405), .QN(n19398) );
  INVX0 U20318 ( .IN(n19339), .QN(n19334) );
  INVX0 U20319 ( .IN(n19306), .QN(n19301) );
  INVX0 U20320 ( .IN(n19273), .QN(n19268) );
  INVX0 U20321 ( .IN(n19335), .QN(n19317) );
  INVX0 U20322 ( .IN(n19302), .QN(n19284) );
  INVX0 U20323 ( .IN(n19269), .QN(n19251) );
  INVX0 U20324 ( .IN(n19335), .QN(n19318) );
  INVX0 U20325 ( .IN(n19302), .QN(n19285) );
  INVX0 U20326 ( .IN(n19269), .QN(n19252) );
  INVX0 U20327 ( .IN(n19335), .QN(n19319) );
  INVX0 U20328 ( .IN(n19302), .QN(n19286) );
  INVX0 U20329 ( .IN(n19269), .QN(n19253) );
  INVX0 U20330 ( .IN(n19306), .QN(n19299) );
  INVX0 U20331 ( .IN(n19273), .QN(n19266) );
  INVX0 U20332 ( .IN(n19207), .QN(n19202) );
  INVX0 U20333 ( .IN(n19174), .QN(n19169) );
  INVX0 U20334 ( .IN(n19141), .QN(n19136) );
  INVX0 U20335 ( .IN(n19203), .QN(n19185) );
  INVX0 U20336 ( .IN(n19170), .QN(n19152) );
  INVX0 U20337 ( .IN(n19137), .QN(n19119) );
  INVX0 U20338 ( .IN(n19203), .QN(n19186) );
  INVX0 U20339 ( .IN(n19170), .QN(n19153) );
  INVX0 U20340 ( .IN(n19137), .QN(n19120) );
  INVX0 U20341 ( .IN(n19203), .QN(n19187) );
  INVX0 U20342 ( .IN(n19170), .QN(n19154) );
  INVX0 U20343 ( .IN(n19137), .QN(n19121) );
  INVX0 U20344 ( .IN(n19174), .QN(n19168) );
  INVX0 U20345 ( .IN(n19141), .QN(n19134) );
  INVX0 U20346 ( .IN(n19075), .QN(n19070) );
  INVX0 U20347 ( .IN(n19071), .QN(n19053) );
  INVX0 U20348 ( .IN(n19005), .QN(n18987) );
  INVX0 U20349 ( .IN(n19071), .QN(n19054) );
  INVX0 U20350 ( .IN(n19042), .QN(n19020) );
  INVX0 U20351 ( .IN(n19005), .QN(n18988) );
  INVX0 U20352 ( .IN(n19071), .QN(n19055) );
  INVX0 U20353 ( .IN(n19005), .QN(n18989) );
  INVX0 U20354 ( .IN(n19041), .QN(n19036) );
  INVX0 U20355 ( .IN(n20789), .QN(n20784) );
  INVX0 U20356 ( .IN(n20756), .QN(n20751) );
  INVX0 U20357 ( .IN(n20785), .QN(n20767) );
  INVX0 U20358 ( .IN(n20752), .QN(n20734) );
  INVX0 U20359 ( .IN(n20719), .QN(n20701) );
  INVX0 U20360 ( .IN(n20785), .QN(n20768) );
  INVX0 U20361 ( .IN(n20752), .QN(n20735) );
  INVX0 U20362 ( .IN(n20719), .QN(n20702) );
  INVX0 U20363 ( .IN(n20785), .QN(n20769) );
  INVX0 U20364 ( .IN(n20752), .QN(n20736) );
  INVX0 U20365 ( .IN(n20719), .QN(n20703) );
  INVX0 U20366 ( .IN(n20756), .QN(n20750) );
  INVX0 U20367 ( .IN(n20657), .QN(n20652) );
  INVX0 U20368 ( .IN(n20621), .QN(n20620) );
  INVX0 U20369 ( .IN(n20591), .QN(n20586) );
  INVX0 U20370 ( .IN(n20653), .QN(n20635) );
  INVX0 U20371 ( .IN(n20621), .QN(n20602) );
  INVX0 U20372 ( .IN(n20587), .QN(n20569) );
  INVX0 U20373 ( .IN(n20653), .QN(n20636) );
  INVX0 U20374 ( .IN(n20621), .QN(n20603) );
  INVX0 U20375 ( .IN(n20587), .QN(n20570) );
  INVX0 U20376 ( .IN(n20653), .QN(n20637) );
  INVX0 U20377 ( .IN(n20621), .QN(n20604) );
  INVX0 U20378 ( .IN(n20587), .QN(n20571) );
  INVX0 U20379 ( .IN(n20657), .QN(n20650) );
  INVX0 U20380 ( .IN(n20624), .QN(n20618) );
  INVX0 U20381 ( .IN(n20591), .QN(n20584) );
  INVX0 U20382 ( .IN(n20525), .QN(n20520) );
  INVX0 U20383 ( .IN(n20489), .QN(n20488) );
  INVX0 U20384 ( .IN(n20459), .QN(n20454) );
  INVX0 U20385 ( .IN(n20521), .QN(n20503) );
  INVX0 U20386 ( .IN(n20489), .QN(n20470) );
  INVX0 U20387 ( .IN(n20455), .QN(n20437) );
  INVX0 U20388 ( .IN(n20521), .QN(n20504) );
  INVX0 U20389 ( .IN(n20489), .QN(n20471) );
  INVX0 U20390 ( .IN(n20455), .QN(n20438) );
  INVX0 U20391 ( .IN(n20521), .QN(n20505) );
  INVX0 U20392 ( .IN(n20489), .QN(n20472) );
  INVX0 U20393 ( .IN(n20455), .QN(n20439) );
  INVX0 U20394 ( .IN(n20525), .QN(n20518) );
  INVX0 U20395 ( .IN(n20492), .QN(n20487) );
  INVX0 U20396 ( .IN(n20459), .QN(n20452) );
  INVX0 U20397 ( .IN(n20393), .QN(n20388) );
  INVX0 U20398 ( .IN(n20360), .QN(n20355) );
  INVX0 U20399 ( .IN(n20327), .QN(n20322) );
  INVX0 U20400 ( .IN(n20389), .QN(n20371) );
  INVX0 U20401 ( .IN(n20356), .QN(n20338) );
  INVX0 U20402 ( .IN(n20323), .QN(n20305) );
  INVX0 U20403 ( .IN(n20389), .QN(n20372) );
  INVX0 U20404 ( .IN(n20356), .QN(n20339) );
  INVX0 U20405 ( .IN(n20323), .QN(n20306) );
  INVX0 U20406 ( .IN(n20389), .QN(n20373) );
  INVX0 U20407 ( .IN(n20356), .QN(n20340) );
  INVX0 U20408 ( .IN(n20323), .QN(n20307) );
  INVX0 U20409 ( .IN(n20393), .QN(n20386) );
  INVX0 U20410 ( .IN(n20360), .QN(n20353) );
  INVX0 U20411 ( .IN(n20327), .QN(n20320) );
  INVX0 U20412 ( .IN(n20261), .QN(n20256) );
  INVX0 U20413 ( .IN(n20228), .QN(n20223) );
  INVX0 U20414 ( .IN(n20195), .QN(n20190) );
  INVX0 U20415 ( .IN(n20257), .QN(n20239) );
  INVX0 U20416 ( .IN(n20224), .QN(n20206) );
  INVX0 U20417 ( .IN(n20191), .QN(n20173) );
  INVX0 U20418 ( .IN(n20257), .QN(n20240) );
  INVX0 U20419 ( .IN(n20224), .QN(n20207) );
  INVX0 U20420 ( .IN(n20191), .QN(n20174) );
  INVX0 U20421 ( .IN(n20257), .QN(n20241) );
  INVX0 U20422 ( .IN(n20224), .QN(n20208) );
  INVX0 U20423 ( .IN(n20191), .QN(n20175) );
  INVX0 U20424 ( .IN(n20261), .QN(n20254) );
  INVX0 U20425 ( .IN(n20228), .QN(n20221) );
  INVX0 U20426 ( .IN(n20195), .QN(n20188) );
  INVX0 U20427 ( .IN(n20129), .QN(n20124) );
  INVX0 U20428 ( .IN(n20125), .QN(n20107) );
  INVX0 U20429 ( .IN(n20093), .QN(n20075) );
  INVX0 U20430 ( .IN(n20060), .QN(n20042) );
  INVX0 U20431 ( .IN(n20125), .QN(n20108) );
  INVX0 U20432 ( .IN(n20093), .QN(n20076) );
  INVX0 U20433 ( .IN(n20060), .QN(n20043) );
  INVX0 U20434 ( .IN(n20125), .QN(n20109) );
  INVX0 U20435 ( .IN(n20093), .QN(n20077) );
  INVX0 U20436 ( .IN(n20060), .QN(n20044) );
  INVX0 U20437 ( .IN(n20095), .QN(n20091) );
  INVX0 U20438 ( .IN(n19998), .QN(n19993) );
  INVX0 U20439 ( .IN(n19962), .QN(n19961) );
  INVX0 U20440 ( .IN(n19994), .QN(n19976) );
  INVX0 U20441 ( .IN(n19962), .QN(n19944) );
  INVX0 U20442 ( .IN(n19929), .QN(n19911) );
  INVX0 U20443 ( .IN(n19994), .QN(n19977) );
  INVX0 U20444 ( .IN(n19962), .QN(n19945) );
  INVX0 U20445 ( .IN(n19929), .QN(n19912) );
  INVX0 U20446 ( .IN(n19994), .QN(n19978) );
  INVX0 U20447 ( .IN(n19962), .QN(n19946) );
  INVX0 U20448 ( .IN(n19929), .QN(n19913) );
  INVX0 U20449 ( .IN(n19962), .QN(n19959) );
  INVX0 U20450 ( .IN(n19867), .QN(n19862) );
  INVX0 U20451 ( .IN(n19863), .QN(n19845) );
  INVX0 U20452 ( .IN(n19797), .QN(n19779) );
  INVX0 U20453 ( .IN(n19863), .QN(n19846) );
  INVX0 U20454 ( .IN(n19834), .QN(n19812) );
  INVX0 U20455 ( .IN(n19797), .QN(n19780) );
  INVX0 U20456 ( .IN(n19863), .QN(n19847) );
  INVX0 U20457 ( .IN(n19797), .QN(n19781) );
  INVX0 U20458 ( .IN(n19833), .QN(n19828) );
  INVX0 U20459 ( .IN(n18943), .QN(n18938) );
  INVX0 U20460 ( .IN(n18939), .QN(n18921) );
  INVX0 U20461 ( .IN(n18873), .QN(n18855) );
  INVX0 U20462 ( .IN(n18939), .QN(n18922) );
  INVX0 U20463 ( .IN(n18910), .QN(n18888) );
  INVX0 U20464 ( .IN(n18873), .QN(n18856) );
  INVX0 U20465 ( .IN(n18939), .QN(n18923) );
  INVX0 U20466 ( .IN(n18873), .QN(n18857) );
  INVX0 U20467 ( .IN(n18909), .QN(n18904) );
  INVX0 U20468 ( .IN(n21075), .QN(n21053) );
  INVX0 U20469 ( .IN(n21073), .QN(n21057) );
  INVX0 U20470 ( .IN(n21074), .QN(n21054) );
  INVX0 U20471 ( .IN(n21072), .QN(n21058) );
  INVX0 U20472 ( .IN(n21074), .QN(n21055) );
  INVX0 U20473 ( .IN(n21073), .QN(n21056) );
  INVX0 U20474 ( .IN(n21072), .QN(n21059) );
  INVX0 U20475 ( .IN(n21075), .QN(n21052) );
  INVX0 U20476 ( .IN(n17885), .QN(n19481) );
  INVX0 U20477 ( .IN(n17886), .QN(n19349) );
  INVX0 U20478 ( .IN(n17887), .QN(n19217) );
  INVX0 U20479 ( .IN(n17888), .QN(n19085) );
  INVX0 U20480 ( .IN(n17889), .QN(n18953) );
  INVX0 U20481 ( .IN(n17890), .QN(n20667) );
  INVX0 U20482 ( .IN(n17891), .QN(n20535) );
  INVX0 U20483 ( .IN(n17892), .QN(n20403) );
  INVX0 U20484 ( .IN(n17893), .QN(n20271) );
  INVX0 U20485 ( .IN(n17894), .QN(n20139) );
  INVX0 U20486 ( .IN(n17895), .QN(n20008) );
  INVX0 U20487 ( .IN(n17896), .QN(n19877) );
  INVX0 U20488 ( .IN(n17897), .QN(n19745) );
  INVX0 U20489 ( .IN(n17898), .QN(n18821) );
  INVX0 U20490 ( .IN(n21071), .QN(n21060) );
  INVX0 U20491 ( .IN(n21069), .QN(n21065) );
  INVX0 U20492 ( .IN(n21070), .QN(n21062) );
  INVX0 U20493 ( .IN(n21069), .QN(n21064) );
  INVX0 U20494 ( .IN(n21070), .QN(n21063) );
  INVX0 U20495 ( .IN(n21071), .QN(n21061) );
  INVX0 U20496 ( .IN(n19481), .QN(n19504) );
  INVX0 U20497 ( .IN(n20139), .QN(n20162) );
  INVX0 U20498 ( .IN(n19349), .QN(n19372) );
  INVX0 U20499 ( .IN(n19217), .QN(n19240) );
  INVX0 U20500 ( .IN(n20008), .QN(n20031) );
  INVX0 U20501 ( .IN(n19877), .QN(n19900) );
  INVX0 U20502 ( .IN(n19085), .QN(n19108) );
  INVX0 U20503 ( .IN(n18953), .QN(n18976) );
  INVX0 U20504 ( .IN(n19745), .QN(n19768) );
  INVX0 U20505 ( .IN(n18821), .QN(n18844) );
  INVX0 U20506 ( .IN(n20667), .QN(n20690) );
  INVX0 U20507 ( .IN(n18297), .QN(n18387) );
  INVX0 U20508 ( .IN(n18291), .QN(n18391) );
  INVX0 U20509 ( .IN(n18296), .QN(n18371) );
  INVX0 U20510 ( .IN(n21068), .QN(n21051) );
  INVX0 U20511 ( .IN(n21077), .QN(n21050) );
  INVX0 U20512 ( .IN(n21076), .QN(n21049) );
  INVX0 U20513 ( .IN(n21076), .QN(n21048) );
  INVX0 U20514 ( .IN(n21077), .QN(n21047) );
  INVX0 U20515 ( .IN(n21077), .QN(n21046) );
  INVX0 U20516 ( .IN(n21076), .QN(n21045) );
  INVX0 U20517 ( .IN(n17780), .QN(n18815) );
  INVX0 U20518 ( .IN(n18815), .QN(n18820) );
  INVX0 U20519 ( .IN(n19712), .QN(n19732) );
  INVX0 U20520 ( .IN(n19679), .QN(n19699) );
  INVX0 U20521 ( .IN(n19646), .QN(n19666) );
  INVX0 U20522 ( .IN(n19712), .QN(n19731) );
  INVX0 U20523 ( .IN(n19679), .QN(n19698) );
  INVX0 U20524 ( .IN(n19646), .QN(n19665) );
  INVX0 U20525 ( .IN(n19714), .QN(n19735) );
  INVX0 U20526 ( .IN(n19715), .QN(n19714) );
  INVX0 U20527 ( .IN(n19648), .QN(n19669) );
  INVX0 U20528 ( .IN(n19649), .QN(n19648) );
  INVX0 U20529 ( .IN(n7178), .QN(n19616) );
  INVX0 U20530 ( .IN(n19681), .QN(n19702) );
  INVX0 U20531 ( .IN(n19682), .QN(n19681) );
  INVX0 U20532 ( .IN(n19618), .QN(n19613) );
  INVX0 U20533 ( .IN(n7178), .QN(n19618) );
  INVX0 U20534 ( .IN(n19744), .QN(n19736) );
  INVX0 U20535 ( .IN(n19711), .QN(n19703) );
  INVX0 U20536 ( .IN(n19678), .QN(n19670) );
  INVX0 U20537 ( .IN(n19645), .QN(n19637) );
  INVX0 U20538 ( .IN(n19683), .QN(n19680) );
  INVX0 U20539 ( .IN(n19650), .QN(n19647) );
  INVX0 U20540 ( .IN(n19716), .QN(n19713) );
  INVX0 U20541 ( .IN(n7178), .QN(n19617) );
  NAND2X0 U20542 ( .IN1(n17781), .IN2(n19744), .QN(n14496) );
  NAND2X0 U20543 ( .IN1(n17782), .IN2(n19711), .QN(n15186) );
  NAND2X0 U20544 ( .IN1(n17783), .IN2(n19678), .QN(n15796) );
  NAND2X0 U20545 ( .IN1(n17784), .IN2(n19645), .QN(n16406) );
  AND2X1 U20546 ( .IN1(n9601), .IN2(n9912), .Q(n18286) );
  AND2X1 U20547 ( .IN1(n9601), .IN2(n9602), .Q(n18287) );
  AND2X1 U20548 ( .IN1(n11770), .IN2(n10841), .Q(n18288) );
  AND2X1 U20549 ( .IN1(n11770), .IN2(n9601), .Q(n18289) );
  AND2X1 U20550 ( .IN1(n11770), .IN2(n11460), .Q(n18290) );
  AND2X1 U20551 ( .IN1(n11770), .IN2(n10222), .Q(n18291) );
  AND2X1 U20552 ( .IN1(n10222), .IN2(n9912), .Q(n18292) );
  AND2X1 U20553 ( .IN1(n10222), .IN2(n9602), .Q(n18293) );
  AND2X1 U20554 ( .IN1(n12080), .IN2(n10841), .Q(n18294) );
  AND2X1 U20555 ( .IN1(n12080), .IN2(n9601), .Q(n18295) );
  AND2X1 U20556 ( .IN1(n12080), .IN2(n11460), .Q(n18296) );
  AND2X1 U20557 ( .IN1(n12080), .IN2(n10222), .Q(n18297) );
  AND2X1 U20558 ( .IN1(n11460), .IN2(n9912), .Q(n18298) );
  AND2X1 U20559 ( .IN1(n9602), .IN2(n11460), .Q(n18299) );
  AND2X1 U20560 ( .IN1(n10841), .IN2(n9912), .Q(n18300) );
  AND2X1 U20561 ( .IN1(n10841), .IN2(n9602), .Q(n18301) );
  INVX0 U20562 ( .IN(n17873), .QN(n18799) );
  INVX0 U20563 ( .IN(n17795), .QN(n18787) );
  INVX0 U20564 ( .IN(n17793), .QN(n18775) );
  INVX0 U20565 ( .IN(n17873), .QN(n18797) );
  INVX0 U20566 ( .IN(n17795), .QN(n18785) );
  INVX0 U20567 ( .IN(n17793), .QN(n18773) );
  INVX0 U20568 ( .IN(n17793), .QN(n18774) );
  INVX0 U20569 ( .IN(n17873), .QN(n18798) );
  INVX0 U20570 ( .IN(n17795), .QN(n18786) );
  INVX0 U20571 ( .IN(n17877), .QN(n18751) );
  INVX0 U20572 ( .IN(n17835), .QN(n18739) );
  INVX0 U20573 ( .IN(n18727), .QN(n18726) );
  INVX0 U20574 ( .IN(n17877), .QN(n18749) );
  INVX0 U20575 ( .IN(n17835), .QN(n18737) );
  INVX0 U20576 ( .IN(n17877), .QN(n18750) );
  INVX0 U20577 ( .IN(n17835), .QN(n18738) );
  INVX0 U20578 ( .IN(n18727), .QN(n18725) );
  INVX0 U20579 ( .IN(n17874), .QN(n18703) );
  INVX0 U20580 ( .IN(n17799), .QN(n18691) );
  INVX0 U20581 ( .IN(n17797), .QN(n18679) );
  INVX0 U20582 ( .IN(n17874), .QN(n18701) );
  INVX0 U20583 ( .IN(n17799), .QN(n18689) );
  INVX0 U20584 ( .IN(n17797), .QN(n18677) );
  INVX0 U20585 ( .IN(n17874), .QN(n18702) );
  INVX0 U20586 ( .IN(n17797), .QN(n18678) );
  INVX0 U20587 ( .IN(n17799), .QN(n18690) );
  INVX0 U20588 ( .IN(n17878), .QN(n18655) );
  INVX0 U20589 ( .IN(n17838), .QN(n18643) );
  INVX0 U20590 ( .IN(n18631), .QN(n18630) );
  INVX0 U20591 ( .IN(n17878), .QN(n18653) );
  INVX0 U20592 ( .IN(n17838), .QN(n18641) );
  INVX0 U20593 ( .IN(n17838), .QN(n18642) );
  INVX0 U20594 ( .IN(n18631), .QN(n18629) );
  INVX0 U20595 ( .IN(n17878), .QN(n18654) );
  INVX0 U20596 ( .IN(n17875), .QN(n18607) );
  INVX0 U20597 ( .IN(n17803), .QN(n18595) );
  INVX0 U20598 ( .IN(n17801), .QN(n18583) );
  INVX0 U20599 ( .IN(n17875), .QN(n18605) );
  INVX0 U20600 ( .IN(n17803), .QN(n18593) );
  INVX0 U20601 ( .IN(n17801), .QN(n18581) );
  INVX0 U20602 ( .IN(n17875), .QN(n18606) );
  INVX0 U20603 ( .IN(n17801), .QN(n18582) );
  INVX0 U20604 ( .IN(n17803), .QN(n18594) );
  INVX0 U20605 ( .IN(n17879), .QN(n18559) );
  INVX0 U20606 ( .IN(n17841), .QN(n18547) );
  INVX0 U20607 ( .IN(n18535), .QN(n18534) );
  INVX0 U20608 ( .IN(n17879), .QN(n18557) );
  INVX0 U20609 ( .IN(n17841), .QN(n18545) );
  INVX0 U20610 ( .IN(n17841), .QN(n18546) );
  INVX0 U20611 ( .IN(n18535), .QN(n18533) );
  INVX0 U20612 ( .IN(n17879), .QN(n18558) );
  INVX0 U20613 ( .IN(n17876), .QN(n18511) );
  INVX0 U20614 ( .IN(n17807), .QN(n18499) );
  INVX0 U20615 ( .IN(n17805), .QN(n18487) );
  INVX0 U20616 ( .IN(n17876), .QN(n18509) );
  INVX0 U20617 ( .IN(n17807), .QN(n18497) );
  INVX0 U20618 ( .IN(n17805), .QN(n18485) );
  INVX0 U20619 ( .IN(n17876), .QN(n18510) );
  INVX0 U20620 ( .IN(n17805), .QN(n18486) );
  INVX0 U20621 ( .IN(n17807), .QN(n18498) );
  INVX0 U20622 ( .IN(n17880), .QN(n18463) );
  INVX0 U20623 ( .IN(n17844), .QN(n18451) );
  INVX0 U20624 ( .IN(n18439), .QN(n18438) );
  INVX0 U20625 ( .IN(n17880), .QN(n18461) );
  INVX0 U20626 ( .IN(n17844), .QN(n18449) );
  INVX0 U20627 ( .IN(n17844), .QN(n18450) );
  INVX0 U20628 ( .IN(n18439), .QN(n18437) );
  INVX0 U20629 ( .IN(n17880), .QN(n18462) );
  INVX0 U20630 ( .IN(n17817), .QN(n18814) );
  INVX0 U20631 ( .IN(n17830), .QN(n18802) );
  INVX0 U20632 ( .IN(n17796), .QN(n18790) );
  INVX0 U20633 ( .IN(n17794), .QN(n18778) );
  INVX0 U20634 ( .IN(n17817), .QN(n18812) );
  INVX0 U20635 ( .IN(n17830), .QN(n18800) );
  INVX0 U20636 ( .IN(n17817), .QN(n18813) );
  INVX0 U20637 ( .IN(n17830), .QN(n18801) );
  INVX0 U20638 ( .IN(n17796), .QN(n18788) );
  INVX0 U20639 ( .IN(n17794), .QN(n18776) );
  INVX0 U20640 ( .IN(n17796), .QN(n18789) );
  INVX0 U20641 ( .IN(n17794), .QN(n18777) );
  INVX0 U20642 ( .IN(n17854), .QN(n18766) );
  INVX0 U20643 ( .IN(n17865), .QN(n18754) );
  INVX0 U20644 ( .IN(n17836), .QN(n18742) );
  INVX0 U20645 ( .IN(n17834), .QN(n18730) );
  INVX0 U20646 ( .IN(n17854), .QN(n18764) );
  INVX0 U20647 ( .IN(n17854), .QN(n18765) );
  INVX0 U20648 ( .IN(n17865), .QN(n18752) );
  INVX0 U20649 ( .IN(n17836), .QN(n18740) );
  INVX0 U20650 ( .IN(n17834), .QN(n18728) );
  INVX0 U20651 ( .IN(n17865), .QN(n18753) );
  INVX0 U20652 ( .IN(n17836), .QN(n18741) );
  INVX0 U20653 ( .IN(n17834), .QN(n18729) );
  INVX0 U20654 ( .IN(n17827), .QN(n18718) );
  INVX0 U20655 ( .IN(n17831), .QN(n18706) );
  INVX0 U20656 ( .IN(n17800), .QN(n18694) );
  INVX0 U20657 ( .IN(n17798), .QN(n18682) );
  INVX0 U20658 ( .IN(n17827), .QN(n18716) );
  INVX0 U20659 ( .IN(n17827), .QN(n18717) );
  INVX0 U20660 ( .IN(n17831), .QN(n18704) );
  INVX0 U20661 ( .IN(n17800), .QN(n18692) );
  INVX0 U20662 ( .IN(n17798), .QN(n18680) );
  INVX0 U20663 ( .IN(n17800), .QN(n18693) );
  INVX0 U20664 ( .IN(n17798), .QN(n18681) );
  INVX0 U20665 ( .IN(n17831), .QN(n18705) );
  INVX0 U20666 ( .IN(n17855), .QN(n18670) );
  INVX0 U20667 ( .IN(n17866), .QN(n18658) );
  INVX0 U20668 ( .IN(n17839), .QN(n18646) );
  INVX0 U20669 ( .IN(n17837), .QN(n18634) );
  INVX0 U20670 ( .IN(n17855), .QN(n18668) );
  INVX0 U20671 ( .IN(n17855), .QN(n18669) );
  INVX0 U20672 ( .IN(n17866), .QN(n18656) );
  INVX0 U20673 ( .IN(n17839), .QN(n18644) );
  INVX0 U20674 ( .IN(n17837), .QN(n18632) );
  INVX0 U20675 ( .IN(n17839), .QN(n18645) );
  INVX0 U20676 ( .IN(n17837), .QN(n18633) );
  INVX0 U20677 ( .IN(n17866), .QN(n18657) );
  INVX0 U20678 ( .IN(n17818), .QN(n18622) );
  INVX0 U20679 ( .IN(n17804), .QN(n18598) );
  INVX0 U20680 ( .IN(n17802), .QN(n18586) );
  INVX0 U20681 ( .IN(n17818), .QN(n18620) );
  INVX0 U20682 ( .IN(n17832), .QN(n18608) );
  INVX0 U20683 ( .IN(n17818), .QN(n18621) );
  INVX0 U20684 ( .IN(n17832), .QN(n18609) );
  INVX0 U20685 ( .IN(n17804), .QN(n18596) );
  INVX0 U20686 ( .IN(n17802), .QN(n18584) );
  INVX0 U20687 ( .IN(n17832), .QN(n18610) );
  INVX0 U20688 ( .IN(n17804), .QN(n18597) );
  INVX0 U20689 ( .IN(n17802), .QN(n18585) );
  INVX0 U20690 ( .IN(n17856), .QN(n18574) );
  INVX0 U20691 ( .IN(n17867), .QN(n18562) );
  INVX0 U20692 ( .IN(n17842), .QN(n18550) );
  INVX0 U20693 ( .IN(n17840), .QN(n18538) );
  INVX0 U20694 ( .IN(n17856), .QN(n18572) );
  INVX0 U20695 ( .IN(n17856), .QN(n18573) );
  INVX0 U20696 ( .IN(n17867), .QN(n18560) );
  INVX0 U20697 ( .IN(n17842), .QN(n18548) );
  INVX0 U20698 ( .IN(n17840), .QN(n18536) );
  INVX0 U20699 ( .IN(n17842), .QN(n18549) );
  INVX0 U20700 ( .IN(n17840), .QN(n18537) );
  INVX0 U20701 ( .IN(n17867), .QN(n18561) );
  INVX0 U20702 ( .IN(n17819), .QN(n18526) );
  INVX0 U20703 ( .IN(n17833), .QN(n18514) );
  INVX0 U20704 ( .IN(n17808), .QN(n18502) );
  INVX0 U20705 ( .IN(n17806), .QN(n18490) );
  INVX0 U20706 ( .IN(n17819), .QN(n18524) );
  INVX0 U20707 ( .IN(n17819), .QN(n18525) );
  INVX0 U20708 ( .IN(n17833), .QN(n18512) );
  INVX0 U20709 ( .IN(n17808), .QN(n18500) );
  INVX0 U20710 ( .IN(n17806), .QN(n18488) );
  INVX0 U20711 ( .IN(n17808), .QN(n18501) );
  INVX0 U20712 ( .IN(n17806), .QN(n18489) );
  INVX0 U20713 ( .IN(n17833), .QN(n18513) );
  INVX0 U20714 ( .IN(n17857), .QN(n18478) );
  INVX0 U20715 ( .IN(n17868), .QN(n18466) );
  INVX0 U20716 ( .IN(n17845), .QN(n18454) );
  INVX0 U20717 ( .IN(n17843), .QN(n18442) );
  INVX0 U20718 ( .IN(n17857), .QN(n18476) );
  INVX0 U20719 ( .IN(n17857), .QN(n18477) );
  INVX0 U20720 ( .IN(n17868), .QN(n18464) );
  INVX0 U20721 ( .IN(n17845), .QN(n18452) );
  INVX0 U20722 ( .IN(n17843), .QN(n18440) );
  INVX0 U20723 ( .IN(n17845), .QN(n18453) );
  INVX0 U20724 ( .IN(n17843), .QN(n18441) );
  INVX0 U20725 ( .IN(n17868), .QN(n18465) );
  INVX0 U20726 ( .IN(n17810), .QN(n18808) );
  INVX0 U20727 ( .IN(n17820), .QN(n18796) );
  INVX0 U20728 ( .IN(n17882), .QN(n18784) );
  INVX0 U20729 ( .IN(n17824), .QN(n18772) );
  INVX0 U20730 ( .IN(n17810), .QN(n18806) );
  INVX0 U20731 ( .IN(n17882), .QN(n18782) );
  INVX0 U20732 ( .IN(n17824), .QN(n18770) );
  INVX0 U20733 ( .IN(n17810), .QN(n18807) );
  INVX0 U20734 ( .IN(n17824), .QN(n18771) );
  INVX0 U20735 ( .IN(n17820), .QN(n18794) );
  INVX0 U20736 ( .IN(n17820), .QN(n18795) );
  INVX0 U20737 ( .IN(n17882), .QN(n18783) );
  INVX0 U20738 ( .IN(n17858), .QN(n18736) );
  INVX0 U20739 ( .IN(n17859), .QN(n18724) );
  INVX0 U20740 ( .IN(n17846), .QN(n18758) );
  INVX0 U20741 ( .IN(n17850), .QN(n18746) );
  INVX0 U20742 ( .IN(n17846), .QN(n18759) );
  INVX0 U20743 ( .IN(n17850), .QN(n18747) );
  INVX0 U20744 ( .IN(n17858), .QN(n18734) );
  INVX0 U20745 ( .IN(n17859), .QN(n18722) );
  INVX0 U20746 ( .IN(n17850), .QN(n18748) );
  INVX0 U20747 ( .IN(n17846), .QN(n18760) );
  INVX0 U20748 ( .IN(n17858), .QN(n18735) );
  INVX0 U20749 ( .IN(n17859), .QN(n18723) );
  INVX0 U20750 ( .IN(n17812), .QN(n18712) );
  INVX0 U20751 ( .IN(n17821), .QN(n18700) );
  INVX0 U20752 ( .IN(n17828), .QN(n18688) );
  INVX0 U20753 ( .IN(n17829), .QN(n18676) );
  INVX0 U20754 ( .IN(n17812), .QN(n18710) );
  INVX0 U20755 ( .IN(n17821), .QN(n18698) );
  INVX0 U20756 ( .IN(n17829), .QN(n18674) );
  INVX0 U20757 ( .IN(n17812), .QN(n18711) );
  INVX0 U20758 ( .IN(n17829), .QN(n18675) );
  INVX0 U20759 ( .IN(n17821), .QN(n18699) );
  INVX0 U20760 ( .IN(n17828), .QN(n18686) );
  INVX0 U20761 ( .IN(n17828), .QN(n18687) );
  INVX0 U20762 ( .IN(n17789), .QN(n18640) );
  INVX0 U20763 ( .IN(n17860), .QN(n18628) );
  INVX0 U20764 ( .IN(n17847), .QN(n18662) );
  INVX0 U20765 ( .IN(n17851), .QN(n18650) );
  INVX0 U20766 ( .IN(n17847), .QN(n18663) );
  INVX0 U20767 ( .IN(n17851), .QN(n18651) );
  INVX0 U20768 ( .IN(n17789), .QN(n18638) );
  INVX0 U20769 ( .IN(n17860), .QN(n18626) );
  INVX0 U20770 ( .IN(n17851), .QN(n18652) );
  INVX0 U20771 ( .IN(n17847), .QN(n18664) );
  INVX0 U20772 ( .IN(n17789), .QN(n18639) );
  INVX0 U20773 ( .IN(n17860), .QN(n18627) );
  INVX0 U20774 ( .IN(n17814), .QN(n18616) );
  INVX0 U20775 ( .IN(n17822), .QN(n18604) );
  INVX0 U20776 ( .IN(n17883), .QN(n18592) );
  INVX0 U20777 ( .IN(n17825), .QN(n18580) );
  INVX0 U20778 ( .IN(n17814), .QN(n18614) );
  INVX0 U20779 ( .IN(n17822), .QN(n18602) );
  INVX0 U20780 ( .IN(n17883), .QN(n18590) );
  INVX0 U20781 ( .IN(n17825), .QN(n18578) );
  INVX0 U20782 ( .IN(n17814), .QN(n18615) );
  INVX0 U20783 ( .IN(n17825), .QN(n18579) );
  INVX0 U20784 ( .IN(n17822), .QN(n18603) );
  INVX0 U20785 ( .IN(n17883), .QN(n18591) );
  INVX0 U20786 ( .IN(n17861), .QN(n18544) );
  INVX0 U20787 ( .IN(n17862), .QN(n18532) );
  INVX0 U20788 ( .IN(n17848), .QN(n18566) );
  INVX0 U20789 ( .IN(n17852), .QN(n18554) );
  INVX0 U20790 ( .IN(n17848), .QN(n18567) );
  INVX0 U20791 ( .IN(n17852), .QN(n18555) );
  INVX0 U20792 ( .IN(n17861), .QN(n18542) );
  INVX0 U20793 ( .IN(n17862), .QN(n18530) );
  INVX0 U20794 ( .IN(n17852), .QN(n18556) );
  INVX0 U20795 ( .IN(n17848), .QN(n18568) );
  INVX0 U20796 ( .IN(n17861), .QN(n18543) );
  INVX0 U20797 ( .IN(n17862), .QN(n18531) );
  INVX0 U20798 ( .IN(n17816), .QN(n18520) );
  INVX0 U20799 ( .IN(n17823), .QN(n18508) );
  INVX0 U20800 ( .IN(n17884), .QN(n18496) );
  INVX0 U20801 ( .IN(n17826), .QN(n18484) );
  INVX0 U20802 ( .IN(n17816), .QN(n18518) );
  INVX0 U20803 ( .IN(n17823), .QN(n18506) );
  INVX0 U20804 ( .IN(n17884), .QN(n18494) );
  INVX0 U20805 ( .IN(n17826), .QN(n18482) );
  INVX0 U20806 ( .IN(n17816), .QN(n18519) );
  INVX0 U20807 ( .IN(n17826), .QN(n18483) );
  INVX0 U20808 ( .IN(n17823), .QN(n18507) );
  INVX0 U20809 ( .IN(n17884), .QN(n18495) );
  INVX0 U20810 ( .IN(n17863), .QN(n18448) );
  INVX0 U20811 ( .IN(n17864), .QN(n18436) );
  INVX0 U20812 ( .IN(n17849), .QN(n18470) );
  INVX0 U20813 ( .IN(n17853), .QN(n18458) );
  INVX0 U20814 ( .IN(n17849), .QN(n18471) );
  INVX0 U20815 ( .IN(n17853), .QN(n18459) );
  INVX0 U20816 ( .IN(n17863), .QN(n18446) );
  INVX0 U20817 ( .IN(n17864), .QN(n18434) );
  INVX0 U20818 ( .IN(n17853), .QN(n18460) );
  INVX0 U20819 ( .IN(n17849), .QN(n18472) );
  INVX0 U20820 ( .IN(n17863), .QN(n18447) );
  INVX0 U20821 ( .IN(n17864), .QN(n18435) );
  INVX0 U20822 ( .IN(n20870), .QN(n20869) );
  INVX0 U20823 ( .IN(n20852), .QN(n20851) );
  INVX0 U20824 ( .IN(n20834), .QN(n20833) );
  INVX0 U20825 ( .IN(n20816), .QN(n20815) );
  INVX0 U20826 ( .IN(n20870), .QN(n20865) );
  INVX0 U20827 ( .IN(n20852), .QN(n20849) );
  INVX0 U20828 ( .IN(n20834), .QN(n20831) );
  INVX0 U20829 ( .IN(n20816), .QN(n20813) );
  INVX0 U20830 ( .IN(n20870), .QN(n20862) );
  INVX0 U20831 ( .IN(n20852), .QN(n20844) );
  INVX0 U20832 ( .IN(n20834), .QN(n20826) );
  INVX0 U20833 ( .IN(n20816), .QN(n20808) );
  INVX0 U20834 ( .IN(n20870), .QN(n20863) );
  INVX0 U20835 ( .IN(n20852), .QN(n20845) );
  INVX0 U20836 ( .IN(n20834), .QN(n20827) );
  INVX0 U20837 ( .IN(n20816), .QN(n20809) );
  INVX0 U20838 ( .IN(n20870), .QN(n20864) );
  INVX0 U20839 ( .IN(n20852), .QN(n20846) );
  INVX0 U20840 ( .IN(n20834), .QN(n20828) );
  INVX0 U20841 ( .IN(n20816), .QN(n20810) );
  INVX0 U20842 ( .IN(n20852), .QN(n20847) );
  INVX0 U20843 ( .IN(n20834), .QN(n20829) );
  INVX0 U20844 ( .IN(n20816), .QN(n20811) );
  INVX0 U20845 ( .IN(n20852), .QN(n20848) );
  INVX0 U20846 ( .IN(n20834), .QN(n20830) );
  INVX0 U20847 ( .IN(n20816), .QN(n20812) );
  INVX0 U20848 ( .IN(n20852), .QN(n20850) );
  INVX0 U20849 ( .IN(n20834), .QN(n20832) );
  INVX0 U20850 ( .IN(n20816), .QN(n20814) );
  INVX0 U20851 ( .IN(n20870), .QN(n20866) );
  INVX0 U20852 ( .IN(n20870), .QN(n20867) );
  INVX0 U20853 ( .IN(n20870), .QN(n20868) );
  INVX0 U20854 ( .IN(n17809), .QN(n18805) );
  INVX0 U20855 ( .IN(n18793), .QN(n18792) );
  INVX0 U20856 ( .IN(n17869), .QN(n18781) );
  INVX0 U20857 ( .IN(n18769), .QN(n18768) );
  INVX0 U20858 ( .IN(n17809), .QN(n18803) );
  INVX0 U20859 ( .IN(n18793), .QN(n18791) );
  INVX0 U20860 ( .IN(n17869), .QN(n18779) );
  INVX0 U20861 ( .IN(n18769), .QN(n18767) );
  INVX0 U20862 ( .IN(n17809), .QN(n18804) );
  INVX0 U20863 ( .IN(n17869), .QN(n18780) );
  INVX0 U20864 ( .IN(n18757), .QN(n18756) );
  INVX0 U20865 ( .IN(n18745), .QN(n18744) );
  INVX0 U20866 ( .IN(n18733), .QN(n18732) );
  INVX0 U20867 ( .IN(n18721), .QN(n18720) );
  INVX0 U20868 ( .IN(n18757), .QN(n18755) );
  INVX0 U20869 ( .IN(n18745), .QN(n18743) );
  INVX0 U20870 ( .IN(n18721), .QN(n18719) );
  INVX0 U20871 ( .IN(n18733), .QN(n18731) );
  INVX0 U20872 ( .IN(n17811), .QN(n18709) );
  INVX0 U20873 ( .IN(n18697), .QN(n18696) );
  INVX0 U20874 ( .IN(n17872), .QN(n18685) );
  INVX0 U20875 ( .IN(n18673), .QN(n18672) );
  INVX0 U20876 ( .IN(n17811), .QN(n18707) );
  INVX0 U20877 ( .IN(n18697), .QN(n18695) );
  INVX0 U20878 ( .IN(n17872), .QN(n18683) );
  INVX0 U20879 ( .IN(n18673), .QN(n18671) );
  INVX0 U20880 ( .IN(n17811), .QN(n18708) );
  INVX0 U20881 ( .IN(n17872), .QN(n18684) );
  INVX0 U20882 ( .IN(n18661), .QN(n18660) );
  INVX0 U20883 ( .IN(n18649), .QN(n18648) );
  INVX0 U20884 ( .IN(n18637), .QN(n18636) );
  INVX0 U20885 ( .IN(n18625), .QN(n18624) );
  INVX0 U20886 ( .IN(n18661), .QN(n18659) );
  INVX0 U20887 ( .IN(n18649), .QN(n18647) );
  INVX0 U20888 ( .IN(n18625), .QN(n18623) );
  INVX0 U20889 ( .IN(n18637), .QN(n18635) );
  INVX0 U20890 ( .IN(n17813), .QN(n18613) );
  INVX0 U20891 ( .IN(n18601), .QN(n18600) );
  INVX0 U20892 ( .IN(n17870), .QN(n18589) );
  INVX0 U20893 ( .IN(n18577), .QN(n18576) );
  INVX0 U20894 ( .IN(n17813), .QN(n18611) );
  INVX0 U20895 ( .IN(n18601), .QN(n18599) );
  INVX0 U20896 ( .IN(n17870), .QN(n18587) );
  INVX0 U20897 ( .IN(n18577), .QN(n18575) );
  INVX0 U20898 ( .IN(n17813), .QN(n18612) );
  INVX0 U20899 ( .IN(n17870), .QN(n18588) );
  INVX0 U20900 ( .IN(n18565), .QN(n18564) );
  INVX0 U20901 ( .IN(n18553), .QN(n18552) );
  INVX0 U20902 ( .IN(n18541), .QN(n18540) );
  INVX0 U20903 ( .IN(n18529), .QN(n18528) );
  INVX0 U20904 ( .IN(n18565), .QN(n18563) );
  INVX0 U20905 ( .IN(n18553), .QN(n18551) );
  INVX0 U20906 ( .IN(n18529), .QN(n18527) );
  INVX0 U20907 ( .IN(n18541), .QN(n18539) );
  INVX0 U20908 ( .IN(n17815), .QN(n18517) );
  INVX0 U20909 ( .IN(n18505), .QN(n18504) );
  INVX0 U20910 ( .IN(n17871), .QN(n18493) );
  INVX0 U20911 ( .IN(n18481), .QN(n18480) );
  INVX0 U20912 ( .IN(n17815), .QN(n18515) );
  INVX0 U20913 ( .IN(n18505), .QN(n18503) );
  INVX0 U20914 ( .IN(n17871), .QN(n18491) );
  INVX0 U20915 ( .IN(n18481), .QN(n18479) );
  INVX0 U20916 ( .IN(n17815), .QN(n18516) );
  INVX0 U20917 ( .IN(n17871), .QN(n18492) );
  INVX0 U20918 ( .IN(n18469), .QN(n18468) );
  INVX0 U20919 ( .IN(n18457), .QN(n18456) );
  INVX0 U20920 ( .IN(n18445), .QN(n18444) );
  INVX0 U20921 ( .IN(n18433), .QN(n18432) );
  INVX0 U20922 ( .IN(n18469), .QN(n18467) );
  INVX0 U20923 ( .IN(n18457), .QN(n18455) );
  INVX0 U20924 ( .IN(n18433), .QN(n18431) );
  INVX0 U20925 ( .IN(n18445), .QN(n18443) );
  INVX0 U20926 ( .IN(n20861), .QN(n20860) );
  INVX0 U20927 ( .IN(n20861), .QN(n20858) );
  INVX0 U20928 ( .IN(n20843), .QN(n20839) );
  INVX0 U20929 ( .IN(n20825), .QN(n20821) );
  INVX0 U20930 ( .IN(n20861), .QN(n20853) );
  INVX0 U20931 ( .IN(n20843), .QN(n20835) );
  INVX0 U20932 ( .IN(n20825), .QN(n20817) );
  INVX0 U20933 ( .IN(n20861), .QN(n20854) );
  INVX0 U20934 ( .IN(n20843), .QN(n20836) );
  INVX0 U20935 ( .IN(n20825), .QN(n20818) );
  INVX0 U20936 ( .IN(n20861), .QN(n20855) );
  INVX0 U20937 ( .IN(n20843), .QN(n20837) );
  INVX0 U20938 ( .IN(n20825), .QN(n20819) );
  INVX0 U20939 ( .IN(n20861), .QN(n20856) );
  INVX0 U20940 ( .IN(n20843), .QN(n20838) );
  INVX0 U20941 ( .IN(n20825), .QN(n20820) );
  INVX0 U20942 ( .IN(n20861), .QN(n20857) );
  INVX0 U20943 ( .IN(n20843), .QN(n20842) );
  INVX0 U20944 ( .IN(n20825), .QN(n20824) );
  INVX0 U20945 ( .IN(n20843), .QN(n20840) );
  INVX0 U20946 ( .IN(n20825), .QN(n20822) );
  INVX0 U20947 ( .IN(n20861), .QN(n20859) );
  INVX0 U20948 ( .IN(n20843), .QN(n20841) );
  INVX0 U20949 ( .IN(n20825), .QN(n20823) );
  INVX0 U20950 ( .IN(n19744), .QN(n19738) );
  INVX0 U20951 ( .IN(n19711), .QN(n19705) );
  INVX0 U20952 ( .IN(n19678), .QN(n19672) );
  INVX0 U20953 ( .IN(n19645), .QN(n19639) );
  INVX0 U20954 ( .IN(n19744), .QN(n19739) );
  INVX0 U20955 ( .IN(n19711), .QN(n19706) );
  INVX0 U20956 ( .IN(n19678), .QN(n19673) );
  INVX0 U20957 ( .IN(n19744), .QN(n19740) );
  INVX0 U20958 ( .IN(n19744), .QN(n19737) );
  INVX0 U20959 ( .IN(n19711), .QN(n19704) );
  INVX0 U20960 ( .IN(n19678), .QN(n19671) );
  INVX0 U20961 ( .IN(n19645), .QN(n19638) );
  INVX0 U20962 ( .IN(n19744), .QN(n19741) );
  INVX0 U20963 ( .IN(n19711), .QN(n19707) );
  INVX0 U20964 ( .IN(n19678), .QN(n19674) );
  INVX0 U20965 ( .IN(n19645), .QN(n19640) );
  INVX0 U20966 ( .IN(n19744), .QN(n19742) );
  INVX0 U20967 ( .IN(n19645), .QN(n19641) );
  INVX0 U20968 ( .IN(n19645), .QN(n19642) );
  INVX0 U20969 ( .IN(n19645), .QN(n19643) );
  INVX0 U20970 ( .IN(n19711), .QN(n19708) );
  INVX0 U20971 ( .IN(n19678), .QN(n19675) );
  INVX0 U20972 ( .IN(n19711), .QN(n19709) );
  INVX0 U20973 ( .IN(n19678), .QN(n19676) );
  INVX0 U20974 ( .IN(n19744), .QN(n19743) );
  INVX0 U20975 ( .IN(n19711), .QN(n19710) );
  INVX0 U20976 ( .IN(n19678), .QN(n19677) );
  INVX0 U20977 ( .IN(n19645), .QN(n19644) );
  INVX0 U20978 ( .IN(n19612), .QN(n19611) );
  INVX0 U20979 ( .IN(n19579), .QN(n19578) );
  INVX0 U20980 ( .IN(n19546), .QN(n19545) );
  INVX0 U20981 ( .IN(n19513), .QN(n19512) );
  INVX0 U20982 ( .IN(n19612), .QN(n19608) );
  INVX0 U20983 ( .IN(n19579), .QN(n19574) );
  INVX0 U20984 ( .IN(n19546), .QN(n19541) );
  INVX0 U20985 ( .IN(n19513), .QN(n19508) );
  INVX0 U20986 ( .IN(n19612), .QN(n19604) );
  INVX0 U20987 ( .IN(n19579), .QN(n19571) );
  INVX0 U20988 ( .IN(n19546), .QN(n19538) );
  INVX0 U20989 ( .IN(n19513), .QN(n19505) );
  INVX0 U20990 ( .IN(n19612), .QN(n19605) );
  INVX0 U20991 ( .IN(n19579), .QN(n19572) );
  INVX0 U20992 ( .IN(n19546), .QN(n19539) );
  INVX0 U20993 ( .IN(n19513), .QN(n19506) );
  INVX0 U20994 ( .IN(n19612), .QN(n19606) );
  INVX0 U20995 ( .IN(n19579), .QN(n19573) );
  INVX0 U20996 ( .IN(n19546), .QN(n19540) );
  INVX0 U20997 ( .IN(n19513), .QN(n19507) );
  INVX0 U20998 ( .IN(n19612), .QN(n19607) );
  INVX0 U20999 ( .IN(n19612), .QN(n19610) );
  INVX0 U21000 ( .IN(n19612), .QN(n19609) );
  INVX0 U21001 ( .IN(n19579), .QN(n19575) );
  INVX0 U21002 ( .IN(n19546), .QN(n19542) );
  INVX0 U21003 ( .IN(n19513), .QN(n19509) );
  INVX0 U21004 ( .IN(n19579), .QN(n19576) );
  INVX0 U21005 ( .IN(n19546), .QN(n19543) );
  INVX0 U21006 ( .IN(n19513), .QN(n19510) );
  INVX0 U21007 ( .IN(n19579), .QN(n19577) );
  INVX0 U21008 ( .IN(n19546), .QN(n19544) );
  INVX0 U21009 ( .IN(n19513), .QN(n19511) );
  INVX0 U21010 ( .IN(n19480), .QN(n19479) );
  INVX0 U21011 ( .IN(n19447), .QN(n19446) );
  INVX0 U21012 ( .IN(n19414), .QN(n19413) );
  INVX0 U21013 ( .IN(n19381), .QN(n19380) );
  INVX0 U21014 ( .IN(n19480), .QN(n19476) );
  INVX0 U21015 ( .IN(n19447), .QN(n19442) );
  INVX0 U21016 ( .IN(n19414), .QN(n19409) );
  INVX0 U21017 ( .IN(n19381), .QN(n19376) );
  INVX0 U21018 ( .IN(n19480), .QN(n19472) );
  INVX0 U21019 ( .IN(n19447), .QN(n19439) );
  INVX0 U21020 ( .IN(n19414), .QN(n19406) );
  INVX0 U21021 ( .IN(n19381), .QN(n19373) );
  INVX0 U21022 ( .IN(n19480), .QN(n19473) );
  INVX0 U21023 ( .IN(n19447), .QN(n19440) );
  INVX0 U21024 ( .IN(n19414), .QN(n19407) );
  INVX0 U21025 ( .IN(n19381), .QN(n19374) );
  INVX0 U21026 ( .IN(n19480), .QN(n19474) );
  INVX0 U21027 ( .IN(n19447), .QN(n19441) );
  INVX0 U21028 ( .IN(n19414), .QN(n19408) );
  INVX0 U21029 ( .IN(n19381), .QN(n19375) );
  INVX0 U21030 ( .IN(n19480), .QN(n19475) );
  INVX0 U21031 ( .IN(n19480), .QN(n19478) );
  INVX0 U21032 ( .IN(n19480), .QN(n19477) );
  INVX0 U21033 ( .IN(n19447), .QN(n19443) );
  INVX0 U21034 ( .IN(n19414), .QN(n19410) );
  INVX0 U21035 ( .IN(n19381), .QN(n19377) );
  INVX0 U21036 ( .IN(n19447), .QN(n19444) );
  INVX0 U21037 ( .IN(n19414), .QN(n19411) );
  INVX0 U21038 ( .IN(n19381), .QN(n19378) );
  INVX0 U21039 ( .IN(n19447), .QN(n19445) );
  INVX0 U21040 ( .IN(n19414), .QN(n19412) );
  INVX0 U21041 ( .IN(n19381), .QN(n19379) );
  INVX0 U21042 ( .IN(n19348), .QN(n19347) );
  INVX0 U21043 ( .IN(n19315), .QN(n19314) );
  INVX0 U21044 ( .IN(n19282), .QN(n19281) );
  INVX0 U21045 ( .IN(n19249), .QN(n19248) );
  INVX0 U21046 ( .IN(n19348), .QN(n19344) );
  INVX0 U21047 ( .IN(n19315), .QN(n19310) );
  INVX0 U21048 ( .IN(n19282), .QN(n19277) );
  INVX0 U21049 ( .IN(n19249), .QN(n19244) );
  INVX0 U21050 ( .IN(n19348), .QN(n19340) );
  INVX0 U21051 ( .IN(n19315), .QN(n19307) );
  INVX0 U21052 ( .IN(n19282), .QN(n19274) );
  INVX0 U21053 ( .IN(n19249), .QN(n19241) );
  INVX0 U21054 ( .IN(n19348), .QN(n19341) );
  INVX0 U21055 ( .IN(n19315), .QN(n19308) );
  INVX0 U21056 ( .IN(n19282), .QN(n19275) );
  INVX0 U21057 ( .IN(n19249), .QN(n19242) );
  INVX0 U21058 ( .IN(n19348), .QN(n19342) );
  INVX0 U21059 ( .IN(n19315), .QN(n19309) );
  INVX0 U21060 ( .IN(n19282), .QN(n19276) );
  INVX0 U21061 ( .IN(n19249), .QN(n19243) );
  INVX0 U21062 ( .IN(n19348), .QN(n19343) );
  INVX0 U21063 ( .IN(n19348), .QN(n19346) );
  INVX0 U21064 ( .IN(n19348), .QN(n19345) );
  INVX0 U21065 ( .IN(n19315), .QN(n19311) );
  INVX0 U21066 ( .IN(n19282), .QN(n19278) );
  INVX0 U21067 ( .IN(n19249), .QN(n19245) );
  INVX0 U21068 ( .IN(n19315), .QN(n19312) );
  INVX0 U21069 ( .IN(n19282), .QN(n19279) );
  INVX0 U21070 ( .IN(n19249), .QN(n19246) );
  INVX0 U21071 ( .IN(n19315), .QN(n19313) );
  INVX0 U21072 ( .IN(n19282), .QN(n19280) );
  INVX0 U21073 ( .IN(n19249), .QN(n19247) );
  INVX0 U21074 ( .IN(n19216), .QN(n19215) );
  INVX0 U21075 ( .IN(n19183), .QN(n19182) );
  INVX0 U21076 ( .IN(n19150), .QN(n19149) );
  INVX0 U21077 ( .IN(n19117), .QN(n19116) );
  INVX0 U21078 ( .IN(n19216), .QN(n19212) );
  INVX0 U21079 ( .IN(n19183), .QN(n19178) );
  INVX0 U21080 ( .IN(n19150), .QN(n19145) );
  INVX0 U21081 ( .IN(n19117), .QN(n19112) );
  INVX0 U21082 ( .IN(n19216), .QN(n19208) );
  INVX0 U21083 ( .IN(n19150), .QN(n19142) );
  INVX0 U21084 ( .IN(n19117), .QN(n19109) );
  INVX0 U21085 ( .IN(n19216), .QN(n19209) );
  INVX0 U21086 ( .IN(n19183), .QN(n19175) );
  INVX0 U21087 ( .IN(n19150), .QN(n19143) );
  INVX0 U21088 ( .IN(n19117), .QN(n19110) );
  INVX0 U21089 ( .IN(n19216), .QN(n19210) );
  INVX0 U21090 ( .IN(n19183), .QN(n19176) );
  INVX0 U21091 ( .IN(n19150), .QN(n19144) );
  INVX0 U21092 ( .IN(n19117), .QN(n19111) );
  INVX0 U21093 ( .IN(n19216), .QN(n19211) );
  INVX0 U21094 ( .IN(n19183), .QN(n19177) );
  INVX0 U21095 ( .IN(n19216), .QN(n19214) );
  INVX0 U21096 ( .IN(n19216), .QN(n19213) );
  INVX0 U21097 ( .IN(n19183), .QN(n19179) );
  INVX0 U21098 ( .IN(n19150), .QN(n19146) );
  INVX0 U21099 ( .IN(n19117), .QN(n19113) );
  INVX0 U21100 ( .IN(n19183), .QN(n19180) );
  INVX0 U21101 ( .IN(n19150), .QN(n19147) );
  INVX0 U21102 ( .IN(n19117), .QN(n19114) );
  INVX0 U21103 ( .IN(n19183), .QN(n19181) );
  INVX0 U21104 ( .IN(n19150), .QN(n19148) );
  INVX0 U21105 ( .IN(n19117), .QN(n19115) );
  INVX0 U21106 ( .IN(n19084), .QN(n19083) );
  INVX0 U21107 ( .IN(n19018), .QN(n19017) );
  INVX0 U21108 ( .IN(n19084), .QN(n19080) );
  INVX0 U21109 ( .IN(n19051), .QN(n19048) );
  INVX0 U21110 ( .IN(n19018), .QN(n19015) );
  INVX0 U21111 ( .IN(n18985), .QN(n18982) );
  INVX0 U21112 ( .IN(n19084), .QN(n19076) );
  INVX0 U21113 ( .IN(n19051), .QN(n19043) );
  INVX0 U21114 ( .IN(n19018), .QN(n19010) );
  INVX0 U21115 ( .IN(n18985), .QN(n18977) );
  INVX0 U21116 ( .IN(n19084), .QN(n19077) );
  INVX0 U21117 ( .IN(n19051), .QN(n19044) );
  INVX0 U21118 ( .IN(n19018), .QN(n19011) );
  INVX0 U21119 ( .IN(n18985), .QN(n18978) );
  INVX0 U21120 ( .IN(n19084), .QN(n19078) );
  INVX0 U21121 ( .IN(n19051), .QN(n19045) );
  INVX0 U21122 ( .IN(n19018), .QN(n19012) );
  INVX0 U21123 ( .IN(n18985), .QN(n18979) );
  INVX0 U21124 ( .IN(n19084), .QN(n19079) );
  INVX0 U21125 ( .IN(n19051), .QN(n19046) );
  INVX0 U21126 ( .IN(n19018), .QN(n19013) );
  INVX0 U21127 ( .IN(n18985), .QN(n18980) );
  INVX0 U21128 ( .IN(n19051), .QN(n19047) );
  INVX0 U21129 ( .IN(n19018), .QN(n19014) );
  INVX0 U21130 ( .IN(n18985), .QN(n18981) );
  INVX0 U21131 ( .IN(n19084), .QN(n19082) );
  INVX0 U21132 ( .IN(n19051), .QN(n19050) );
  INVX0 U21133 ( .IN(n19018), .QN(n19016) );
  INVX0 U21134 ( .IN(n18985), .QN(n18984) );
  INVX0 U21135 ( .IN(n19051), .QN(n19049) );
  INVX0 U21136 ( .IN(n18985), .QN(n18983) );
  INVX0 U21137 ( .IN(n19084), .QN(n19081) );
  INVX0 U21138 ( .IN(n20798), .QN(n20797) );
  INVX0 U21139 ( .IN(n20732), .QN(n20731) );
  INVX0 U21140 ( .IN(n20765), .QN(n20761) );
  INVX0 U21141 ( .IN(n20732), .QN(n20728) );
  INVX0 U21142 ( .IN(n20699), .QN(n20695) );
  INVX0 U21143 ( .IN(n20798), .QN(n20790) );
  INVX0 U21144 ( .IN(n20765), .QN(n20757) );
  INVX0 U21145 ( .IN(n20732), .QN(n20724) );
  INVX0 U21146 ( .IN(n20699), .QN(n20691) );
  INVX0 U21147 ( .IN(n20798), .QN(n20791) );
  INVX0 U21148 ( .IN(n20765), .QN(n20758) );
  INVX0 U21149 ( .IN(n20732), .QN(n20725) );
  INVX0 U21150 ( .IN(n20699), .QN(n20692) );
  INVX0 U21151 ( .IN(n20798), .QN(n20792) );
  INVX0 U21152 ( .IN(n20765), .QN(n20759) );
  INVX0 U21153 ( .IN(n20732), .QN(n20726) );
  INVX0 U21154 ( .IN(n20699), .QN(n20693) );
  INVX0 U21155 ( .IN(n20798), .QN(n20793) );
  INVX0 U21156 ( .IN(n20765), .QN(n20760) );
  INVX0 U21157 ( .IN(n20732), .QN(n20727) );
  INVX0 U21158 ( .IN(n20699), .QN(n20694) );
  INVX0 U21159 ( .IN(n20798), .QN(n20796) );
  INVX0 U21160 ( .IN(n20765), .QN(n20764) );
  INVX0 U21161 ( .IN(n20798), .QN(n20794) );
  INVX0 U21162 ( .IN(n20732), .QN(n20729) );
  INVX0 U21163 ( .IN(n20699), .QN(n20696) );
  INVX0 U21164 ( .IN(n20765), .QN(n20762) );
  INVX0 U21165 ( .IN(n20732), .QN(n20730) );
  INVX0 U21166 ( .IN(n20699), .QN(n20697) );
  INVX0 U21167 ( .IN(n20798), .QN(n20795) );
  INVX0 U21168 ( .IN(n20765), .QN(n20763) );
  INVX0 U21169 ( .IN(n20699), .QN(n20698) );
  INVX0 U21170 ( .IN(n20666), .QN(n20665) );
  INVX0 U21171 ( .IN(n20600), .QN(n20599) );
  INVX0 U21172 ( .IN(n20567), .QN(n20566) );
  INVX0 U21173 ( .IN(n20666), .QN(n20662) );
  INVX0 U21174 ( .IN(n20633), .QN(n20628) );
  INVX0 U21175 ( .IN(n20600), .QN(n20595) );
  INVX0 U21176 ( .IN(n20567), .QN(n20562) );
  INVX0 U21177 ( .IN(n20666), .QN(n20658) );
  INVX0 U21178 ( .IN(n20633), .QN(n20625) );
  INVX0 U21179 ( .IN(n20600), .QN(n20592) );
  INVX0 U21180 ( .IN(n20666), .QN(n20659) );
  INVX0 U21181 ( .IN(n20633), .QN(n20626) );
  INVX0 U21182 ( .IN(n20600), .QN(n20593) );
  INVX0 U21183 ( .IN(n20567), .QN(n20559) );
  INVX0 U21184 ( .IN(n20666), .QN(n20660) );
  INVX0 U21185 ( .IN(n20633), .QN(n20627) );
  INVX0 U21186 ( .IN(n20600), .QN(n20594) );
  INVX0 U21187 ( .IN(n20567), .QN(n20560) );
  INVX0 U21188 ( .IN(n20666), .QN(n20661) );
  INVX0 U21189 ( .IN(n20567), .QN(n20561) );
  INVX0 U21190 ( .IN(n20666), .QN(n20664) );
  INVX0 U21191 ( .IN(n20567), .QN(n20565) );
  INVX0 U21192 ( .IN(n20666), .QN(n20663) );
  INVX0 U21193 ( .IN(n20633), .QN(n20629) );
  INVX0 U21194 ( .IN(n20600), .QN(n20596) );
  INVX0 U21195 ( .IN(n20567), .QN(n20563) );
  INVX0 U21196 ( .IN(n20633), .QN(n20630) );
  INVX0 U21197 ( .IN(n20600), .QN(n20597) );
  INVX0 U21198 ( .IN(n20633), .QN(n20631) );
  INVX0 U21199 ( .IN(n20633), .QN(n20632) );
  INVX0 U21200 ( .IN(n20600), .QN(n20598) );
  INVX0 U21201 ( .IN(n20567), .QN(n20564) );
  INVX0 U21202 ( .IN(n20534), .QN(n20533) );
  INVX0 U21203 ( .IN(n20501), .QN(n20500) );
  INVX0 U21204 ( .IN(n20468), .QN(n20467) );
  INVX0 U21205 ( .IN(n20435), .QN(n20434) );
  INVX0 U21206 ( .IN(n20534), .QN(n20530) );
  INVX0 U21207 ( .IN(n20501), .QN(n20497) );
  INVX0 U21208 ( .IN(n20468), .QN(n20463) );
  INVX0 U21209 ( .IN(n20435), .QN(n20430) );
  INVX0 U21210 ( .IN(n20534), .QN(n20526) );
  INVX0 U21211 ( .IN(n20501), .QN(n20493) );
  INVX0 U21212 ( .IN(n20468), .QN(n20460) );
  INVX0 U21213 ( .IN(n20534), .QN(n20527) );
  INVX0 U21214 ( .IN(n20501), .QN(n20494) );
  INVX0 U21215 ( .IN(n20468), .QN(n20461) );
  INVX0 U21216 ( .IN(n20435), .QN(n20427) );
  INVX0 U21217 ( .IN(n20534), .QN(n20528) );
  INVX0 U21218 ( .IN(n20501), .QN(n20495) );
  INVX0 U21219 ( .IN(n20468), .QN(n20462) );
  INVX0 U21220 ( .IN(n20435), .QN(n20428) );
  INVX0 U21221 ( .IN(n20534), .QN(n20529) );
  INVX0 U21222 ( .IN(n20501), .QN(n20496) );
  INVX0 U21223 ( .IN(n20435), .QN(n20429) );
  INVX0 U21224 ( .IN(n20534), .QN(n20532) );
  INVX0 U21225 ( .IN(n20501), .QN(n20499) );
  INVX0 U21226 ( .IN(n20435), .QN(n20433) );
  INVX0 U21227 ( .IN(n20534), .QN(n20531) );
  INVX0 U21228 ( .IN(n20501), .QN(n20498) );
  INVX0 U21229 ( .IN(n20468), .QN(n20464) );
  INVX0 U21230 ( .IN(n20435), .QN(n20431) );
  INVX0 U21231 ( .IN(n20468), .QN(n20465) );
  INVX0 U21232 ( .IN(n20468), .QN(n20466) );
  INVX0 U21233 ( .IN(n20435), .QN(n20432) );
  INVX0 U21234 ( .IN(n20402), .QN(n20401) );
  INVX0 U21235 ( .IN(n20369), .QN(n20368) );
  INVX0 U21236 ( .IN(n20336), .QN(n20335) );
  INVX0 U21237 ( .IN(n20303), .QN(n20302) );
  INVX0 U21238 ( .IN(n20402), .QN(n20398) );
  INVX0 U21239 ( .IN(n20369), .QN(n20364) );
  INVX0 U21240 ( .IN(n20336), .QN(n20331) );
  INVX0 U21241 ( .IN(n20303), .QN(n20298) );
  INVX0 U21242 ( .IN(n20402), .QN(n20394) );
  INVX0 U21243 ( .IN(n20369), .QN(n20361) );
  INVX0 U21244 ( .IN(n20336), .QN(n20328) );
  INVX0 U21245 ( .IN(n20402), .QN(n20395) );
  INVX0 U21246 ( .IN(n20369), .QN(n20362) );
  INVX0 U21247 ( .IN(n20336), .QN(n20329) );
  INVX0 U21248 ( .IN(n20303), .QN(n20295) );
  INVX0 U21249 ( .IN(n20402), .QN(n20396) );
  INVX0 U21250 ( .IN(n20369), .QN(n20363) );
  INVX0 U21251 ( .IN(n20336), .QN(n20330) );
  INVX0 U21252 ( .IN(n20303), .QN(n20296) );
  INVX0 U21253 ( .IN(n20402), .QN(n20397) );
  INVX0 U21254 ( .IN(n20303), .QN(n20297) );
  INVX0 U21255 ( .IN(n20402), .QN(n20400) );
  INVX0 U21256 ( .IN(n20303), .QN(n20301) );
  INVX0 U21257 ( .IN(n20402), .QN(n20399) );
  INVX0 U21258 ( .IN(n20369), .QN(n20365) );
  INVX0 U21259 ( .IN(n20336), .QN(n20332) );
  INVX0 U21260 ( .IN(n20303), .QN(n20299) );
  INVX0 U21261 ( .IN(n20369), .QN(n20366) );
  INVX0 U21262 ( .IN(n20336), .QN(n20333) );
  INVX0 U21263 ( .IN(n20369), .QN(n20367) );
  INVX0 U21264 ( .IN(n20336), .QN(n20334) );
  INVX0 U21265 ( .IN(n20303), .QN(n20300) );
  INVX0 U21266 ( .IN(n20270), .QN(n20269) );
  INVX0 U21267 ( .IN(n20237), .QN(n20236) );
  INVX0 U21268 ( .IN(n20204), .QN(n20203) );
  INVX0 U21269 ( .IN(n20171), .QN(n20170) );
  INVX0 U21270 ( .IN(n20270), .QN(n20266) );
  INVX0 U21271 ( .IN(n20237), .QN(n20232) );
  INVX0 U21272 ( .IN(n20204), .QN(n20199) );
  INVX0 U21273 ( .IN(n20171), .QN(n20166) );
  INVX0 U21274 ( .IN(n20270), .QN(n20262) );
  INVX0 U21275 ( .IN(n20237), .QN(n20229) );
  INVX0 U21276 ( .IN(n20204), .QN(n20196) );
  INVX0 U21277 ( .IN(n20171), .QN(n20163) );
  INVX0 U21278 ( .IN(n20270), .QN(n20263) );
  INVX0 U21279 ( .IN(n20237), .QN(n20230) );
  INVX0 U21280 ( .IN(n20204), .QN(n20197) );
  INVX0 U21281 ( .IN(n20171), .QN(n20164) );
  INVX0 U21282 ( .IN(n20270), .QN(n20264) );
  INVX0 U21283 ( .IN(n20237), .QN(n20231) );
  INVX0 U21284 ( .IN(n20204), .QN(n20198) );
  INVX0 U21285 ( .IN(n20171), .QN(n20165) );
  INVX0 U21286 ( .IN(n20270), .QN(n20265) );
  INVX0 U21287 ( .IN(n20270), .QN(n20268) );
  INVX0 U21288 ( .IN(n20270), .QN(n20267) );
  INVX0 U21289 ( .IN(n20237), .QN(n20233) );
  INVX0 U21290 ( .IN(n20204), .QN(n20200) );
  INVX0 U21291 ( .IN(n20171), .QN(n20167) );
  INVX0 U21292 ( .IN(n20237), .QN(n20234) );
  INVX0 U21293 ( .IN(n20204), .QN(n20201) );
  INVX0 U21294 ( .IN(n20171), .QN(n20168) );
  INVX0 U21295 ( .IN(n20237), .QN(n20235) );
  INVX0 U21296 ( .IN(n20204), .QN(n20202) );
  INVX0 U21297 ( .IN(n20171), .QN(n20169) );
  INVX0 U21298 ( .IN(n20138), .QN(n20137) );
  INVX0 U21299 ( .IN(n20073), .QN(n20072) );
  INVX0 U21300 ( .IN(n20138), .QN(n20134) );
  INVX0 U21301 ( .IN(n20105), .QN(n20102) );
  INVX0 U21302 ( .IN(n20073), .QN(n20069) );
  INVX0 U21303 ( .IN(n20040), .QN(n20036) );
  INVX0 U21304 ( .IN(n20138), .QN(n20130) );
  INVX0 U21305 ( .IN(n20105), .QN(n20097) );
  INVX0 U21306 ( .IN(n20073), .QN(n20065) );
  INVX0 U21307 ( .IN(n20040), .QN(n20032) );
  INVX0 U21308 ( .IN(n20138), .QN(n20131) );
  INVX0 U21309 ( .IN(n20105), .QN(n20098) );
  INVX0 U21310 ( .IN(n20073), .QN(n20066) );
  INVX0 U21311 ( .IN(n20040), .QN(n20033) );
  INVX0 U21312 ( .IN(n20138), .QN(n20132) );
  INVX0 U21313 ( .IN(n20105), .QN(n20099) );
  INVX0 U21314 ( .IN(n20073), .QN(n20067) );
  INVX0 U21315 ( .IN(n20040), .QN(n20034) );
  INVX0 U21316 ( .IN(n20138), .QN(n20133) );
  INVX0 U21317 ( .IN(n20105), .QN(n20100) );
  INVX0 U21318 ( .IN(n20073), .QN(n20068) );
  INVX0 U21319 ( .IN(n20040), .QN(n20035) );
  INVX0 U21320 ( .IN(n20105), .QN(n20101) );
  INVX0 U21321 ( .IN(n20138), .QN(n20136) );
  INVX0 U21322 ( .IN(n20105), .QN(n20104) );
  INVX0 U21323 ( .IN(n20073), .QN(n20071) );
  INVX0 U21324 ( .IN(n20040), .QN(n20039) );
  INVX0 U21325 ( .IN(n20105), .QN(n20103) );
  INVX0 U21326 ( .IN(n20138), .QN(n20135) );
  INVX0 U21327 ( .IN(n20073), .QN(n20070) );
  INVX0 U21328 ( .IN(n20040), .QN(n20037) );
  INVX0 U21329 ( .IN(n20040), .QN(n20038) );
  INVX0 U21330 ( .IN(n20007), .QN(n20006) );
  INVX0 U21331 ( .IN(n19942), .QN(n19941) );
  INVX0 U21332 ( .IN(n19974), .QN(n19970) );
  INVX0 U21333 ( .IN(n19942), .QN(n19938) );
  INVX0 U21334 ( .IN(n19909), .QN(n19905) );
  INVX0 U21335 ( .IN(n20007), .QN(n19999) );
  INVX0 U21336 ( .IN(n19974), .QN(n19966) );
  INVX0 U21337 ( .IN(n19942), .QN(n19934) );
  INVX0 U21338 ( .IN(n19909), .QN(n19901) );
  INVX0 U21339 ( .IN(n20007), .QN(n20000) );
  INVX0 U21340 ( .IN(n19974), .QN(n19967) );
  INVX0 U21341 ( .IN(n19942), .QN(n19935) );
  INVX0 U21342 ( .IN(n19909), .QN(n19902) );
  INVX0 U21343 ( .IN(n20007), .QN(n20001) );
  INVX0 U21344 ( .IN(n19974), .QN(n19968) );
  INVX0 U21345 ( .IN(n19942), .QN(n19936) );
  INVX0 U21346 ( .IN(n19909), .QN(n19903) );
  INVX0 U21347 ( .IN(n20007), .QN(n20002) );
  INVX0 U21348 ( .IN(n19974), .QN(n19969) );
  INVX0 U21349 ( .IN(n19942), .QN(n19937) );
  INVX0 U21350 ( .IN(n19909), .QN(n19904) );
  INVX0 U21351 ( .IN(n20007), .QN(n20005) );
  INVX0 U21352 ( .IN(n19974), .QN(n19973) );
  INVX0 U21353 ( .IN(n20007), .QN(n20003) );
  INVX0 U21354 ( .IN(n19942), .QN(n19939) );
  INVX0 U21355 ( .IN(n19909), .QN(n19906) );
  INVX0 U21356 ( .IN(n19974), .QN(n19971) );
  INVX0 U21357 ( .IN(n19942), .QN(n19940) );
  INVX0 U21358 ( .IN(n19909), .QN(n19907) );
  INVX0 U21359 ( .IN(n20007), .QN(n20004) );
  INVX0 U21360 ( .IN(n19974), .QN(n19972) );
  INVX0 U21361 ( .IN(n19909), .QN(n19908) );
  INVX0 U21362 ( .IN(n19876), .QN(n19875) );
  INVX0 U21363 ( .IN(n19810), .QN(n19809) );
  INVX0 U21364 ( .IN(n19876), .QN(n19872) );
  INVX0 U21365 ( .IN(n19843), .QN(n19840) );
  INVX0 U21366 ( .IN(n19810), .QN(n19807) );
  INVX0 U21367 ( .IN(n19777), .QN(n19773) );
  INVX0 U21368 ( .IN(n19876), .QN(n19868) );
  INVX0 U21369 ( .IN(n19843), .QN(n19835) );
  INVX0 U21370 ( .IN(n19810), .QN(n19802) );
  INVX0 U21371 ( .IN(n19777), .QN(n19769) );
  INVX0 U21372 ( .IN(n19876), .QN(n19869) );
  INVX0 U21373 ( .IN(n19843), .QN(n19836) );
  INVX0 U21374 ( .IN(n19810), .QN(n19803) );
  INVX0 U21375 ( .IN(n19777), .QN(n19770) );
  INVX0 U21376 ( .IN(n19876), .QN(n19870) );
  INVX0 U21377 ( .IN(n19843), .QN(n19837) );
  INVX0 U21378 ( .IN(n19810), .QN(n19804) );
  INVX0 U21379 ( .IN(n19777), .QN(n19771) );
  INVX0 U21380 ( .IN(n19876), .QN(n19871) );
  INVX0 U21381 ( .IN(n19843), .QN(n19838) );
  INVX0 U21382 ( .IN(n19810), .QN(n19805) );
  INVX0 U21383 ( .IN(n19777), .QN(n19772) );
  INVX0 U21384 ( .IN(n19843), .QN(n19839) );
  INVX0 U21385 ( .IN(n19810), .QN(n19806) );
  INVX0 U21386 ( .IN(n19876), .QN(n19874) );
  INVX0 U21387 ( .IN(n19843), .QN(n19842) );
  INVX0 U21388 ( .IN(n19810), .QN(n19808) );
  INVX0 U21389 ( .IN(n19777), .QN(n19776) );
  INVX0 U21390 ( .IN(n19843), .QN(n19841) );
  INVX0 U21391 ( .IN(n19876), .QN(n19873) );
  INVX0 U21392 ( .IN(n19777), .QN(n19774) );
  INVX0 U21393 ( .IN(n19777), .QN(n19775) );
  INVX0 U21394 ( .IN(n18952), .QN(n18951) );
  INVX0 U21395 ( .IN(n18886), .QN(n18885) );
  INVX0 U21396 ( .IN(n18952), .QN(n18948) );
  INVX0 U21397 ( .IN(n18919), .QN(n18916) );
  INVX0 U21398 ( .IN(n18886), .QN(n18883) );
  INVX0 U21399 ( .IN(n18853), .QN(n18849) );
  INVX0 U21400 ( .IN(n18952), .QN(n18944) );
  INVX0 U21401 ( .IN(n18919), .QN(n18911) );
  INVX0 U21402 ( .IN(n18886), .QN(n18878) );
  INVX0 U21403 ( .IN(n18853), .QN(n18845) );
  INVX0 U21404 ( .IN(n18952), .QN(n18945) );
  INVX0 U21405 ( .IN(n18919), .QN(n18912) );
  INVX0 U21406 ( .IN(n18886), .QN(n18879) );
  INVX0 U21407 ( .IN(n18853), .QN(n18846) );
  INVX0 U21408 ( .IN(n18952), .QN(n18946) );
  INVX0 U21409 ( .IN(n18919), .QN(n18913) );
  INVX0 U21410 ( .IN(n18886), .QN(n18880) );
  INVX0 U21411 ( .IN(n18853), .QN(n18847) );
  INVX0 U21412 ( .IN(n18952), .QN(n18947) );
  INVX0 U21413 ( .IN(n18919), .QN(n18914) );
  INVX0 U21414 ( .IN(n18886), .QN(n18881) );
  INVX0 U21415 ( .IN(n18853), .QN(n18848) );
  INVX0 U21416 ( .IN(n18919), .QN(n18915) );
  INVX0 U21417 ( .IN(n18886), .QN(n18882) );
  INVX0 U21418 ( .IN(n18952), .QN(n18950) );
  INVX0 U21419 ( .IN(n18919), .QN(n18918) );
  INVX0 U21420 ( .IN(n18886), .QN(n18884) );
  INVX0 U21421 ( .IN(n18853), .QN(n18852) );
  INVX0 U21422 ( .IN(n18919), .QN(n18917) );
  INVX0 U21423 ( .IN(n18952), .QN(n18949) );
  INVX0 U21424 ( .IN(n18853), .QN(n18850) );
  INVX0 U21425 ( .IN(n18853), .QN(n18851) );
  INVX0 U21426 ( .IN(n4514), .QN(n20807) );
  INVX0 U21427 ( .IN(n19580), .QN(n19599) );
  INVX0 U21428 ( .IN(n7358), .QN(n19567) );
  INVX0 U21429 ( .IN(n19514), .QN(n19533) );
  INVX0 U21430 ( .IN(n19448), .QN(n19467) );
  INVX0 U21431 ( .IN(n19415), .QN(n19434) );
  INVX0 U21432 ( .IN(n19382), .QN(n19401) );
  INVX0 U21433 ( .IN(n19316), .QN(n19335) );
  INVX0 U21434 ( .IN(n19283), .QN(n19302) );
  INVX0 U21435 ( .IN(n19250), .QN(n19269) );
  INVX0 U21436 ( .IN(n19184), .QN(n19203) );
  INVX0 U21437 ( .IN(n19151), .QN(n19170) );
  INVX0 U21438 ( .IN(n19118), .QN(n19137) );
  INVX0 U21439 ( .IN(n19052), .QN(n19071) );
  INVX0 U21440 ( .IN(n18986), .QN(n19005) );
  INVX0 U21441 ( .IN(n20766), .QN(n20785) );
  INVX0 U21442 ( .IN(n20733), .QN(n20752) );
  INVX0 U21443 ( .IN(n20700), .QN(n20719) );
  INVX0 U21444 ( .IN(n20634), .QN(n20653) );
  INVX0 U21445 ( .IN(n20601), .QN(n20621) );
  INVX0 U21446 ( .IN(n20568), .QN(n20587) );
  INVX0 U21447 ( .IN(n20502), .QN(n20521) );
  INVX0 U21448 ( .IN(n5398), .QN(n20489) );
  INVX0 U21449 ( .IN(n20436), .QN(n20455) );
  INVX0 U21450 ( .IN(n20370), .QN(n20389) );
  INVX0 U21451 ( .IN(n20337), .QN(n20356) );
  INVX0 U21452 ( .IN(n20304), .QN(n20323) );
  INVX0 U21453 ( .IN(n20238), .QN(n20257) );
  INVX0 U21454 ( .IN(n20205), .QN(n20224) );
  INVX0 U21455 ( .IN(n20172), .QN(n20191) );
  INVX0 U21456 ( .IN(n20106), .QN(n20125) );
  INVX0 U21457 ( .IN(n6286), .QN(n20093) );
  INVX0 U21458 ( .IN(n20041), .QN(n20060) );
  INVX0 U21459 ( .IN(n19975), .QN(n19994) );
  INVX0 U21460 ( .IN(n6582), .QN(n19962) );
  INVX0 U21461 ( .IN(n19910), .QN(n19929) );
  INVX0 U21462 ( .IN(n19844), .QN(n19863) );
  INVX0 U21463 ( .IN(n19778), .QN(n19797) );
  INVX0 U21464 ( .IN(n18920), .QN(n18939) );
  INVX0 U21465 ( .IN(n18854), .QN(n18873) );
  INVX0 U21466 ( .IN(n21081), .QN(n21074) );
  INVX0 U21467 ( .IN(n21081), .QN(n21073) );
  INVX0 U21468 ( .IN(n21082), .QN(n21072) );
  INVX0 U21469 ( .IN(n21080), .QN(n21075) );
  INVX0 U21470 ( .IN(n21083), .QN(n21069) );
  INVX0 U21471 ( .IN(n21083), .QN(n21070) );
  INVX0 U21472 ( .IN(n21082), .QN(n21071) );
  INVX0 U21473 ( .IN(n19570), .QN(n19547) );
  INVX0 U21474 ( .IN(n17899), .QN(n19514) );
  INVX0 U21475 ( .IN(n17901), .QN(n19415) );
  INVX0 U21476 ( .IN(n17900), .QN(n19382) );
  INVX0 U21477 ( .IN(n17903), .QN(n19283) );
  INVX0 U21478 ( .IN(n17902), .QN(n19250) );
  INVX0 U21479 ( .IN(n17905), .QN(n19151) );
  INVX0 U21480 ( .IN(n17904), .QN(n19118) );
  INVX0 U21481 ( .IN(n17906), .QN(n18986) );
  INVX0 U21482 ( .IN(n17790), .QN(n19019) );
  INVX0 U21483 ( .IN(n17907), .QN(n20733) );
  INVX0 U21484 ( .IN(n17908), .QN(n20700) );
  INVX0 U21485 ( .IN(n17881), .QN(n20601) );
  INVX0 U21486 ( .IN(n17909), .QN(n20568) );
  INVX0 U21487 ( .IN(n20489), .QN(n20469) );
  INVX0 U21488 ( .IN(n17910), .QN(n20436) );
  INVX0 U21489 ( .IN(n17912), .QN(n20337) );
  INVX0 U21490 ( .IN(n17911), .QN(n20304) );
  INVX0 U21491 ( .IN(n17914), .QN(n20205) );
  INVX0 U21492 ( .IN(n17913), .QN(n20172) );
  INVX0 U21493 ( .IN(n17915), .QN(n20041) );
  INVX0 U21494 ( .IN(n17916), .QN(n19910) );
  INVX0 U21495 ( .IN(n19962), .QN(n19943) );
  INVX0 U21496 ( .IN(n17917), .QN(n19778) );
  INVX0 U21497 ( .IN(n17791), .QN(n19811) );
  INVX0 U21498 ( .IN(n17918), .QN(n18854) );
  INVX0 U21499 ( .IN(n17792), .QN(n18887) );
  INVX0 U21500 ( .IN(n21068), .QN(n21066) );
  INVX0 U21501 ( .IN(n21068), .QN(n21067) );
  INVX0 U21502 ( .IN(n20634), .QN(n20657) );
  INVX0 U21503 ( .IN(n17929), .QN(n20634) );
  INVX0 U21504 ( .IN(n20568), .QN(n20591) );
  INVX0 U21505 ( .IN(n20502), .QN(n20525) );
  INVX0 U21506 ( .IN(n17930), .QN(n20502) );
  INVX0 U21507 ( .IN(n20436), .QN(n20459) );
  INVX0 U21508 ( .IN(n19580), .QN(n19603) );
  INVX0 U21509 ( .IN(n17925), .QN(n19580) );
  INVX0 U21510 ( .IN(n19514), .QN(n19537) );
  INVX0 U21511 ( .IN(n20337), .QN(n20360) );
  INVX0 U21512 ( .IN(n20370), .QN(n20393) );
  INVX0 U21513 ( .IN(n17931), .QN(n20370) );
  INVX0 U21514 ( .IN(n20304), .QN(n20327) );
  INVX0 U21515 ( .IN(n20205), .QN(n20228) );
  INVX0 U21516 ( .IN(n20238), .QN(n20261) );
  INVX0 U21517 ( .IN(n17932), .QN(n20238) );
  INVX0 U21518 ( .IN(n20172), .QN(n20195) );
  INVX0 U21519 ( .IN(n19415), .QN(n19438) );
  INVX0 U21520 ( .IN(n19448), .QN(n19471) );
  INVX0 U21521 ( .IN(n17926), .QN(n19448) );
  INVX0 U21522 ( .IN(n19382), .QN(n19405) );
  INVX0 U21523 ( .IN(n19283), .QN(n19306) );
  INVX0 U21524 ( .IN(n19316), .QN(n19339) );
  INVX0 U21525 ( .IN(n17927), .QN(n19316) );
  INVX0 U21526 ( .IN(n19250), .QN(n19273) );
  INVX0 U21527 ( .IN(n20106), .QN(n20129) );
  INVX0 U21528 ( .IN(n17921), .QN(n20106) );
  INVX0 U21529 ( .IN(n19975), .QN(n19998) );
  INVX0 U21530 ( .IN(n17922), .QN(n19975) );
  INVX0 U21531 ( .IN(n19151), .QN(n19174) );
  INVX0 U21532 ( .IN(n19184), .QN(n19207) );
  INVX0 U21533 ( .IN(n17928), .QN(n19184) );
  INVX0 U21534 ( .IN(n19118), .QN(n19141) );
  INVX0 U21535 ( .IN(n19052), .QN(n19075) );
  INVX0 U21536 ( .IN(n17919), .QN(n19052) );
  INVX0 U21537 ( .IN(n19844), .QN(n19867) );
  INVX0 U21538 ( .IN(n17923), .QN(n19844) );
  INVX0 U21539 ( .IN(n18920), .QN(n18943) );
  INVX0 U21540 ( .IN(n17924), .QN(n18920) );
  INVX0 U21541 ( .IN(n20733), .QN(n20756) );
  INVX0 U21542 ( .IN(n20766), .QN(n20789) );
  INVX0 U21543 ( .IN(n17920), .QN(n20766) );
  NAND2X0 U21544 ( .IN1(n17873), .IN2(n20870), .QN(n4519) );
  NAND2X0 U21545 ( .IN1(n17874), .IN2(n20852), .QN(n4521) );
  NAND2X0 U21546 ( .IN1(n17875), .IN2(n20834), .QN(n4523) );
  NAND2X0 U21547 ( .IN1(n17876), .IN2(n20816), .QN(n4525) );
  NAND2X0 U21548 ( .IN1(n17877), .IN2(n20861), .QN(n4520) );
  NAND2X0 U21549 ( .IN1(n17878), .IN2(n20843), .QN(n4522) );
  NAND2X0 U21550 ( .IN1(n17879), .IN2(n20825), .QN(n4524) );
  NAND2X0 U21551 ( .IN1(n17880), .IN2(n20807), .QN(n4526) );
  NAND2X0 U21552 ( .IN1(n17824), .IN2(n19876), .QN(n6887) );
  NAND2X0 U21553 ( .IN1(n17793), .IN2(n20138), .QN(n6295) );
  NAND2X0 U21554 ( .IN1(n18793), .IN2(n19084), .QN(n8551) );
  NAND2X0 U21555 ( .IN1(n17829), .IN2(n19843), .QN(n6889) );
  NAND2X0 U21556 ( .IN1(n17797), .IN2(n20105), .QN(n6297) );
  NAND2X0 U21557 ( .IN1(n18697), .IN2(n19051), .QN(n8553) );
  NAND2X0 U21558 ( .IN1(n17825), .IN2(n19810), .QN(n6891) );
  NAND2X0 U21559 ( .IN1(n17801), .IN2(n20073), .QN(n6299) );
  NAND2X0 U21560 ( .IN1(n18601), .IN2(n19018), .QN(n8555) );
  NAND2X0 U21561 ( .IN1(n17826), .IN2(n19777), .QN(n6893) );
  NAND2X0 U21562 ( .IN1(n17805), .IN2(n20040), .QN(n6301) );
  NAND2X0 U21563 ( .IN1(n18505), .IN2(n18985), .QN(n8557) );
  NAND2X0 U21564 ( .IN1(n17859), .IN2(n17923), .QN(n6888) );
  NAND2X0 U21565 ( .IN1(n18727), .IN2(n17921), .QN(n6296) );
  NAND2X0 U21566 ( .IN1(n18745), .IN2(n17919), .QN(n8552) );
  NAND2X0 U21567 ( .IN1(n17860), .IN2(n17791), .QN(n6890) );
  NAND2X0 U21568 ( .IN1(n18631), .IN2(n20074), .QN(n6298) );
  NAND2X0 U21569 ( .IN1(n18649), .IN2(n17790), .QN(n8554) );
  NAND2X0 U21570 ( .IN1(n17862), .IN2(n17917), .QN(n6892) );
  NAND2X0 U21571 ( .IN1(n18535), .IN2(n17915), .QN(n6300) );
  NAND2X0 U21572 ( .IN1(n18553), .IN2(n17906), .QN(n8556) );
  NAND2X0 U21573 ( .IN1(n17864), .IN2(n17897), .QN(n6894) );
  NAND2X0 U21574 ( .IN1(n18439), .IN2(n17895), .QN(n6302) );
  NAND2X0 U21575 ( .IN1(n18457), .IN2(n17889), .QN(n8558) );
  NAND2X0 U21576 ( .IN1(n17830), .IN2(n20798), .QN(n4815) );
  NAND2X0 U21577 ( .IN1(n17794), .IN2(n20007), .QN(n6591) );
  NAND2X0 U21578 ( .IN1(n18769), .IN2(n18952), .QN(n8847) );
  NAND2X0 U21579 ( .IN1(n17831), .IN2(n20765), .QN(n4817) );
  NAND2X0 U21580 ( .IN1(n17798), .IN2(n19974), .QN(n6593) );
  NAND2X0 U21581 ( .IN1(n18673), .IN2(n18919), .QN(n8849) );
  NAND2X0 U21582 ( .IN1(n17832), .IN2(n20732), .QN(n4819) );
  NAND2X0 U21583 ( .IN1(n17802), .IN2(n19942), .QN(n6595) );
  NAND2X0 U21584 ( .IN1(n18577), .IN2(n18886), .QN(n8851) );
  NAND2X0 U21585 ( .IN1(n17833), .IN2(n20699), .QN(n4821) );
  NAND2X0 U21586 ( .IN1(n17806), .IN2(n19909), .QN(n6597) );
  NAND2X0 U21587 ( .IN1(n18481), .IN2(n18853), .QN(n8853) );
  NAND2X0 U21588 ( .IN1(n17865), .IN2(n17920), .QN(n4816) );
  NAND2X0 U21589 ( .IN1(n17834), .IN2(n17922), .QN(n6592) );
  NAND2X0 U21590 ( .IN1(n18721), .IN2(n17924), .QN(n8848) );
  NAND2X0 U21591 ( .IN1(n17866), .IN2(n17907), .QN(n4818) );
  NAND2X0 U21592 ( .IN1(n17837), .IN2(n19962), .QN(n6594) );
  NAND2X0 U21593 ( .IN1(n18625), .IN2(n17792), .QN(n8850) );
  NAND2X0 U21594 ( .IN1(n17867), .IN2(n17908), .QN(n4820) );
  NAND2X0 U21595 ( .IN1(n17840), .IN2(n17916), .QN(n6596) );
  NAND2X0 U21596 ( .IN1(n18529), .IN2(n17918), .QN(n8852) );
  NAND2X0 U21597 ( .IN1(n17868), .IN2(n17890), .QN(n4822) );
  NAND2X0 U21598 ( .IN1(n17843), .IN2(n17896), .QN(n6598) );
  NAND2X0 U21599 ( .IN1(n18433), .IN2(n17898), .QN(n8854) );
  NAND2X0 U21600 ( .IN1(n17882), .IN2(n20666), .QN(n5111) );
  NAND2X0 U21601 ( .IN1(n17795), .IN2(n20402), .QN(n5703) );
  NAND2X0 U21602 ( .IN1(n17809), .IN2(n19348), .QN(n7959) );
  NAND2X0 U21603 ( .IN1(n17817), .IN2(n19612), .QN(n7367) );
  NAND2X0 U21604 ( .IN1(n17827), .IN2(n19579), .QN(n7369) );
  NAND2X0 U21605 ( .IN1(n17818), .IN2(n19546), .QN(n7371) );
  NAND2X0 U21606 ( .IN1(n17819), .IN2(n19513), .QN(n7373) );
  NAND2X0 U21607 ( .IN1(n17811), .IN2(n19315), .QN(n7961) );
  NAND2X0 U21608 ( .IN1(n17813), .IN2(n19282), .QN(n7963) );
  NAND2X0 U21609 ( .IN1(n17815), .IN2(n19249), .QN(n7965) );
  NAND2X0 U21610 ( .IN1(n17828), .IN2(n20633), .QN(n5113) );
  NAND2X0 U21611 ( .IN1(n17883), .IN2(n20600), .QN(n5115) );
  NAND2X0 U21612 ( .IN1(n17884), .IN2(n20567), .QN(n5117) );
  NAND2X0 U21613 ( .IN1(n17799), .IN2(n20369), .QN(n5705) );
  NAND2X0 U21614 ( .IN1(n17803), .IN2(n20336), .QN(n5707) );
  NAND2X0 U21615 ( .IN1(n17807), .IN2(n20303), .QN(n5709) );
  NAND2X0 U21616 ( .IN1(n17858), .IN2(n17929), .QN(n5112) );
  NAND2X0 U21617 ( .IN1(n17835), .IN2(n17931), .QN(n5704) );
  NAND2X0 U21618 ( .IN1(n18757), .IN2(n17927), .QN(n7960) );
  NAND2X0 U21619 ( .IN1(n17854), .IN2(n17925), .QN(n7368) );
  NAND2X0 U21620 ( .IN1(n17855), .IN2(n19567), .QN(n7370) );
  NAND2X0 U21621 ( .IN1(n17856), .IN2(n17899), .QN(n7372) );
  NAND2X0 U21622 ( .IN1(n17857), .IN2(n17885), .QN(n7374) );
  NAND2X0 U21623 ( .IN1(n18661), .IN2(n17903), .QN(n7962) );
  NAND2X0 U21624 ( .IN1(n18565), .IN2(n17902), .QN(n7964) );
  NAND2X0 U21625 ( .IN1(n18469), .IN2(n17887), .QN(n7966) );
  NAND2X0 U21626 ( .IN1(n17789), .IN2(n17881), .QN(n5114) );
  NAND2X0 U21627 ( .IN1(n17861), .IN2(n17909), .QN(n5116) );
  NAND2X0 U21628 ( .IN1(n17863), .IN2(n17891), .QN(n5118) );
  NAND2X0 U21629 ( .IN1(n17838), .IN2(n17912), .QN(n5706) );
  NAND2X0 U21630 ( .IN1(n17841), .IN2(n17911), .QN(n5708) );
  NAND2X0 U21631 ( .IN1(n17844), .IN2(n17893), .QN(n5710) );
  NAND2X0 U21632 ( .IN1(n17869), .IN2(n20534), .QN(n5407) );
  NAND2X0 U21633 ( .IN1(n17796), .IN2(n20270), .QN(n5999) );
  NAND2X0 U21634 ( .IN1(n17820), .IN2(n19216), .QN(n8255) );
  NAND2X0 U21635 ( .IN1(n17810), .IN2(n19480), .QN(n7663) );
  NAND2X0 U21636 ( .IN1(n17812), .IN2(n19447), .QN(n7665) );
  NAND2X0 U21637 ( .IN1(n17814), .IN2(n19414), .QN(n7667) );
  NAND2X0 U21638 ( .IN1(n17816), .IN2(n19381), .QN(n7669) );
  NAND2X0 U21639 ( .IN1(n17821), .IN2(n19183), .QN(n8257) );
  NAND2X0 U21640 ( .IN1(n17822), .IN2(n19150), .QN(n8259) );
  NAND2X0 U21641 ( .IN1(n17823), .IN2(n19117), .QN(n8261) );
  NAND2X0 U21642 ( .IN1(n17872), .IN2(n20501), .QN(n5409) );
  NAND2X0 U21643 ( .IN1(n17870), .IN2(n20468), .QN(n5411) );
  NAND2X0 U21644 ( .IN1(n17871), .IN2(n20435), .QN(n5413) );
  NAND2X0 U21645 ( .IN1(n17800), .IN2(n20237), .QN(n6001) );
  NAND2X0 U21646 ( .IN1(n17804), .IN2(n20204), .QN(n6003) );
  NAND2X0 U21647 ( .IN1(n17808), .IN2(n20171), .QN(n6005) );
  NAND2X0 U21648 ( .IN1(n18733), .IN2(n17930), .QN(n5408) );
  NAND2X0 U21649 ( .IN1(n17836), .IN2(n17932), .QN(n6000) );
  NAND2X0 U21650 ( .IN1(n17850), .IN2(n17928), .QN(n8256) );
  NAND2X0 U21651 ( .IN1(n17846), .IN2(n17926), .QN(n7664) );
  NAND2X0 U21652 ( .IN1(n17847), .IN2(n17901), .QN(n7666) );
  NAND2X0 U21653 ( .IN1(n17848), .IN2(n17900), .QN(n7668) );
  NAND2X0 U21654 ( .IN1(n17849), .IN2(n17886), .QN(n7670) );
  NAND2X0 U21655 ( .IN1(n17851), .IN2(n17905), .QN(n8258) );
  NAND2X0 U21656 ( .IN1(n17852), .IN2(n17904), .QN(n8260) );
  NAND2X0 U21657 ( .IN1(n17853), .IN2(n17888), .QN(n8262) );
  NAND2X0 U21658 ( .IN1(n18637), .IN2(n20489), .QN(n5410) );
  NAND2X0 U21659 ( .IN1(n18541), .IN2(n17910), .QN(n5412) );
  NAND2X0 U21660 ( .IN1(n18445), .IN2(n17892), .QN(n5414) );
  NAND2X0 U21661 ( .IN1(n17839), .IN2(n17914), .QN(n6002) );
  NAND2X0 U21662 ( .IN1(n17842), .IN2(n17913), .QN(n6004) );
  NAND2X0 U21663 ( .IN1(n17845), .IN2(n17894), .QN(n6006) );
  INVX0 U21664 ( .IN(n21079), .QN(n21076) );
  INVX0 U21665 ( .IN(n21079), .QN(n21077) );
  NAND2X0 U21666 ( .IN1(n11273), .IN2(n3264), .QN(n11292) );
  NAND2X0 U21667 ( .IN1(n10654), .IN2(n3280), .QN(n10673) );
  NAND2X0 U21668 ( .IN1(n10035), .IN2(n3296), .QN(n10054) );
  NAND2X0 U21669 ( .IN1(n9414), .IN2(n3312), .QN(n9433) );
  NAND2X0 U21670 ( .IN1(n13439), .IN2(n3328), .QN(n13458) );
  NAND2X0 U21671 ( .IN1(n10964), .IN2(n3272), .QN(n10983) );
  NAND2X0 U21672 ( .IN1(n10345), .IN2(n3288), .QN(n10364) );
  NAND2X0 U21673 ( .IN1(n9725), .IN2(n3304), .QN(n9744) );
  NAND3X0 U21674 ( .IN1(n11281), .IN2(n3403), .IN3(n3263), .QN(n11268) );
  NAND3X0 U21675 ( .IN1(n10662), .IN2(n3411), .IN3(n3279), .QN(n10649) );
  NAND3X0 U21676 ( .IN1(n10043), .IN2(n3419), .IN3(n3295), .QN(n10030) );
  NAND3X0 U21677 ( .IN1(n9422), .IN2(n3427), .IN3(n3311), .QN(n9409) );
  NAND3X0 U21678 ( .IN1(n13756), .IN2(n3431), .IN3(n3319), .QN(n13743) );
  NAND3X0 U21679 ( .IN1(n13447), .IN2(n3435), .IN3(n3327), .QN(n13434) );
  NAND3X0 U21680 ( .IN1(n13138), .IN2(n3439), .IN3(n3335), .QN(n13125) );
  NAND3X0 U21681 ( .IN1(n12829), .IN2(n3443), .IN3(n3343), .QN(n12816) );
  NAND3X0 U21682 ( .IN1(n10972), .IN2(n3407), .IN3(n3271), .QN(n10959) );
  NAND3X0 U21683 ( .IN1(n12520), .IN2(n3447), .IN3(n3351), .QN(n12507) );
  NAND3X0 U21684 ( .IN1(n12211), .IN2(n3451), .IN3(n3359), .QN(n12198) );
  NAND3X0 U21685 ( .IN1(n10353), .IN2(n3415), .IN3(n3287), .QN(n10340) );
  NAND3X0 U21686 ( .IN1(n11901), .IN2(n3455), .IN3(n3367), .QN(n11888) );
  NAND3X0 U21687 ( .IN1(n11591), .IN2(n3459), .IN3(n3375), .QN(n11578) );
  NAND3X0 U21688 ( .IN1(n9733), .IN2(n3423), .IN3(n3303), .QN(n9720) );
  NAND3X0 U21689 ( .IN1(n14020), .IN2(n3398), .IN3(n3253), .QN(n14007) );
  NAND3X0 U21690 ( .IN1(n13814), .IN2(n3432), .IN3(n3321), .QN(n13820) );
  NAND3X0 U21691 ( .IN1(n13689), .IN2(n3430), .IN3(n3317), .QN(n13694) );
  NAND3X0 U21692 ( .IN1(n13505), .IN2(n3436), .IN3(n3329), .QN(n13511) );
  NAND3X0 U21693 ( .IN1(n13380), .IN2(n3434), .IN3(n3325), .QN(n13385) );
  NAND3X0 U21694 ( .IN1(n11339), .IN2(n3404), .IN3(n3265), .QN(n11345) );
  NAND3X0 U21695 ( .IN1(n11214), .IN2(n3402), .IN3(n3261), .QN(n11219) );
  NAND3X0 U21696 ( .IN1(n13196), .IN2(n3440), .IN3(n3337), .QN(n13202) );
  NAND3X0 U21697 ( .IN1(n13071), .IN2(n3438), .IN3(n3333), .QN(n13076) );
  NAND3X0 U21698 ( .IN1(n12887), .IN2(n3444), .IN3(n3345), .QN(n12893) );
  NAND3X0 U21699 ( .IN1(n12762), .IN2(n3442), .IN3(n3341), .QN(n12767) );
  NAND3X0 U21700 ( .IN1(n11030), .IN2(n3408), .IN3(n3273), .QN(n11036) );
  NAND3X0 U21701 ( .IN1(n10905), .IN2(n3406), .IN3(n3269), .QN(n10910) );
  NAND3X0 U21702 ( .IN1(n10720), .IN2(n3412), .IN3(n3281), .QN(n10726) );
  NAND3X0 U21703 ( .IN1(n10595), .IN2(n3410), .IN3(n3277), .QN(n10600) );
  NAND3X0 U21704 ( .IN1(n12578), .IN2(n3448), .IN3(n3353), .QN(n12584) );
  NAND3X0 U21705 ( .IN1(n12453), .IN2(n3446), .IN3(n3349), .QN(n12458) );
  NAND3X0 U21706 ( .IN1(n12269), .IN2(n3452), .IN3(n3361), .QN(n12275) );
  NAND3X0 U21707 ( .IN1(n12144), .IN2(n3450), .IN3(n3357), .QN(n12149) );
  NAND3X0 U21708 ( .IN1(n10411), .IN2(n3416), .IN3(n3289), .QN(n10417) );
  NAND3X0 U21709 ( .IN1(n10286), .IN2(n3414), .IN3(n3285), .QN(n10291) );
  NAND3X0 U21710 ( .IN1(n10101), .IN2(n3420), .IN3(n3297), .QN(n10107) );
  NAND3X0 U21711 ( .IN1(n9976), .IN2(n3418), .IN3(n3293), .QN(n9981) );
  NAND3X0 U21712 ( .IN1(n11959), .IN2(n3456), .IN3(n3369), .QN(n11965) );
  NAND3X0 U21713 ( .IN1(n11834), .IN2(n3454), .IN3(n3365), .QN(n11839) );
  NAND3X0 U21714 ( .IN1(n11649), .IN2(n3460), .IN3(n3377), .QN(n11655) );
  NAND3X0 U21715 ( .IN1(n11524), .IN2(n3458), .IN3(n3373), .QN(n11529) );
  NAND3X0 U21716 ( .IN1(n9791), .IN2(n3424), .IN3(n3305), .QN(n9797) );
  NAND3X0 U21717 ( .IN1(n9666), .IN2(n3422), .IN3(n3301), .QN(n9671) );
  NAND3X0 U21718 ( .IN1(n9480), .IN2(n3428), .IN3(n3313), .QN(n9486) );
  NAND3X0 U21719 ( .IN1(n9355), .IN2(n3426), .IN3(n3309), .QN(n9360) );
  OA21X1 U21720 ( .IN1(n13753), .IN2(n13767), .IN3(n13768), .Q(n13762) );
  OA21X1 U21721 ( .IN1(n13135), .IN2(n13149), .IN3(n13150), .Q(n13144) );
  OA21X1 U21722 ( .IN1(n12826), .IN2(n12840), .IN3(n12841), .Q(n12835) );
  OA21X1 U21723 ( .IN1(n12517), .IN2(n12531), .IN3(n12532), .Q(n12526) );
  OA21X1 U21724 ( .IN1(n12208), .IN2(n12222), .IN3(n12223), .Q(n12217) );
  OA21X1 U21725 ( .IN1(n11898), .IN2(n11912), .IN3(n11913), .Q(n11907) );
  OA21X1 U21726 ( .IN1(n11588), .IN2(n11602), .IN3(n11603), .Q(n11597) );
  OA21X1 U21727 ( .IN1(n14017), .IN2(n14031), .IN3(n14032), .Q(n14026) );
  OA21X1 U21728 ( .IN1(n13827), .IN2(n13828), .IN3(n13829), .Q(n13826) );
  OA21X1 U21729 ( .IN1(n13701), .IN2(n13702), .IN3(n13703), .Q(n13700) );
  OA21X1 U21730 ( .IN1(n13518), .IN2(n13519), .IN3(n13520), .Q(n13517) );
  OA21X1 U21731 ( .IN1(n13455), .IN2(n13456), .IN3(n13457), .Q(n13454) );
  OA21X1 U21732 ( .IN1(n13392), .IN2(n13393), .IN3(n13394), .Q(n13391) );
  OA21X1 U21733 ( .IN1(n11352), .IN2(n11353), .IN3(n11354), .Q(n11351) );
  OA21X1 U21734 ( .IN1(n11226), .IN2(n11227), .IN3(n11228), .Q(n11225) );
  OA21X1 U21735 ( .IN1(n13209), .IN2(n13210), .IN3(n13211), .Q(n13208) );
  OA21X1 U21736 ( .IN1(n13083), .IN2(n13084), .IN3(n13085), .Q(n13082) );
  OA21X1 U21737 ( .IN1(n12900), .IN2(n12901), .IN3(n12902), .Q(n12899) );
  OA21X1 U21738 ( .IN1(n12774), .IN2(n12775), .IN3(n12776), .Q(n12773) );
  OA21X1 U21739 ( .IN1(n11043), .IN2(n11044), .IN3(n11045), .Q(n11042) );
  OA21X1 U21740 ( .IN1(n10980), .IN2(n10981), .IN3(n10982), .Q(n10979) );
  OA21X1 U21741 ( .IN1(n10917), .IN2(n10918), .IN3(n10919), .Q(n10916) );
  OA21X1 U21742 ( .IN1(n10733), .IN2(n10734), .IN3(n10735), .Q(n10732) );
  OA21X1 U21743 ( .IN1(n10607), .IN2(n10608), .IN3(n10609), .Q(n10606) );
  OA21X1 U21744 ( .IN1(n12591), .IN2(n12592), .IN3(n12593), .Q(n12590) );
  OA21X1 U21745 ( .IN1(n12465), .IN2(n12466), .IN3(n12467), .Q(n12464) );
  OA21X1 U21746 ( .IN1(n12282), .IN2(n12283), .IN3(n12284), .Q(n12281) );
  OA21X1 U21747 ( .IN1(n12156), .IN2(n12157), .IN3(n12158), .Q(n12155) );
  OA21X1 U21748 ( .IN1(n10424), .IN2(n10425), .IN3(n10426), .Q(n10423) );
  OA21X1 U21749 ( .IN1(n10361), .IN2(n10362), .IN3(n10363), .Q(n10360) );
  OA21X1 U21750 ( .IN1(n10298), .IN2(n10299), .IN3(n10300), .Q(n10297) );
  OA21X1 U21751 ( .IN1(n10114), .IN2(n10115), .IN3(n10116), .Q(n10113) );
  OA21X1 U21752 ( .IN1(n9988), .IN2(n9989), .IN3(n9990), .Q(n9987) );
  OA21X1 U21753 ( .IN1(n11972), .IN2(n11973), .IN3(n11974), .Q(n11971) );
  OA21X1 U21754 ( .IN1(n11846), .IN2(n11847), .IN3(n11848), .Q(n11845) );
  OA21X1 U21755 ( .IN1(n11662), .IN2(n11663), .IN3(n11664), .Q(n11661) );
  OA21X1 U21756 ( .IN1(n11536), .IN2(n11537), .IN3(n11538), .Q(n11535) );
  OA21X1 U21757 ( .IN1(n9804), .IN2(n9805), .IN3(n9806), .Q(n9803) );
  OA21X1 U21758 ( .IN1(n9741), .IN2(n9742), .IN3(n9743), .Q(n9740) );
  OA21X1 U21759 ( .IN1(n9678), .IN2(n9679), .IN3(n9680), .Q(n9677) );
  OA21X1 U21760 ( .IN1(n9493), .IN2(n9494), .IN3(n9495), .Q(n9492) );
  OA21X1 U21761 ( .IN1(n9367), .IN2(n9368), .IN3(n9369), .Q(n9366) );
  OA21X1 U21762 ( .IN1(n11278), .IN2(n11292), .IN3(n11293), .Q(n11287) );
  OA21X1 U21763 ( .IN1(n10659), .IN2(n10673), .IN3(n10674), .Q(n10668) );
  OA21X1 U21764 ( .IN1(n10040), .IN2(n10054), .IN3(n10055), .Q(n10049) );
  OA21X1 U21765 ( .IN1(n9419), .IN2(n9433), .IN3(n9434), .Q(n9428) );
  INVX0 U21766 ( .IN(n13428), .QN(n2986) );
  INVX0 U21767 ( .IN(n10953), .QN(n2874) );
  INVX0 U21768 ( .IN(n10334), .QN(n2906) );
  INVX0 U21769 ( .IN(n9714), .QN(n2938) );
  INVX0 U21770 ( .IN(n13737), .QN(n2970) );
  INVX0 U21771 ( .IN(n11262), .QN(n2858) );
  INVX0 U21772 ( .IN(n13119), .QN(n3002) );
  INVX0 U21773 ( .IN(n12810), .QN(n3018) );
  INVX0 U21774 ( .IN(n10643), .QN(n2890) );
  INVX0 U21775 ( .IN(n12501), .QN(n3034) );
  INVX0 U21776 ( .IN(n12192), .QN(n3050) );
  INVX0 U21777 ( .IN(n10024), .QN(n2922) );
  INVX0 U21778 ( .IN(n11882), .QN(n3066) );
  INVX0 U21779 ( .IN(n11572), .QN(n3082) );
  INVX0 U21780 ( .IN(n9403), .QN(n2954) );
  AOI21X1 U21781 ( .IN1(n4170), .IN2(n11273), .IN3(n11314), .QN(n11293) );
  AOI21X1 U21782 ( .IN1(n4080), .IN2(n10654), .IN3(n10695), .QN(n10674) );
  AOI21X1 U21783 ( .IN1(n3990), .IN2(n10035), .IN3(n10076), .QN(n10055) );
  AOI21X1 U21784 ( .IN1(n3900), .IN2(n9414), .IN3(n9455), .QN(n9434) );
  INVX0 U21785 ( .IN(n13821), .QN(n3145) );
  INVX0 U21786 ( .IN(n13695), .QN(n3142) );
  INVX0 U21787 ( .IN(n13512), .QN(n3151) );
  INVX0 U21788 ( .IN(n13386), .QN(n3148) );
  INVX0 U21789 ( .IN(n11346), .QN(n3103) );
  INVX0 U21790 ( .IN(n11220), .QN(n3100) );
  INVX0 U21791 ( .IN(n13203), .QN(n3157) );
  INVX0 U21792 ( .IN(n13077), .QN(n3154) );
  INVX0 U21793 ( .IN(n12894), .QN(n3163) );
  INVX0 U21794 ( .IN(n12768), .QN(n3160) );
  INVX0 U21795 ( .IN(n11037), .QN(n3109) );
  INVX0 U21796 ( .IN(n10911), .QN(n3106) );
  INVX0 U21797 ( .IN(n10727), .QN(n3115) );
  INVX0 U21798 ( .IN(n10601), .QN(n3112) );
  INVX0 U21799 ( .IN(n12585), .QN(n3169) );
  INVX0 U21800 ( .IN(n12459), .QN(n3166) );
  INVX0 U21801 ( .IN(n12276), .QN(n3175) );
  INVX0 U21802 ( .IN(n12150), .QN(n3172) );
  INVX0 U21803 ( .IN(n10418), .QN(n3121) );
  INVX0 U21804 ( .IN(n10292), .QN(n3118) );
  INVX0 U21805 ( .IN(n10108), .QN(n3127) );
  INVX0 U21806 ( .IN(n9982), .QN(n3124) );
  INVX0 U21807 ( .IN(n11966), .QN(n3181) );
  INVX0 U21808 ( .IN(n11840), .QN(n3178) );
  INVX0 U21809 ( .IN(n11656), .QN(n3187) );
  INVX0 U21810 ( .IN(n11530), .QN(n3184) );
  INVX0 U21811 ( .IN(n9798), .QN(n3133) );
  INVX0 U21812 ( .IN(n9672), .QN(n3130) );
  INVX0 U21813 ( .IN(n9487), .QN(n3139) );
  INVX0 U21814 ( .IN(n9361), .QN(n3136) );
  NAND2X0 U21815 ( .IN1(n2976), .IN2(n13634), .QN(n13843) );
  NAND2X0 U21816 ( .IN1(n2968), .IN2(n13670), .QN(n13714) );
  NAND2X0 U21817 ( .IN1(n2992), .IN2(n13325), .QN(n13534) );
  NAND2X0 U21818 ( .IN1(n2984), .IN2(n13361), .QN(n13405) );
  NAND2X0 U21819 ( .IN1(n2864), .IN2(n11159), .QN(n11368) );
  NAND2X0 U21820 ( .IN1(n2856), .IN2(n11195), .QN(n11239) );
  NAND2X0 U21821 ( .IN1(n3008), .IN2(n13016), .QN(n13225) );
  NAND2X0 U21822 ( .IN1(n3000), .IN2(n13052), .QN(n13096) );
  NAND2X0 U21823 ( .IN1(n3024), .IN2(n12707), .QN(n12916) );
  NAND2X0 U21824 ( .IN1(n3016), .IN2(n12743), .QN(n12787) );
  NAND2X0 U21825 ( .IN1(n2880), .IN2(n10850), .QN(n11059) );
  NAND2X0 U21826 ( .IN1(n2872), .IN2(n10886), .QN(n10930) );
  NAND2X0 U21827 ( .IN1(n2896), .IN2(n10540), .QN(n10749) );
  NAND2X0 U21828 ( .IN1(n2888), .IN2(n10576), .QN(n10620) );
  NAND2X0 U21829 ( .IN1(n3040), .IN2(n12398), .QN(n12607) );
  NAND2X0 U21830 ( .IN1(n3032), .IN2(n12434), .QN(n12478) );
  NAND2X0 U21831 ( .IN1(n3056), .IN2(n12089), .QN(n12298) );
  NAND2X0 U21832 ( .IN1(n3048), .IN2(n12125), .QN(n12169) );
  NAND2X0 U21833 ( .IN1(n2912), .IN2(n10231), .QN(n10440) );
  NAND2X0 U21834 ( .IN1(n2904), .IN2(n10267), .QN(n10311) );
  NAND2X0 U21835 ( .IN1(n2928), .IN2(n9921), .QN(n10130) );
  NAND2X0 U21836 ( .IN1(n2920), .IN2(n9957), .QN(n10001) );
  NAND2X0 U21837 ( .IN1(n3072), .IN2(n11779), .QN(n11988) );
  NAND2X0 U21838 ( .IN1(n3064), .IN2(n11815), .QN(n11859) );
  NAND2X0 U21839 ( .IN1(n3088), .IN2(n11469), .QN(n11678) );
  NAND2X0 U21840 ( .IN1(n3080), .IN2(n11505), .QN(n11549) );
  NAND2X0 U21841 ( .IN1(n2944), .IN2(n9611), .QN(n9820) );
  NAND2X0 U21842 ( .IN1(n2936), .IN2(n9647), .QN(n9691) );
  NAND2X0 U21843 ( .IN1(n2960), .IN2(n9300), .QN(n9509) );
  NAND2X0 U21844 ( .IN1(n2952), .IN2(n9336), .QN(n9380) );
  NAND3X0 U21845 ( .IN1(n13946), .IN2(n3400), .IN3(n3257), .QN(n13953) );
  NAND3X0 U21846 ( .IN1(n14086), .IN2(n3401), .IN3(n3259), .QN(n14093) );
  ISOLANDX1 U21847 ( .D(n13921), .ISO(n3323), .Q(n13922) );
  ISOLANDX1 U21848 ( .D(n13612), .ISO(n3331), .Q(n13613) );
  ISOLANDX1 U21849 ( .D(n11446), .ISO(n3267), .Q(n11447) );
  ISOLANDX1 U21850 ( .D(n13303), .ISO(n3339), .Q(n13304) );
  ISOLANDX1 U21851 ( .D(n12994), .ISO(n3347), .Q(n12995) );
  ISOLANDX1 U21852 ( .D(n11137), .ISO(n3275), .Q(n11138) );
  ISOLANDX1 U21853 ( .D(n10827), .ISO(n3283), .Q(n10828) );
  ISOLANDX1 U21854 ( .D(n12685), .ISO(n3355), .Q(n12686) );
  ISOLANDX1 U21855 ( .D(n12376), .ISO(n3363), .Q(n12377) );
  ISOLANDX1 U21856 ( .D(n10518), .ISO(n3291), .Q(n10519) );
  ISOLANDX1 U21857 ( .D(n10208), .ISO(n3299), .Q(n10209) );
  ISOLANDX1 U21858 ( .D(n12066), .ISO(n3371), .Q(n12067) );
  ISOLANDX1 U21859 ( .D(n11756), .ISO(n3379), .Q(n11757) );
  ISOLANDX1 U21860 ( .D(n9898), .ISO(n3307), .Q(n9899) );
  ISOLANDX1 U21861 ( .D(n9587), .ISO(n3315), .Q(n9588) );
  ISOLANDX1 U21862 ( .D(n14195), .ISO(n3255), .Q(n14196) );
  OA21X1 U21863 ( .IN1(n13812), .IN2(n13634), .IN3(n13813), .Q(n13811) );
  AOI21X1 U21864 ( .IN1(n3322), .IN2(n13814), .IN3(n2976), .QN(n13812) );
  OA21X1 U21865 ( .IN1(n13687), .IN2(n13670), .IN3(n13688), .Q(n13686) );
  AOI21X1 U21866 ( .IN1(n3318), .IN2(n13689), .IN3(n2968), .QN(n13687) );
  OA21X1 U21867 ( .IN1(n13503), .IN2(n13325), .IN3(n13504), .Q(n13502) );
  AOI21X1 U21868 ( .IN1(n3330), .IN2(n13505), .IN3(n2992), .QN(n13503) );
  OA21X1 U21869 ( .IN1(n13378), .IN2(n13361), .IN3(n13379), .Q(n13377) );
  AOI21X1 U21870 ( .IN1(n3326), .IN2(n13380), .IN3(n2984), .QN(n13378) );
  OA21X1 U21871 ( .IN1(n11337), .IN2(n11159), .IN3(n11338), .Q(n11336) );
  AOI21X1 U21872 ( .IN1(n3266), .IN2(n11339), .IN3(n2864), .QN(n11337) );
  OA21X1 U21873 ( .IN1(n11212), .IN2(n11195), .IN3(n11213), .Q(n11211) );
  AOI21X1 U21874 ( .IN1(n3262), .IN2(n11214), .IN3(n2856), .QN(n11212) );
  OA21X1 U21875 ( .IN1(n13194), .IN2(n13016), .IN3(n13195), .Q(n13193) );
  AOI21X1 U21876 ( .IN1(n3338), .IN2(n13196), .IN3(n3008), .QN(n13194) );
  OA21X1 U21877 ( .IN1(n13069), .IN2(n13052), .IN3(n13070), .Q(n13068) );
  AOI21X1 U21878 ( .IN1(n3334), .IN2(n13071), .IN3(n3000), .QN(n13069) );
  OA21X1 U21879 ( .IN1(n12885), .IN2(n12707), .IN3(n12886), .Q(n12884) );
  AOI21X1 U21880 ( .IN1(n3346), .IN2(n12887), .IN3(n3024), .QN(n12885) );
  OA21X1 U21881 ( .IN1(n12760), .IN2(n12743), .IN3(n12761), .Q(n12759) );
  AOI21X1 U21882 ( .IN1(n3342), .IN2(n12762), .IN3(n3016), .QN(n12760) );
  OA21X1 U21883 ( .IN1(n11028), .IN2(n10850), .IN3(n11029), .Q(n11027) );
  AOI21X1 U21884 ( .IN1(n3274), .IN2(n11030), .IN3(n2880), .QN(n11028) );
  OA21X1 U21885 ( .IN1(n10903), .IN2(n10886), .IN3(n10904), .Q(n10902) );
  AOI21X1 U21886 ( .IN1(n3270), .IN2(n10905), .IN3(n2872), .QN(n10903) );
  OA21X1 U21887 ( .IN1(n10718), .IN2(n10540), .IN3(n10719), .Q(n10717) );
  AOI21X1 U21888 ( .IN1(n3282), .IN2(n10720), .IN3(n2896), .QN(n10718) );
  OA21X1 U21889 ( .IN1(n10593), .IN2(n10576), .IN3(n10594), .Q(n10592) );
  AOI21X1 U21890 ( .IN1(n3278), .IN2(n10595), .IN3(n2888), .QN(n10593) );
  OA21X1 U21891 ( .IN1(n12576), .IN2(n12398), .IN3(n12577), .Q(n12575) );
  AOI21X1 U21892 ( .IN1(n3354), .IN2(n12578), .IN3(n3040), .QN(n12576) );
  OA21X1 U21893 ( .IN1(n12451), .IN2(n12434), .IN3(n12452), .Q(n12450) );
  AOI21X1 U21894 ( .IN1(n3350), .IN2(n12453), .IN3(n3032), .QN(n12451) );
  OA21X1 U21895 ( .IN1(n12267), .IN2(n12089), .IN3(n12268), .Q(n12266) );
  AOI21X1 U21896 ( .IN1(n3362), .IN2(n12269), .IN3(n3056), .QN(n12267) );
  OA21X1 U21897 ( .IN1(n12142), .IN2(n12125), .IN3(n12143), .Q(n12141) );
  AOI21X1 U21898 ( .IN1(n3358), .IN2(n12144), .IN3(n3048), .QN(n12142) );
  OA21X1 U21899 ( .IN1(n10409), .IN2(n10231), .IN3(n10410), .Q(n10408) );
  AOI21X1 U21900 ( .IN1(n3290), .IN2(n10411), .IN3(n2912), .QN(n10409) );
  OA21X1 U21901 ( .IN1(n10284), .IN2(n10267), .IN3(n10285), .Q(n10283) );
  AOI21X1 U21902 ( .IN1(n3286), .IN2(n10286), .IN3(n2904), .QN(n10284) );
  OA21X1 U21903 ( .IN1(n10099), .IN2(n9921), .IN3(n10100), .Q(n10098) );
  AOI21X1 U21904 ( .IN1(n3298), .IN2(n10101), .IN3(n2928), .QN(n10099) );
  OA21X1 U21905 ( .IN1(n9974), .IN2(n9957), .IN3(n9975), .Q(n9973) );
  AOI21X1 U21906 ( .IN1(n3294), .IN2(n9976), .IN3(n2920), .QN(n9974) );
  OA21X1 U21907 ( .IN1(n11957), .IN2(n11779), .IN3(n11958), .Q(n11956) );
  AOI21X1 U21908 ( .IN1(n3370), .IN2(n11959), .IN3(n3072), .QN(n11957) );
  OA21X1 U21909 ( .IN1(n11832), .IN2(n11815), .IN3(n11833), .Q(n11831) );
  AOI21X1 U21910 ( .IN1(n3366), .IN2(n11834), .IN3(n3064), .QN(n11832) );
  OA21X1 U21911 ( .IN1(n11647), .IN2(n11469), .IN3(n11648), .Q(n11646) );
  AOI21X1 U21912 ( .IN1(n3378), .IN2(n11649), .IN3(n3088), .QN(n11647) );
  OA21X1 U21913 ( .IN1(n11522), .IN2(n11505), .IN3(n11523), .Q(n11521) );
  AOI21X1 U21914 ( .IN1(n3374), .IN2(n11524), .IN3(n3080), .QN(n11522) );
  OA21X1 U21915 ( .IN1(n9789), .IN2(n9611), .IN3(n9790), .Q(n9788) );
  AOI21X1 U21916 ( .IN1(n3306), .IN2(n9791), .IN3(n2944), .QN(n9789) );
  OA21X1 U21917 ( .IN1(n9664), .IN2(n9647), .IN3(n9665), .Q(n9663) );
  AOI21X1 U21918 ( .IN1(n3302), .IN2(n9666), .IN3(n2936), .QN(n9664) );
  OA21X1 U21919 ( .IN1(n9478), .IN2(n9300), .IN3(n9479), .Q(n9477) );
  AOI21X1 U21920 ( .IN1(n3314), .IN2(n9480), .IN3(n2960), .QN(n9478) );
  OA21X1 U21921 ( .IN1(n9353), .IN2(n9336), .IN3(n9354), .Q(n9352) );
  AOI21X1 U21922 ( .IN1(n3310), .IN2(n9355), .IN3(n2952), .QN(n9353) );
  OA21X1 U21923 ( .IN1(n13895), .IN2(n13896), .IN3(n13897), .Q(n13893) );
  OA21X1 U21924 ( .IN1(n13586), .IN2(n13587), .IN3(n13588), .Q(n13584) );
  OA21X1 U21925 ( .IN1(n11420), .IN2(n11421), .IN3(n11422), .Q(n11418) );
  OA21X1 U21926 ( .IN1(n13277), .IN2(n13278), .IN3(n13279), .Q(n13275) );
  OA21X1 U21927 ( .IN1(n12968), .IN2(n12969), .IN3(n12970), .Q(n12966) );
  OA21X1 U21928 ( .IN1(n11111), .IN2(n11112), .IN3(n11113), .Q(n11109) );
  OA21X1 U21929 ( .IN1(n10801), .IN2(n10802), .IN3(n10803), .Q(n10799) );
  OA21X1 U21930 ( .IN1(n12659), .IN2(n12660), .IN3(n12661), .Q(n12657) );
  OA21X1 U21931 ( .IN1(n12350), .IN2(n12351), .IN3(n12352), .Q(n12348) );
  OA21X1 U21932 ( .IN1(n10492), .IN2(n10493), .IN3(n10494), .Q(n10490) );
  OA21X1 U21933 ( .IN1(n10182), .IN2(n10183), .IN3(n10184), .Q(n10180) );
  OA21X1 U21934 ( .IN1(n12040), .IN2(n12041), .IN3(n12042), .Q(n12038) );
  OA21X1 U21935 ( .IN1(n11730), .IN2(n11731), .IN3(n11732), .Q(n11728) );
  OA21X1 U21936 ( .IN1(n9872), .IN2(n9873), .IN3(n9874), .Q(n9870) );
  OA21X1 U21937 ( .IN1(n9561), .IN2(n9562), .IN3(n9563), .Q(n9559) );
  OA21X1 U21938 ( .IN1(n13960), .IN2(n13961), .IN3(n13962), .Q(n13959) );
  OA21X1 U21939 ( .IN1(n14169), .IN2(n14170), .IN3(n14171), .Q(n14167) );
  OA21X1 U21940 ( .IN1(n14100), .IN2(n14101), .IN3(n14102), .Q(n14099) );
  OA21X1 U21941 ( .IN1(n2979), .IN2(n13915), .IN3(n13916), .Q(n13908) );
  OA21X1 U21942 ( .IN1(n3433), .IN2(n13898), .IN3(n13895), .Q(n13915) );
  OA21X1 U21943 ( .IN1(n2995), .IN2(n13606), .IN3(n13607), .Q(n13599) );
  OA21X1 U21944 ( .IN1(n3437), .IN2(n13589), .IN3(n13586), .Q(n13606) );
  OA21X1 U21945 ( .IN1(n2867), .IN2(n11440), .IN3(n11441), .Q(n11433) );
  OA21X1 U21946 ( .IN1(n3405), .IN2(n11423), .IN3(n11420), .Q(n11440) );
  OA21X1 U21947 ( .IN1(n3011), .IN2(n13297), .IN3(n13298), .Q(n13290) );
  OA21X1 U21948 ( .IN1(n3441), .IN2(n13280), .IN3(n13277), .Q(n13297) );
  OA21X1 U21949 ( .IN1(n3027), .IN2(n12988), .IN3(n12989), .Q(n12981) );
  OA21X1 U21950 ( .IN1(n3445), .IN2(n12971), .IN3(n12968), .Q(n12988) );
  OA21X1 U21951 ( .IN1(n2883), .IN2(n11131), .IN3(n11132), .Q(n11124) );
  OA21X1 U21952 ( .IN1(n3409), .IN2(n11114), .IN3(n11111), .Q(n11131) );
  OA21X1 U21953 ( .IN1(n2899), .IN2(n10821), .IN3(n10822), .Q(n10814) );
  OA21X1 U21954 ( .IN1(n3413), .IN2(n10804), .IN3(n10801), .Q(n10821) );
  OA21X1 U21955 ( .IN1(n3043), .IN2(n12679), .IN3(n12680), .Q(n12672) );
  OA21X1 U21956 ( .IN1(n3449), .IN2(n12662), .IN3(n12659), .Q(n12679) );
  OA21X1 U21957 ( .IN1(n3059), .IN2(n12370), .IN3(n12371), .Q(n12363) );
  OA21X1 U21958 ( .IN1(n3453), .IN2(n12353), .IN3(n12350), .Q(n12370) );
  OA21X1 U21959 ( .IN1(n2915), .IN2(n10512), .IN3(n10513), .Q(n10505) );
  OA21X1 U21960 ( .IN1(n3417), .IN2(n10495), .IN3(n10492), .Q(n10512) );
  OA21X1 U21961 ( .IN1(n2931), .IN2(n10202), .IN3(n10203), .Q(n10195) );
  OA21X1 U21962 ( .IN1(n3421), .IN2(n10185), .IN3(n10182), .Q(n10202) );
  OA21X1 U21963 ( .IN1(n3075), .IN2(n12060), .IN3(n12061), .Q(n12053) );
  OA21X1 U21964 ( .IN1(n3457), .IN2(n12043), .IN3(n12040), .Q(n12060) );
  OA21X1 U21965 ( .IN1(n3091), .IN2(n11750), .IN3(n11751), .Q(n11743) );
  OA21X1 U21966 ( .IN1(n3461), .IN2(n11733), .IN3(n11730), .Q(n11750) );
  OA21X1 U21967 ( .IN1(n2947), .IN2(n9892), .IN3(n9893), .Q(n9885) );
  OA21X1 U21968 ( .IN1(n3425), .IN2(n9875), .IN3(n9872), .Q(n9892) );
  OA21X1 U21969 ( .IN1(n2963), .IN2(n9581), .IN3(n9582), .Q(n9574) );
  OA21X1 U21970 ( .IN1(n3429), .IN2(n9564), .IN3(n9561), .Q(n9581) );
  OA21X1 U21971 ( .IN1(n2842), .IN2(n14189), .IN3(n14190), .Q(n14182) );
  OA21X1 U21972 ( .IN1(n3399), .IN2(n14172), .IN3(n14169), .Q(n14189) );
  NAND3X0 U21973 ( .IN1(n3433), .IN2(n13887), .IN3(n3324), .QN(n13878) );
  NAND3X0 U21974 ( .IN1(n3437), .IN2(n13578), .IN3(n3332), .QN(n13569) );
  NAND3X0 U21975 ( .IN1(n3405), .IN2(n11412), .IN3(n3268), .QN(n11403) );
  NAND3X0 U21976 ( .IN1(n3441), .IN2(n13269), .IN3(n3340), .QN(n13260) );
  NAND3X0 U21977 ( .IN1(n3445), .IN2(n12960), .IN3(n3348), .QN(n12951) );
  NAND3X0 U21978 ( .IN1(n3409), .IN2(n11103), .IN3(n3276), .QN(n11094) );
  NAND3X0 U21979 ( .IN1(n3413), .IN2(n10793), .IN3(n3284), .QN(n10784) );
  NAND3X0 U21980 ( .IN1(n3449), .IN2(n12651), .IN3(n3356), .QN(n12642) );
  NAND3X0 U21981 ( .IN1(n3453), .IN2(n12342), .IN3(n3364), .QN(n12333) );
  NAND3X0 U21982 ( .IN1(n3417), .IN2(n10484), .IN3(n3292), .QN(n10475) );
  NAND3X0 U21983 ( .IN1(n3421), .IN2(n10174), .IN3(n3300), .QN(n10165) );
  NAND3X0 U21984 ( .IN1(n3457), .IN2(n12032), .IN3(n3372), .QN(n12023) );
  NAND3X0 U21985 ( .IN1(n3461), .IN2(n11722), .IN3(n3380), .QN(n11713) );
  NAND3X0 U21986 ( .IN1(n3425), .IN2(n9864), .IN3(n3308), .QN(n9855) );
  NAND3X0 U21987 ( .IN1(n3429), .IN2(n9553), .IN3(n3316), .QN(n9544) );
  NAND3X0 U21988 ( .IN1(n3399), .IN2(n14161), .IN3(n3256), .QN(n14152) );
  AOI21X1 U21989 ( .IN1(n3879), .IN2(n13880), .IN3(n13918), .QN(n13899) );
  AOI21X1 U21990 ( .IN1(n3834), .IN2(n13571), .IN3(n13609), .QN(n13590) );
  AOI21X1 U21991 ( .IN1(n4194), .IN2(n11405), .IN3(n11443), .QN(n11424) );
  AOI21X1 U21992 ( .IN1(n3789), .IN2(n13262), .IN3(n13300), .QN(n13281) );
  AOI21X1 U21993 ( .IN1(n3744), .IN2(n12953), .IN3(n12991), .QN(n12972) );
  AOI21X1 U21994 ( .IN1(n4149), .IN2(n11096), .IN3(n11134), .QN(n11115) );
  AOI21X1 U21995 ( .IN1(n4104), .IN2(n10786), .IN3(n10824), .QN(n10805) );
  AOI21X1 U21996 ( .IN1(n3699), .IN2(n12644), .IN3(n12682), .QN(n12663) );
  AOI21X1 U21997 ( .IN1(n3654), .IN2(n12335), .IN3(n12373), .QN(n12354) );
  AOI21X1 U21998 ( .IN1(n4059), .IN2(n10477), .IN3(n10515), .QN(n10496) );
  AOI21X1 U21999 ( .IN1(n4014), .IN2(n10167), .IN3(n10205), .QN(n10186) );
  AOI21X1 U22000 ( .IN1(n3609), .IN2(n12025), .IN3(n12063), .QN(n12044) );
  AOI21X1 U22001 ( .IN1(n3564), .IN2(n11715), .IN3(n11753), .QN(n11734) );
  AOI21X1 U22002 ( .IN1(n3969), .IN2(n9857), .IN3(n9895), .QN(n9876) );
  AOI21X1 U22003 ( .IN1(n3924), .IN2(n9546), .IN3(n9584), .QN(n9565) );
  AOI21X1 U22004 ( .IN1(n4239), .IN2(n14154), .IN3(n14192), .QN(n14173) );
  INVX0 U22005 ( .IN(n13954), .QN(n3096) );
  INVX0 U22006 ( .IN(n14094), .QN(n3098) );
  INVX0 U22007 ( .IN(n13898), .QN(n3324) );
  INVX0 U22008 ( .IN(n13589), .QN(n3332) );
  INVX0 U22009 ( .IN(n11423), .QN(n3268) );
  INVX0 U22010 ( .IN(n12662), .QN(n3356) );
  INVX0 U22011 ( .IN(n12353), .QN(n3364) );
  INVX0 U22012 ( .IN(n9875), .QN(n3308) );
  INVX0 U22013 ( .IN(n14172), .QN(n3256) );
  INVX0 U22014 ( .IN(n14103), .QN(n3259) );
  OA21X1 U22015 ( .IN1(n14084), .IN2(n3382), .IN3(n14085), .Q(n14083) );
  AOI21X1 U22016 ( .IN1(n3260), .IN2(n14086), .IN3(n2851), .QN(n14084) );
  INVX0 U22017 ( .IN(n13868), .QN(n2977) );
  INVX0 U22018 ( .IN(n13559), .QN(n2993) );
  INVX0 U22019 ( .IN(n11393), .QN(n2865) );
  INVX0 U22020 ( .IN(n12632), .QN(n3041) );
  INVX0 U22021 ( .IN(n12323), .QN(n3057) );
  INVX0 U22022 ( .IN(n9845), .QN(n2945) );
  INVX0 U22023 ( .IN(n14142), .QN(n2840) );
  INVX0 U22024 ( .IN(n14076), .QN(n2848) );
  OR2X1 U22025 ( .IN1(n13881), .IN2(n3390), .Q(n13910) );
  OR2X1 U22026 ( .IN1(n13572), .IN2(n3391), .Q(n13601) );
  OR2X1 U22027 ( .IN1(n11406), .IN2(n3383), .Q(n11435) );
  OR2X1 U22028 ( .IN1(n13263), .IN2(n3392), .Q(n13292) );
  OR2X1 U22029 ( .IN1(n12954), .IN2(n3393), .Q(n12983) );
  OR2X1 U22030 ( .IN1(n11097), .IN2(n3384), .Q(n11126) );
  OR2X1 U22031 ( .IN1(n10787), .IN2(n3385), .Q(n10816) );
  OR2X1 U22032 ( .IN1(n12645), .IN2(n3394), .Q(n12674) );
  OR2X1 U22033 ( .IN1(n12336), .IN2(n3395), .Q(n12365) );
  OR2X1 U22034 ( .IN1(n10478), .IN2(n3386), .Q(n10507) );
  OR2X1 U22035 ( .IN1(n10168), .IN2(n3387), .Q(n10197) );
  OR2X1 U22036 ( .IN1(n12026), .IN2(n3396), .Q(n12055) );
  OR2X1 U22037 ( .IN1(n11716), .IN2(n3397), .Q(n11745) );
  OR2X1 U22038 ( .IN1(n9858), .IN2(n3388), .Q(n9887) );
  OR2X1 U22039 ( .IN1(n9547), .IN2(n3389), .Q(n9576) );
  INVX0 U22040 ( .IN(n19717), .QN(n19712) );
  INVX0 U22041 ( .IN(n7172), .QN(n19717) );
  INVX0 U22042 ( .IN(n19651), .QN(n19646) );
  INVX0 U22043 ( .IN(n7176), .QN(n19651) );
  INVX0 U22044 ( .IN(n7174), .QN(n19682) );
  INVX0 U22045 ( .IN(n7172), .QN(n19715) );
  INVX0 U22046 ( .IN(n7176), .QN(n19649) );
  INVX0 U22047 ( .IN(n19684), .QN(n19679) );
  INVX0 U22048 ( .IN(n7174), .QN(n19684) );
  NAND3X0 U22049 ( .IN1(n4205), .IN2(n4210), .IN3(n4211), .QN(n7178) );
  NOR2X0 U22050 ( .IN1(s15_addr_o[3]), .IN2(s15_addr_o[4]), .QN(n9601) );
  NOR2X0 U22051 ( .IN1(s15_addr_o[2]), .IN2(s15_addr_o[5]), .QN(n11770) );
  NOR2X0 U22052 ( .IN1(n1698), .IN2(s15_addr_o[4]), .QN(n10222) );
  NOR2X0 U22053 ( .IN1(n1700), .IN2(s15_addr_o[5]), .QN(n12080) );
  INVX0 U22054 ( .IN(s15_addr_o[2]), .QN(n1700) );
  INVX0 U22055 ( .IN(s15_addr_o[3]), .QN(n1698) );
  ISOLANDX1 U22056 ( .D(s15_addr_o[5]), .ISO(n1700), .Q(n9912) );
  ISOLANDX1 U22057 ( .D(s15_addr_o[5]), .ISO(s15_addr_o[2]), .Q(n9602) );
  ISOLANDX1 U22058 ( .D(s15_addr_o[4]), .ISO(n1698), .Q(n11460) );
  ISOLANDX1 U22059 ( .D(s15_addr_o[4]), .ISO(s15_addr_o[3]), .Q(n10841) );
  INVX0 U22060 ( .IN(n14208), .QN(n1692) );
  INVX0 U22061 ( .IN(n11459), .QN(n1680) );
  INVX0 U22062 ( .IN(n11150), .QN(n1693) );
  INVX0 U22063 ( .IN(n10840), .QN(n1681) );
  INVX0 U22064 ( .IN(n10531), .QN(n1694) );
  INVX0 U22065 ( .IN(n10221), .QN(n1682) );
  INVX0 U22066 ( .IN(n9911), .QN(n1695) );
  INVX0 U22067 ( .IN(n9600), .QN(n1683) );
  INVX0 U22068 ( .IN(n13934), .QN(n1688) );
  INVX0 U22069 ( .IN(n13625), .QN(n1684) );
  INVX0 U22070 ( .IN(n13316), .QN(n1689) );
  INVX0 U22071 ( .IN(n13007), .QN(n1685) );
  INVX0 U22072 ( .IN(n12698), .QN(n1690) );
  INVX0 U22073 ( .IN(n12389), .QN(n1686) );
  INVX0 U22074 ( .IN(n12079), .QN(n1691) );
  INVX0 U22075 ( .IN(n11769), .QN(n1687) );
  INVX0 U22076 ( .IN(n7173), .QN(n19711) );
  INVX0 U22077 ( .IN(n7171), .QN(n19744) );
  INVX0 U22078 ( .IN(n7175), .QN(n19678) );
  INVX0 U22079 ( .IN(n7177), .QN(n19645) );
  INVX0 U22080 ( .IN(n7174), .QN(n19683) );
  INVX0 U22081 ( .IN(n7176), .QN(n19650) );
  INVX0 U22082 ( .IN(n7172), .QN(n19716) );
  NBUFFX2 U22083 ( .IN(n14208), .Q(n18337) );
  NBUFFX2 U22084 ( .IN(n14208), .Q(n18336) );
  NBUFFX2 U22085 ( .IN(n11459), .Q(n18405) );
  NBUFFX2 U22086 ( .IN(n11459), .Q(n18404) );
  NBUFFX2 U22087 ( .IN(n11150), .Q(n18409) );
  NBUFFX2 U22088 ( .IN(n11150), .Q(n18408) );
  NBUFFX2 U22089 ( .IN(n10840), .Q(n18413) );
  NBUFFX2 U22090 ( .IN(n10840), .Q(n18412) );
  NBUFFX2 U22091 ( .IN(n10531), .Q(n18417) );
  NBUFFX2 U22092 ( .IN(n10531), .Q(n18416) );
  NBUFFX2 U22093 ( .IN(n10221), .Q(n18421) );
  NBUFFX2 U22094 ( .IN(n10221), .Q(n18420) );
  NBUFFX2 U22095 ( .IN(n9911), .Q(n18425) );
  NBUFFX2 U22096 ( .IN(n9911), .Q(n18424) );
  NBUFFX2 U22097 ( .IN(n9600), .Q(n18429) );
  NBUFFX2 U22098 ( .IN(n9600), .Q(n18428) );
  NBUFFX2 U22099 ( .IN(n13934), .Q(n18373) );
  NBUFFX2 U22100 ( .IN(n13934), .Q(n18372) );
  NBUFFX2 U22101 ( .IN(n13625), .Q(n18377) );
  NBUFFX2 U22102 ( .IN(n13625), .Q(n18376) );
  NBUFFX2 U22103 ( .IN(n13316), .Q(n18381) );
  NBUFFX2 U22104 ( .IN(n13316), .Q(n18380) );
  NBUFFX2 U22105 ( .IN(n13007), .Q(n18385) );
  NBUFFX2 U22106 ( .IN(n13007), .Q(n18384) );
  OR2X1 U22107 ( .IN1(n14155), .IN2(n3381), .Q(n14184) );
  NAND2X0 U22108 ( .IN1(n2851), .IN2(n3382), .QN(n14116) );
  NAND3X0 U22109 ( .IN1(n3935), .IN2(n3940), .IN3(n3941), .QN(n4514) );
  INVX0 U22110 ( .IN(n7357), .QN(n19579) );
  INVX0 U22111 ( .IN(n7359), .QN(n19546) );
  INVX0 U22112 ( .IN(n7361), .QN(n19513) );
  INVX0 U22113 ( .IN(n7355), .QN(n19612) );
  INVX0 U22114 ( .IN(n7653), .QN(n19447) );
  INVX0 U22115 ( .IN(n7655), .QN(n19414) );
  INVX0 U22116 ( .IN(n7657), .QN(n19381) );
  INVX0 U22117 ( .IN(n7651), .QN(n19480) );
  INVX0 U22118 ( .IN(n7949), .QN(n19315) );
  INVX0 U22119 ( .IN(n7951), .QN(n19282) );
  INVX0 U22120 ( .IN(n7953), .QN(n19249) );
  INVX0 U22121 ( .IN(n7947), .QN(n19348) );
  INVX0 U22122 ( .IN(n8245), .QN(n19183) );
  INVX0 U22123 ( .IN(n8247), .QN(n19150) );
  INVX0 U22124 ( .IN(n8249), .QN(n19117) );
  INVX0 U22125 ( .IN(n8243), .QN(n19216) );
  INVX0 U22126 ( .IN(n8541), .QN(n19051) );
  INVX0 U22127 ( .IN(n8543), .QN(n19018) );
  INVX0 U22128 ( .IN(n8545), .QN(n18985) );
  INVX0 U22129 ( .IN(n8539), .QN(n19084) );
  INVX0 U22130 ( .IN(n4509), .QN(n20852) );
  INVX0 U22131 ( .IN(n4511), .QN(n20834) );
  INVX0 U22132 ( .IN(n4513), .QN(n20816) );
  INVX0 U22133 ( .IN(n4507), .QN(n20870) );
  INVX0 U22134 ( .IN(n4510), .QN(n20843) );
  INVX0 U22135 ( .IN(n4512), .QN(n20825) );
  INVX0 U22136 ( .IN(n4805), .QN(n20765) );
  INVX0 U22137 ( .IN(n4807), .QN(n20732) );
  INVX0 U22138 ( .IN(n4809), .QN(n20699) );
  INVX0 U22139 ( .IN(n4803), .QN(n20798) );
  INVX0 U22140 ( .IN(n5101), .QN(n20633) );
  INVX0 U22141 ( .IN(n5103), .QN(n20600) );
  INVX0 U22142 ( .IN(n5105), .QN(n20567) );
  INVX0 U22143 ( .IN(n5099), .QN(n20666) );
  INVX0 U22144 ( .IN(n5397), .QN(n20501) );
  INVX0 U22145 ( .IN(n5399), .QN(n20468) );
  INVX0 U22146 ( .IN(n5401), .QN(n20435) );
  INVX0 U22147 ( .IN(n5395), .QN(n20534) );
  INVX0 U22148 ( .IN(n5693), .QN(n20369) );
  INVX0 U22149 ( .IN(n5695), .QN(n20336) );
  INVX0 U22150 ( .IN(n5697), .QN(n20303) );
  INVX0 U22151 ( .IN(n5691), .QN(n20402) );
  INVX0 U22152 ( .IN(n5989), .QN(n20237) );
  INVX0 U22153 ( .IN(n5991), .QN(n20204) );
  INVX0 U22154 ( .IN(n5993), .QN(n20171) );
  INVX0 U22155 ( .IN(n5987), .QN(n20270) );
  INVX0 U22156 ( .IN(n6285), .QN(n20105) );
  INVX0 U22157 ( .IN(n6287), .QN(n20073) );
  INVX0 U22158 ( .IN(n6289), .QN(n20040) );
  INVX0 U22159 ( .IN(n6283), .QN(n20138) );
  INVX0 U22160 ( .IN(n6581), .QN(n19974) );
  INVX0 U22161 ( .IN(n6583), .QN(n19942) );
  INVX0 U22162 ( .IN(n6585), .QN(n19909) );
  INVX0 U22163 ( .IN(n6579), .QN(n20007) );
  INVX0 U22164 ( .IN(n6877), .QN(n19843) );
  INVX0 U22165 ( .IN(n6879), .QN(n19810) );
  INVX0 U22166 ( .IN(n6881), .QN(n19777) );
  INVX0 U22167 ( .IN(n6875), .QN(n19876) );
  INVX0 U22168 ( .IN(n8837), .QN(n18919) );
  INVX0 U22169 ( .IN(n8839), .QN(n18886) );
  INVX0 U22170 ( .IN(n8841), .QN(n18853) );
  INVX0 U22171 ( .IN(n8835), .QN(n18952) );
  INVX0 U22172 ( .IN(n14523), .QN(n18793) );
  INVX0 U22173 ( .IN(n14533), .QN(n18769) );
  INVX0 U22174 ( .IN(n14900), .QN(n18757) );
  INVX0 U22175 ( .IN(n14905), .QN(n18745) );
  INVX0 U22176 ( .IN(n14910), .QN(n18733) );
  INVX0 U22177 ( .IN(n14915), .QN(n18721) );
  INVX0 U22178 ( .IN(n15210), .QN(n18697) );
  INVX0 U22179 ( .IN(n15220), .QN(n18673) );
  INVX0 U22180 ( .IN(n15510), .QN(n18661) );
  INVX0 U22181 ( .IN(n15515), .QN(n18649) );
  INVX0 U22182 ( .IN(n15520), .QN(n18637) );
  INVX0 U22183 ( .IN(n15525), .QN(n18625) );
  INVX0 U22184 ( .IN(n15820), .QN(n18601) );
  INVX0 U22185 ( .IN(n15830), .QN(n18577) );
  INVX0 U22186 ( .IN(n16120), .QN(n18565) );
  INVX0 U22187 ( .IN(n16125), .QN(n18553) );
  INVX0 U22188 ( .IN(n16130), .QN(n18541) );
  INVX0 U22189 ( .IN(n16135), .QN(n18529) );
  INVX0 U22190 ( .IN(n16430), .QN(n18505) );
  INVX0 U22191 ( .IN(n16440), .QN(n18481) );
  INVX0 U22192 ( .IN(n16730), .QN(n18469) );
  INVX0 U22193 ( .IN(n16735), .QN(n18457) );
  INVX0 U22194 ( .IN(n16740), .QN(n18445) );
  INVX0 U22195 ( .IN(n16745), .QN(n18433) );
  INVX0 U22196 ( .IN(n14912), .QN(n18727) );
  INVX0 U22197 ( .IN(n15522), .QN(n18631) );
  INVX0 U22198 ( .IN(n16132), .QN(n18535) );
  INVX0 U22199 ( .IN(n16742), .QN(n18439) );
  INVX0 U22200 ( .IN(n4508), .QN(n20861) );
  INVX0 U22201 ( .IN(n21086), .QN(n21081) );
  INVX0 U22202 ( .IN(n21086), .QN(n21082) );
  INVX0 U22203 ( .IN(n21087), .QN(n21080) );
  INVX0 U22204 ( .IN(n21085), .QN(n21083) );
  INVX0 U22205 ( .IN(n21084), .QN(n21068) );
  INVX0 U22206 ( .IN(n21085), .QN(n21084) );
  INVX0 U22207 ( .IN(n6286), .QN(n20074) );
  NBUFFX2 U22208 ( .IN(n21105), .Q(n18341) );
  NBUFFX2 U22209 ( .IN(n21104), .Q(n18343) );
  NBUFFX2 U22210 ( .IN(n21103), .Q(n18345) );
  NBUFFX2 U22211 ( .IN(n21102), .Q(n18347) );
  NBUFFX2 U22212 ( .IN(n21101), .Q(n18349) );
  NBUFFX2 U22213 ( .IN(n21100), .Q(n18351) );
  NBUFFX2 U22214 ( .IN(n21099), .Q(n18353) );
  NBUFFX2 U22215 ( .IN(n21098), .Q(n18355) );
  NBUFFX2 U22216 ( .IN(n21097), .Q(n18357) );
  NBUFFX2 U22217 ( .IN(n21096), .Q(n18359) );
  NBUFFX2 U22218 ( .IN(n21095), .Q(n18361) );
  NBUFFX2 U22219 ( .IN(n21094), .Q(n18363) );
  NBUFFX2 U22220 ( .IN(n21093), .Q(n18365) );
  NBUFFX2 U22221 ( .IN(n21092), .Q(n18367) );
  NBUFFX2 U22222 ( .IN(n21091), .Q(n18369) );
  NBUFFX2 U22223 ( .IN(n21090), .Q(n18339) );
  NBUFFX2 U22224 ( .IN(n21105), .Q(s15_data_o[0]) );
  NBUFFX2 U22225 ( .IN(n21104), .Q(s15_data_o[1]) );
  NBUFFX2 U22226 ( .IN(n21103), .Q(s15_data_o[2]) );
  NBUFFX2 U22227 ( .IN(n21102), .Q(s15_data_o[3]) );
  NBUFFX2 U22228 ( .IN(n21101), .Q(s15_data_o[4]) );
  NBUFFX2 U22229 ( .IN(n21100), .Q(s15_data_o[5]) );
  NBUFFX2 U22230 ( .IN(n21099), .Q(s15_data_o[6]) );
  NBUFFX2 U22231 ( .IN(n21098), .Q(s15_data_o[7]) );
  NBUFFX2 U22232 ( .IN(n21097), .Q(s15_data_o[8]) );
  NBUFFX2 U22233 ( .IN(n21096), .Q(s15_data_o[9]) );
  NBUFFX2 U22234 ( .IN(n21095), .Q(s15_data_o[10]) );
  NBUFFX2 U22235 ( .IN(n21094), .Q(s15_data_o[11]) );
  NBUFFX2 U22236 ( .IN(n21093), .Q(s15_data_o[12]) );
  NBUFFX2 U22237 ( .IN(n21092), .Q(s15_data_o[13]) );
  NBUFFX2 U22238 ( .IN(n21091), .Q(s15_data_o[14]) );
  NBUFFX2 U22239 ( .IN(n21090), .Q(s15_data_o[15]) );
  NBUFFX2 U22240 ( .IN(n12698), .Q(n18389) );
  NBUFFX2 U22241 ( .IN(n12698), .Q(n18388) );
  NBUFFX2 U22242 ( .IN(n12389), .Q(n18393) );
  NBUFFX2 U22243 ( .IN(n12389), .Q(n18392) );
  NBUFFX2 U22244 ( .IN(n12079), .Q(n18397) );
  NBUFFX2 U22245 ( .IN(n12079), .Q(n18396) );
  NBUFFX2 U22246 ( .IN(n11769), .Q(n18401) );
  NBUFFX2 U22247 ( .IN(n11769), .Q(n18400) );
  NOR2X0 U22248 ( .IN1(n13896), .IN2(n3224), .QN(n13887) );
  NOR2X0 U22249 ( .IN1(n13587), .IN2(n3228), .QN(n13578) );
  NOR2X0 U22250 ( .IN1(n11421), .IN2(n3196), .QN(n11412) );
  NOR2X0 U22251 ( .IN1(n13278), .IN2(n3232), .QN(n13269) );
  NOR2X0 U22252 ( .IN1(n12969), .IN2(n3236), .QN(n12960) );
  NOR2X0 U22253 ( .IN1(n11112), .IN2(n3200), .QN(n11103) );
  NOR2X0 U22254 ( .IN1(n10802), .IN2(n3204), .QN(n10793) );
  NOR2X0 U22255 ( .IN1(n12660), .IN2(n3240), .QN(n12651) );
  NOR2X0 U22256 ( .IN1(n12351), .IN2(n3244), .QN(n12342) );
  NOR2X0 U22257 ( .IN1(n10493), .IN2(n3208), .QN(n10484) );
  NOR2X0 U22258 ( .IN1(n10183), .IN2(n3212), .QN(n10174) );
  NOR2X0 U22259 ( .IN1(n12041), .IN2(n3248), .QN(n12032) );
  NOR2X0 U22260 ( .IN1(n11731), .IN2(n3252), .QN(n11722) );
  NOR2X0 U22261 ( .IN1(n9873), .IN2(n3216), .QN(n9864) );
  NOR2X0 U22262 ( .IN1(n9562), .IN2(n3220), .QN(n9553) );
  NOR2X0 U22263 ( .IN1(n14170), .IN2(n3190), .QN(n14161) );
  NOR2X0 U22264 ( .IN1(n3857), .IN2(n3854), .QN(n13744) );
  NOR2X0 U22265 ( .IN1(n3812), .IN2(n3809), .QN(n13435) );
  NOR2X0 U22266 ( .IN1(n4172), .IN2(n4169), .QN(n11269) );
  NOR2X0 U22267 ( .IN1(n3767), .IN2(n3764), .QN(n13126) );
  NOR2X0 U22268 ( .IN1(n3722), .IN2(n3719), .QN(n12817) );
  NOR2X0 U22269 ( .IN1(n4127), .IN2(n4124), .QN(n10960) );
  NOR2X0 U22270 ( .IN1(n4082), .IN2(n4079), .QN(n10650) );
  NOR2X0 U22271 ( .IN1(n3677), .IN2(n3674), .QN(n12508) );
  NOR2X0 U22272 ( .IN1(n3632), .IN2(n3629), .QN(n12199) );
  NOR2X0 U22273 ( .IN1(n4037), .IN2(n4034), .QN(n10341) );
  NOR2X0 U22274 ( .IN1(n3992), .IN2(n3989), .QN(n10031) );
  NOR2X0 U22275 ( .IN1(n3587), .IN2(n3584), .QN(n11889) );
  NOR2X0 U22276 ( .IN1(n3542), .IN2(n3539), .QN(n11579) );
  NOR2X0 U22277 ( .IN1(n3947), .IN2(n3944), .QN(n9721) );
  NOR2X0 U22278 ( .IN1(n3902), .IN2(n3899), .QN(n9410) );
  NOR2X0 U22279 ( .IN1(n4217), .IN2(n4214), .QN(n14008) );
  NOR2X0 U22280 ( .IN1(n3881), .IN2(n3878), .QN(n13875) );
  NOR2X0 U22281 ( .IN1(n3836), .IN2(n3833), .QN(n13566) );
  NOR2X0 U22282 ( .IN1(n4196), .IN2(n4193), .QN(n11400) );
  NOR2X0 U22283 ( .IN1(n3791), .IN2(n3788), .QN(n13257) );
  NOR2X0 U22284 ( .IN1(n3746), .IN2(n3743), .QN(n12948) );
  NOR2X0 U22285 ( .IN1(n4151), .IN2(n4148), .QN(n11091) );
  NOR2X0 U22286 ( .IN1(n4106), .IN2(n4103), .QN(n10781) );
  NOR2X0 U22287 ( .IN1(n3701), .IN2(n3698), .QN(n12639) );
  NOR2X0 U22288 ( .IN1(n3656), .IN2(n3653), .QN(n12330) );
  NOR2X0 U22289 ( .IN1(n4061), .IN2(n4058), .QN(n10472) );
  NOR2X0 U22290 ( .IN1(n4016), .IN2(n4013), .QN(n10162) );
  NOR2X0 U22291 ( .IN1(n3611), .IN2(n3608), .QN(n12020) );
  NOR2X0 U22292 ( .IN1(n3566), .IN2(n3563), .QN(n11710) );
  NOR2X0 U22293 ( .IN1(n3971), .IN2(n3968), .QN(n9852) );
  NOR2X0 U22294 ( .IN1(n3926), .IN2(n3923), .QN(n9541) );
  NOR2X0 U22295 ( .IN1(n4241), .IN2(n4238), .QN(n14149) );
  NOR2X0 U22296 ( .IN1(n3865), .IN2(n3862), .QN(n13809) );
  NOR2X0 U22297 ( .IN1(n3873), .IN2(n3870), .QN(n13684) );
  NOR2X0 U22298 ( .IN1(n3820), .IN2(n3817), .QN(n13500) );
  NOR2X0 U22299 ( .IN1(n3828), .IN2(n3825), .QN(n13375) );
  NOR2X0 U22300 ( .IN1(n4180), .IN2(n4177), .QN(n11334) );
  NOR2X0 U22301 ( .IN1(n4188), .IN2(n4185), .QN(n11209) );
  NOR2X0 U22302 ( .IN1(n3775), .IN2(n3772), .QN(n13191) );
  NOR2X0 U22303 ( .IN1(n3783), .IN2(n3780), .QN(n13066) );
  NOR2X0 U22304 ( .IN1(n3730), .IN2(n3727), .QN(n12882) );
  NOR2X0 U22305 ( .IN1(n3738), .IN2(n3735), .QN(n12757) );
  NOR2X0 U22306 ( .IN1(n4135), .IN2(n4132), .QN(n11025) );
  NOR2X0 U22307 ( .IN1(n4143), .IN2(n4140), .QN(n10900) );
  NOR2X0 U22308 ( .IN1(n4090), .IN2(n4087), .QN(n10715) );
  NOR2X0 U22309 ( .IN1(n4098), .IN2(n4095), .QN(n10590) );
  NOR2X0 U22310 ( .IN1(n3685), .IN2(n3682), .QN(n12573) );
  NOR2X0 U22311 ( .IN1(n3693), .IN2(n3690), .QN(n12448) );
  NOR2X0 U22312 ( .IN1(n3640), .IN2(n3637), .QN(n12264) );
  NOR2X0 U22313 ( .IN1(n3648), .IN2(n3645), .QN(n12139) );
  NOR2X0 U22314 ( .IN1(n4045), .IN2(n4042), .QN(n10406) );
  NOR2X0 U22315 ( .IN1(n4053), .IN2(n4050), .QN(n10281) );
  NOR2X0 U22316 ( .IN1(n4000), .IN2(n3997), .QN(n10096) );
  NOR2X0 U22317 ( .IN1(n4008), .IN2(n4005), .QN(n9971) );
  NOR2X0 U22318 ( .IN1(n3595), .IN2(n3592), .QN(n11954) );
  NOR2X0 U22319 ( .IN1(n3603), .IN2(n3600), .QN(n11829) );
  NOR2X0 U22320 ( .IN1(n3550), .IN2(n3547), .QN(n11644) );
  NOR2X0 U22321 ( .IN1(n3558), .IN2(n3555), .QN(n11519) );
  NOR2X0 U22322 ( .IN1(n3955), .IN2(n3952), .QN(n9786) );
  NOR2X0 U22323 ( .IN1(n3963), .IN2(n3960), .QN(n9661) );
  NOR2X0 U22324 ( .IN1(n3910), .IN2(n3907), .QN(n9475) );
  NOR2X0 U22325 ( .IN1(n3918), .IN2(n3915), .QN(n9350) );
  NOR2X0 U22326 ( .IN1(n4225), .IN2(n4222), .QN(n13940) );
  NOR2X0 U22327 ( .IN1(n4233), .IN2(n4230), .QN(n14081) );
  NAND2X0 U22328 ( .IN1(n2974), .IN2(n3144), .QN(n13828) );
  NAND2X0 U22329 ( .IN1(n2990), .IN2(n3150), .QN(n13519) );
  NAND2X0 U22330 ( .IN1(n2862), .IN2(n3102), .QN(n11353) );
  NAND2X0 U22331 ( .IN1(n3006), .IN2(n3156), .QN(n13210) );
  NAND2X0 U22332 ( .IN1(n3022), .IN2(n3162), .QN(n12901) );
  NAND2X0 U22333 ( .IN1(n2878), .IN2(n3108), .QN(n11044) );
  NAND2X0 U22334 ( .IN1(n2894), .IN2(n3114), .QN(n10734) );
  NAND2X0 U22335 ( .IN1(n3038), .IN2(n3168), .QN(n12592) );
  NAND2X0 U22336 ( .IN1(n3054), .IN2(n3174), .QN(n12283) );
  NAND2X0 U22337 ( .IN1(n2910), .IN2(n3120), .QN(n10425) );
  NAND2X0 U22338 ( .IN1(n2926), .IN2(n3126), .QN(n10115) );
  NAND2X0 U22339 ( .IN1(n3070), .IN2(n3180), .QN(n11973) );
  NAND2X0 U22340 ( .IN1(n3086), .IN2(n3186), .QN(n11663) );
  NAND2X0 U22341 ( .IN1(n2942), .IN2(n3132), .QN(n9805) );
  NAND2X0 U22342 ( .IN1(n2958), .IN2(n3138), .QN(n9494) );
  NAND2X0 U22343 ( .IN1(n2844), .IN2(n3095), .QN(n13961) );
  NAND2X0 U22344 ( .IN1(n2966), .IN2(n3141), .QN(n13702) );
  NAND2X0 U22345 ( .IN1(n2982), .IN2(n3147), .QN(n13393) );
  NAND2X0 U22346 ( .IN1(n2854), .IN2(n3099), .QN(n11227) );
  NAND2X0 U22347 ( .IN1(n2998), .IN2(n3153), .QN(n13084) );
  NAND2X0 U22348 ( .IN1(n3014), .IN2(n3159), .QN(n12775) );
  NAND2X0 U22349 ( .IN1(n2870), .IN2(n3105), .QN(n10918) );
  NAND2X0 U22350 ( .IN1(n2886), .IN2(n3111), .QN(n10608) );
  NAND2X0 U22351 ( .IN1(n3030), .IN2(n3165), .QN(n12466) );
  NAND2X0 U22352 ( .IN1(n3046), .IN2(n3171), .QN(n12157) );
  NAND2X0 U22353 ( .IN1(n2902), .IN2(n3117), .QN(n10299) );
  NAND2X0 U22354 ( .IN1(n2918), .IN2(n3123), .QN(n9989) );
  NAND2X0 U22355 ( .IN1(n3062), .IN2(n3177), .QN(n11847) );
  NAND2X0 U22356 ( .IN1(n3078), .IN2(n3183), .QN(n11537) );
  NAND2X0 U22357 ( .IN1(n2934), .IN2(n3129), .QN(n9679) );
  NAND2X0 U22358 ( .IN1(n2950), .IN2(n3135), .QN(n9368) );
  NAND2X0 U22359 ( .IN1(n2849), .IN2(n3097), .QN(n14101) );
  NAND2X0 U22360 ( .IN1(n2971), .IN2(n3143), .QN(n13765) );
  NAND2X0 U22361 ( .IN1(n2987), .IN2(n3149), .QN(n13456) );
  NAND2X0 U22362 ( .IN1(n2859), .IN2(n3101), .QN(n11290) );
  NAND2X0 U22363 ( .IN1(n3003), .IN2(n3155), .QN(n13147) );
  NAND2X0 U22364 ( .IN1(n3019), .IN2(n3161), .QN(n12838) );
  NAND2X0 U22365 ( .IN1(n2875), .IN2(n3107), .QN(n10981) );
  NAND2X0 U22366 ( .IN1(n2891), .IN2(n3113), .QN(n10671) );
  NAND2X0 U22367 ( .IN1(n3035), .IN2(n3167), .QN(n12529) );
  NAND2X0 U22368 ( .IN1(n3051), .IN2(n3173), .QN(n12220) );
  NAND2X0 U22369 ( .IN1(n2907), .IN2(n3119), .QN(n10362) );
  NAND2X0 U22370 ( .IN1(n2923), .IN2(n3125), .QN(n10052) );
  NAND2X0 U22371 ( .IN1(n3067), .IN2(n3179), .QN(n11910) );
  NAND2X0 U22372 ( .IN1(n3083), .IN2(n3185), .QN(n11600) );
  NAND2X0 U22373 ( .IN1(n2939), .IN2(n3131), .QN(n9742) );
  NAND2X0 U22374 ( .IN1(n2955), .IN2(n3137), .QN(n9431) );
  NAND2X0 U22375 ( .IN1(n2838), .IN2(n3093), .QN(n14029) );
  INVX0 U22376 ( .IN(n13819), .QN(n2976) );
  INVX0 U22377 ( .IN(n13693), .QN(n2968) );
  INVX0 U22378 ( .IN(n13510), .QN(n2992) );
  INVX0 U22379 ( .IN(n13384), .QN(n2984) );
  INVX0 U22380 ( .IN(n11344), .QN(n2864) );
  INVX0 U22381 ( .IN(n11218), .QN(n2856) );
  INVX0 U22382 ( .IN(n13201), .QN(n3008) );
  INVX0 U22383 ( .IN(n13075), .QN(n3000) );
  INVX0 U22384 ( .IN(n12892), .QN(n3024) );
  INVX0 U22385 ( .IN(n12766), .QN(n3016) );
  INVX0 U22386 ( .IN(n11035), .QN(n2880) );
  INVX0 U22387 ( .IN(n10909), .QN(n2872) );
  INVX0 U22388 ( .IN(n10725), .QN(n2896) );
  INVX0 U22389 ( .IN(n10599), .QN(n2888) );
  INVX0 U22390 ( .IN(n12583), .QN(n3040) );
  INVX0 U22391 ( .IN(n12457), .QN(n3032) );
  INVX0 U22392 ( .IN(n12274), .QN(n3056) );
  INVX0 U22393 ( .IN(n12148), .QN(n3048) );
  INVX0 U22394 ( .IN(n10416), .QN(n2912) );
  INVX0 U22395 ( .IN(n10290), .QN(n2904) );
  INVX0 U22396 ( .IN(n10106), .QN(n2928) );
  INVX0 U22397 ( .IN(n9980), .QN(n2920) );
  INVX0 U22398 ( .IN(n11964), .QN(n3072) );
  INVX0 U22399 ( .IN(n11838), .QN(n3064) );
  INVX0 U22400 ( .IN(n11654), .QN(n3088) );
  INVX0 U22401 ( .IN(n11528), .QN(n3080) );
  INVX0 U22402 ( .IN(n9796), .QN(n2944) );
  INVX0 U22403 ( .IN(n9670), .QN(n2936) );
  INVX0 U22404 ( .IN(n9485), .QN(n2960) );
  INVX0 U22405 ( .IN(n9359), .QN(n2952) );
  INVX0 U22406 ( .IN(n13951), .QN(n2846) );
  INVX0 U22407 ( .IN(n14091), .QN(n2851) );
  INVX0 U22408 ( .IN(n21068), .QN(n21079) );
  INVX0 U22409 ( .IN(n21021), .QN(n21078) );
  NAND2X0 U22410 ( .IN1(n17964), .IN2(n18152), .QN(n13666) );
  NAND2X0 U22411 ( .IN1(n18155), .IN2(n17947), .QN(n13357) );
  NAND2X0 U22412 ( .IN1(n18156), .IN2(n17948), .QN(n11191) );
  NAND2X0 U22413 ( .IN1(n18063), .IN2(n17935), .QN(n13048) );
  NAND2X0 U22414 ( .IN1(n17934), .IN2(n18066), .QN(n12739) );
  NAND2X0 U22415 ( .IN1(n18062), .IN2(n17936), .QN(n10882) );
  NAND2X0 U22416 ( .IN1(n17958), .IN2(n18083), .QN(n10572) );
  NAND2X0 U22417 ( .IN1(n17945), .IN2(n18151), .QN(n12430) );
  NAND2X0 U22418 ( .IN1(n18154), .IN2(n17946), .QN(n12121) );
  NAND2X0 U22419 ( .IN1(n18061), .IN2(n17937), .QN(n10263) );
  NAND2X0 U22420 ( .IN1(n17957), .IN2(n18084), .QN(n9953) );
  NAND2X0 U22421 ( .IN1(n18064), .IN2(n17938), .QN(n11811) );
  NAND2X0 U22422 ( .IN1(n17959), .IN2(n18085), .QN(n11501) );
  NAND2X0 U22423 ( .IN1(n18153), .IN2(n17940), .QN(n9643) );
  NAND2X0 U22424 ( .IN1(n17933), .IN2(n18065), .QN(n9332) );
  OA22X1 U22425 ( .IN1(n13471), .IN2(n13448), .IN3(n13473), .IN4(n13475), .Q(
        n13493) );
  OA22X1 U22426 ( .IN1(n10996), .IN2(n10973), .IN3(n10998), .IN4(n11000), .Q(
        n11018) );
  OA22X1 U22427 ( .IN1(n10377), .IN2(n10354), .IN3(n10379), .IN4(n10381), .Q(
        n10399) );
  OA22X1 U22428 ( .IN1(n9757), .IN2(n9734), .IN3(n9759), .IN4(n9761), .Q(n9779) );
  AND2X1 U22429 ( .IN1(n13471), .IN2(n13475), .Q(n13439) );
  AND2X1 U22430 ( .IN1(n10996), .IN2(n11000), .Q(n10964) );
  AND2X1 U22431 ( .IN1(n10377), .IN2(n10381), .Q(n10345) );
  AND2X1 U22432 ( .IN1(n9757), .IN2(n9761), .Q(n9725) );
  AND2X1 U22433 ( .IN1(n11305), .IN2(n11309), .Q(n11273) );
  AND2X1 U22434 ( .IN1(n10686), .IN2(n10690), .Q(n10654) );
  AND2X1 U22435 ( .IN1(n10067), .IN2(n10071), .Q(n10035) );
  AND2X1 U22436 ( .IN1(n9446), .IN2(n9450), .Q(n9414) );
  OA22X1 U22437 ( .IN1(n3149), .IN2(n13465), .IN3(n13464), .IN4(n2987), .Q(
        n13491) );
  OA22X1 U22438 ( .IN1(n13443), .IN2(n3328), .IN3(n13462), .IN4(n3226), .Q(
        n13492) );
  OA22X1 U22439 ( .IN1(n3499), .IN2(n13490), .IN3(n13449), .IN4(n3435), .Q(
        n13494) );
  OA22X1 U22440 ( .IN1(n3107), .IN2(n10990), .IN3(n10989), .IN4(n2875), .Q(
        n11016) );
  OA22X1 U22441 ( .IN1(n10968), .IN2(n3272), .IN3(n10987), .IN4(n3198), .Q(
        n11017) );
  OA22X1 U22442 ( .IN1(n3471), .IN2(n11015), .IN3(n10974), .IN4(n3407), .Q(
        n11019) );
  OA22X1 U22443 ( .IN1(n3119), .IN2(n10371), .IN3(n10370), .IN4(n2907), .Q(
        n10397) );
  OA22X1 U22444 ( .IN1(n10349), .IN2(n3288), .IN3(n10368), .IN4(n3206), .Q(
        n10398) );
  OA22X1 U22445 ( .IN1(n3479), .IN2(n10396), .IN3(n10355), .IN4(n3415), .Q(
        n10400) );
  OA22X1 U22446 ( .IN1(n3131), .IN2(n9751), .IN3(n9750), .IN4(n2939), .Q(n9777) );
  OA22X1 U22447 ( .IN1(n9729), .IN2(n3304), .IN3(n9748), .IN4(n3214), .Q(n9778) );
  OA22X1 U22448 ( .IN1(n3487), .IN2(n9776), .IN3(n9735), .IN4(n3423), .Q(n9780) );
  OA22X1 U22449 ( .IN1(n3143), .IN2(n13774), .IN3(n13773), .IN4(n2971), .Q(
        n13800) );
  OA22X1 U22450 ( .IN1(n13752), .IN2(n3320), .IN3(n13771), .IN4(n3222), .Q(
        n13801) );
  OA22X1 U22451 ( .IN1(n3495), .IN2(n13799), .IN3(n13758), .IN4(n3431), .Q(
        n13803) );
  OA22X1 U22452 ( .IN1(n3101), .IN2(n11299), .IN3(n11298), .IN4(n2859), .Q(
        n11325) );
  OA22X1 U22453 ( .IN1(n11277), .IN2(n3264), .IN3(n11296), .IN4(n3194), .Q(
        n11326) );
  OA22X1 U22454 ( .IN1(n3467), .IN2(n11324), .IN3(n11283), .IN4(n3403), .Q(
        n11328) );
  OA22X1 U22455 ( .IN1(n3155), .IN2(n13156), .IN3(n13155), .IN4(n3003), .Q(
        n13182) );
  OA22X1 U22456 ( .IN1(n13134), .IN2(n3336), .IN3(n13153), .IN4(n3230), .Q(
        n13183) );
  OA22X1 U22457 ( .IN1(n3503), .IN2(n13181), .IN3(n13140), .IN4(n3439), .Q(
        n13185) );
  OA22X1 U22458 ( .IN1(n3161), .IN2(n12847), .IN3(n12846), .IN4(n3019), .Q(
        n12873) );
  OA22X1 U22459 ( .IN1(n12825), .IN2(n3344), .IN3(n12844), .IN4(n3234), .Q(
        n12874) );
  OA22X1 U22460 ( .IN1(n3507), .IN2(n12872), .IN3(n12831), .IN4(n3443), .Q(
        n12876) );
  OA22X1 U22461 ( .IN1(n3113), .IN2(n10680), .IN3(n10679), .IN4(n2891), .Q(
        n10706) );
  OA22X1 U22462 ( .IN1(n10658), .IN2(n3280), .IN3(n10677), .IN4(n3202), .Q(
        n10707) );
  OA22X1 U22463 ( .IN1(n3475), .IN2(n10705), .IN3(n10664), .IN4(n3411), .Q(
        n10709) );
  OA22X1 U22464 ( .IN1(n3167), .IN2(n12538), .IN3(n12537), .IN4(n3035), .Q(
        n12564) );
  OA22X1 U22465 ( .IN1(n12516), .IN2(n3352), .IN3(n12535), .IN4(n3238), .Q(
        n12565) );
  OA22X1 U22466 ( .IN1(n3511), .IN2(n12563), .IN3(n12522), .IN4(n3447), .Q(
        n12567) );
  OA22X1 U22467 ( .IN1(n3173), .IN2(n12229), .IN3(n12228), .IN4(n3051), .Q(
        n12255) );
  OA22X1 U22468 ( .IN1(n12207), .IN2(n3360), .IN3(n12226), .IN4(n3242), .Q(
        n12256) );
  OA22X1 U22469 ( .IN1(n3515), .IN2(n12254), .IN3(n12213), .IN4(n3451), .Q(
        n12258) );
  OA22X1 U22470 ( .IN1(n3125), .IN2(n10061), .IN3(n10060), .IN4(n2923), .Q(
        n10087) );
  OA22X1 U22471 ( .IN1(n10039), .IN2(n3296), .IN3(n10058), .IN4(n3210), .Q(
        n10088) );
  OA22X1 U22472 ( .IN1(n3483), .IN2(n10086), .IN3(n10045), .IN4(n3419), .Q(
        n10090) );
  OA22X1 U22473 ( .IN1(n3179), .IN2(n11919), .IN3(n11918), .IN4(n3067), .Q(
        n11945) );
  OA22X1 U22474 ( .IN1(n11897), .IN2(n3368), .IN3(n11916), .IN4(n3246), .Q(
        n11946) );
  OA22X1 U22475 ( .IN1(n3519), .IN2(n11944), .IN3(n11903), .IN4(n3455), .Q(
        n11948) );
  OA22X1 U22476 ( .IN1(n3185), .IN2(n11609), .IN3(n11608), .IN4(n3083), .Q(
        n11635) );
  OA22X1 U22477 ( .IN1(n11587), .IN2(n3376), .IN3(n11606), .IN4(n3250), .Q(
        n11636) );
  OA22X1 U22478 ( .IN1(n3523), .IN2(n11634), .IN3(n11593), .IN4(n3459), .Q(
        n11638) );
  OA22X1 U22479 ( .IN1(n3137), .IN2(n9440), .IN3(n9439), .IN4(n2955), .Q(n9466) );
  OA22X1 U22480 ( .IN1(n9418), .IN2(n3312), .IN3(n9437), .IN4(n3218), .Q(n9467) );
  OA22X1 U22481 ( .IN1(n3491), .IN2(n9465), .IN3(n9424), .IN4(n3427), .Q(n9469) );
  AO221X1 U22482 ( .IN1(n13856), .IN2(n13857), .IN3(n13854), .IN4(n3866), 
        .IN5(n13858), .Q(n13821) );
  NOR2X0 U22483 ( .IN1(n13835), .IN2(n13832), .QN(n13856) );
  AO22X1 U22484 ( .IN1(n3864), .IN2(n13857), .IN3(n3863), .IN4(n13859), .Q(
        n13858) );
  INVX0 U22485 ( .IN(n13834), .QN(n3864) );
  AO221X1 U22486 ( .IN1(n13725), .IN2(n13726), .IN3(n13678), .IN4(n3874), 
        .IN5(n13727), .Q(n13695) );
  NOR2X0 U22487 ( .IN1(n13675), .IN2(n13673), .QN(n13725) );
  AO22X1 U22488 ( .IN1(n3872), .IN2(n13726), .IN3(n3871), .IN4(n13728), .Q(
        n13727) );
  INVX0 U22489 ( .IN(n13707), .QN(n3872) );
  AO221X1 U22490 ( .IN1(n13547), .IN2(n13548), .IN3(n13545), .IN4(n3821), 
        .IN5(n13549), .Q(n13512) );
  NOR2X0 U22491 ( .IN1(n13526), .IN2(n13523), .QN(n13547) );
  AO22X1 U22492 ( .IN1(n3819), .IN2(n13548), .IN3(n3818), .IN4(n13550), .Q(
        n13549) );
  INVX0 U22493 ( .IN(n13525), .QN(n3819) );
  AO221X1 U22494 ( .IN1(n13416), .IN2(n13417), .IN3(n13369), .IN4(n3829), 
        .IN5(n13418), .Q(n13386) );
  NOR2X0 U22495 ( .IN1(n13366), .IN2(n13364), .QN(n13416) );
  AO22X1 U22496 ( .IN1(n3827), .IN2(n13417), .IN3(n3826), .IN4(n13419), .Q(
        n13418) );
  INVX0 U22497 ( .IN(n13398), .QN(n3827) );
  AO221X1 U22498 ( .IN1(n11381), .IN2(n11382), .IN3(n11379), .IN4(n4181), 
        .IN5(n11383), .Q(n11346) );
  NOR2X0 U22499 ( .IN1(n11360), .IN2(n11357), .QN(n11381) );
  AO22X1 U22500 ( .IN1(n4179), .IN2(n11382), .IN3(n4178), .IN4(n11384), .Q(
        n11383) );
  INVX0 U22501 ( .IN(n11359), .QN(n4179) );
  AO221X1 U22502 ( .IN1(n11250), .IN2(n11251), .IN3(n11203), .IN4(n4189), 
        .IN5(n11252), .Q(n11220) );
  NOR2X0 U22503 ( .IN1(n11200), .IN2(n11198), .QN(n11250) );
  AO22X1 U22504 ( .IN1(n4187), .IN2(n11251), .IN3(n4186), .IN4(n11253), .Q(
        n11252) );
  INVX0 U22505 ( .IN(n11232), .QN(n4187) );
  AO221X1 U22506 ( .IN1(n13238), .IN2(n13239), .IN3(n13236), .IN4(n3776), 
        .IN5(n13240), .Q(n13203) );
  NOR2X0 U22507 ( .IN1(n13217), .IN2(n13214), .QN(n13238) );
  AO22X1 U22508 ( .IN1(n3774), .IN2(n13239), .IN3(n3773), .IN4(n13241), .Q(
        n13240) );
  INVX0 U22509 ( .IN(n13216), .QN(n3774) );
  AO221X1 U22510 ( .IN1(n13107), .IN2(n13108), .IN3(n13060), .IN4(n3784), 
        .IN5(n13109), .Q(n13077) );
  NOR2X0 U22511 ( .IN1(n13057), .IN2(n13055), .QN(n13107) );
  AO22X1 U22512 ( .IN1(n3782), .IN2(n13108), .IN3(n3781), .IN4(n13110), .Q(
        n13109) );
  INVX0 U22513 ( .IN(n13089), .QN(n3782) );
  AO221X1 U22514 ( .IN1(n12929), .IN2(n12930), .IN3(n12927), .IN4(n3731), 
        .IN5(n12931), .Q(n12894) );
  NOR2X0 U22515 ( .IN1(n12908), .IN2(n12905), .QN(n12929) );
  AO22X1 U22516 ( .IN1(n3729), .IN2(n12930), .IN3(n3728), .IN4(n12932), .Q(
        n12931) );
  INVX0 U22517 ( .IN(n12907), .QN(n3729) );
  AO221X1 U22518 ( .IN1(n12798), .IN2(n12799), .IN3(n12751), .IN4(n3739), 
        .IN5(n12800), .Q(n12768) );
  NOR2X0 U22519 ( .IN1(n12748), .IN2(n12746), .QN(n12798) );
  AO22X1 U22520 ( .IN1(n3737), .IN2(n12799), .IN3(n3736), .IN4(n12801), .Q(
        n12800) );
  INVX0 U22521 ( .IN(n12780), .QN(n3737) );
  AO221X1 U22522 ( .IN1(n11072), .IN2(n11073), .IN3(n11070), .IN4(n4136), 
        .IN5(n11074), .Q(n11037) );
  NOR2X0 U22523 ( .IN1(n11051), .IN2(n11048), .QN(n11072) );
  AO22X1 U22524 ( .IN1(n4134), .IN2(n11073), .IN3(n4133), .IN4(n11075), .Q(
        n11074) );
  INVX0 U22525 ( .IN(n11050), .QN(n4134) );
  AO221X1 U22526 ( .IN1(n10941), .IN2(n10942), .IN3(n10894), .IN4(n4144), 
        .IN5(n10943), .Q(n10911) );
  NOR2X0 U22527 ( .IN1(n10891), .IN2(n10889), .QN(n10941) );
  AO22X1 U22528 ( .IN1(n4142), .IN2(n10942), .IN3(n4141), .IN4(n10944), .Q(
        n10943) );
  INVX0 U22529 ( .IN(n10923), .QN(n4142) );
  AO221X1 U22530 ( .IN1(n10762), .IN2(n10763), .IN3(n10760), .IN4(n4091), 
        .IN5(n10764), .Q(n10727) );
  NOR2X0 U22531 ( .IN1(n10741), .IN2(n10738), .QN(n10762) );
  AO22X1 U22532 ( .IN1(n4089), .IN2(n10763), .IN3(n4088), .IN4(n10765), .Q(
        n10764) );
  INVX0 U22533 ( .IN(n10740), .QN(n4089) );
  AO221X1 U22534 ( .IN1(n10631), .IN2(n10632), .IN3(n10584), .IN4(n4099), 
        .IN5(n10633), .Q(n10601) );
  NOR2X0 U22535 ( .IN1(n10581), .IN2(n10579), .QN(n10631) );
  AO22X1 U22536 ( .IN1(n4097), .IN2(n10632), .IN3(n4096), .IN4(n10634), .Q(
        n10633) );
  INVX0 U22537 ( .IN(n10613), .QN(n4097) );
  AO221X1 U22538 ( .IN1(n12620), .IN2(n12621), .IN3(n12618), .IN4(n3686), 
        .IN5(n12622), .Q(n12585) );
  NOR2X0 U22539 ( .IN1(n12599), .IN2(n12596), .QN(n12620) );
  AO22X1 U22540 ( .IN1(n3684), .IN2(n12621), .IN3(n3683), .IN4(n12623), .Q(
        n12622) );
  INVX0 U22541 ( .IN(n12598), .QN(n3684) );
  AO221X1 U22542 ( .IN1(n12489), .IN2(n12490), .IN3(n12442), .IN4(n3694), 
        .IN5(n12491), .Q(n12459) );
  NOR2X0 U22543 ( .IN1(n12439), .IN2(n12437), .QN(n12489) );
  AO22X1 U22544 ( .IN1(n3692), .IN2(n12490), .IN3(n3691), .IN4(n12492), .Q(
        n12491) );
  INVX0 U22545 ( .IN(n12471), .QN(n3692) );
  AO221X1 U22546 ( .IN1(n12311), .IN2(n12312), .IN3(n12309), .IN4(n3641), 
        .IN5(n12313), .Q(n12276) );
  NOR2X0 U22547 ( .IN1(n12290), .IN2(n12287), .QN(n12311) );
  AO22X1 U22548 ( .IN1(n3639), .IN2(n12312), .IN3(n3638), .IN4(n12314), .Q(
        n12313) );
  INVX0 U22549 ( .IN(n12289), .QN(n3639) );
  AO221X1 U22550 ( .IN1(n12180), .IN2(n12181), .IN3(n12133), .IN4(n3649), 
        .IN5(n12182), .Q(n12150) );
  NOR2X0 U22551 ( .IN1(n12130), .IN2(n12128), .QN(n12180) );
  AO22X1 U22552 ( .IN1(n3647), .IN2(n12181), .IN3(n3646), .IN4(n12183), .Q(
        n12182) );
  INVX0 U22553 ( .IN(n12162), .QN(n3647) );
  AO221X1 U22554 ( .IN1(n10453), .IN2(n10454), .IN3(n10451), .IN4(n4046), 
        .IN5(n10455), .Q(n10418) );
  NOR2X0 U22555 ( .IN1(n10432), .IN2(n10429), .QN(n10453) );
  AO22X1 U22556 ( .IN1(n4044), .IN2(n10454), .IN3(n4043), .IN4(n10456), .Q(
        n10455) );
  INVX0 U22557 ( .IN(n10431), .QN(n4044) );
  AO221X1 U22558 ( .IN1(n10322), .IN2(n10323), .IN3(n10275), .IN4(n4054), 
        .IN5(n10324), .Q(n10292) );
  NOR2X0 U22559 ( .IN1(n10272), .IN2(n10270), .QN(n10322) );
  AO22X1 U22560 ( .IN1(n4052), .IN2(n10323), .IN3(n4051), .IN4(n10325), .Q(
        n10324) );
  INVX0 U22561 ( .IN(n10304), .QN(n4052) );
  AO221X1 U22562 ( .IN1(n10143), .IN2(n10144), .IN3(n10141), .IN4(n4001), 
        .IN5(n10145), .Q(n10108) );
  NOR2X0 U22563 ( .IN1(n10122), .IN2(n10119), .QN(n10143) );
  AO22X1 U22564 ( .IN1(n3999), .IN2(n10144), .IN3(n3998), .IN4(n10146), .Q(
        n10145) );
  INVX0 U22565 ( .IN(n10121), .QN(n3999) );
  AO221X1 U22566 ( .IN1(n10012), .IN2(n10013), .IN3(n9965), .IN4(n4009), .IN5(
        n10014), .Q(n9982) );
  NOR2X0 U22567 ( .IN1(n9962), .IN2(n9960), .QN(n10012) );
  AO22X1 U22568 ( .IN1(n4007), .IN2(n10013), .IN3(n4006), .IN4(n10015), .Q(
        n10014) );
  INVX0 U22569 ( .IN(n9994), .QN(n4007) );
  AO221X1 U22570 ( .IN1(n12001), .IN2(n12002), .IN3(n11999), .IN4(n3596), 
        .IN5(n12003), .Q(n11966) );
  NOR2X0 U22571 ( .IN1(n11980), .IN2(n11977), .QN(n12001) );
  AO22X1 U22572 ( .IN1(n3594), .IN2(n12002), .IN3(n3593), .IN4(n12004), .Q(
        n12003) );
  INVX0 U22573 ( .IN(n11979), .QN(n3594) );
  AO221X1 U22574 ( .IN1(n11870), .IN2(n11871), .IN3(n11823), .IN4(n3604), 
        .IN5(n11872), .Q(n11840) );
  NOR2X0 U22575 ( .IN1(n11820), .IN2(n11818), .QN(n11870) );
  AO22X1 U22576 ( .IN1(n3602), .IN2(n11871), .IN3(n3601), .IN4(n11873), .Q(
        n11872) );
  INVX0 U22577 ( .IN(n11852), .QN(n3602) );
  AO221X1 U22578 ( .IN1(n11691), .IN2(n11692), .IN3(n11689), .IN4(n3551), 
        .IN5(n11693), .Q(n11656) );
  NOR2X0 U22579 ( .IN1(n11670), .IN2(n11667), .QN(n11691) );
  AO22X1 U22580 ( .IN1(n3549), .IN2(n11692), .IN3(n3548), .IN4(n11694), .Q(
        n11693) );
  INVX0 U22581 ( .IN(n11669), .QN(n3549) );
  AO221X1 U22582 ( .IN1(n11560), .IN2(n11561), .IN3(n11513), .IN4(n3559), 
        .IN5(n11562), .Q(n11530) );
  NOR2X0 U22583 ( .IN1(n11510), .IN2(n11508), .QN(n11560) );
  AO22X1 U22584 ( .IN1(n3557), .IN2(n11561), .IN3(n3556), .IN4(n11563), .Q(
        n11562) );
  INVX0 U22585 ( .IN(n11542), .QN(n3557) );
  AO221X1 U22586 ( .IN1(n9833), .IN2(n9834), .IN3(n9831), .IN4(n3956), .IN5(
        n9835), .Q(n9798) );
  NOR2X0 U22587 ( .IN1(n9812), .IN2(n9809), .QN(n9833) );
  AO22X1 U22588 ( .IN1(n3954), .IN2(n9834), .IN3(n3953), .IN4(n9836), .Q(n9835) );
  INVX0 U22589 ( .IN(n9811), .QN(n3954) );
  AO221X1 U22590 ( .IN1(n9702), .IN2(n9703), .IN3(n9655), .IN4(n3964), .IN5(
        n9704), .Q(n9672) );
  NOR2X0 U22591 ( .IN1(n9652), .IN2(n9650), .QN(n9702) );
  AO22X1 U22592 ( .IN1(n3962), .IN2(n9703), .IN3(n3961), .IN4(n9705), .Q(n9704) );
  INVX0 U22593 ( .IN(n9684), .QN(n3962) );
  AO221X1 U22594 ( .IN1(n9522), .IN2(n9523), .IN3(n9520), .IN4(n3911), .IN5(
        n9524), .Q(n9487) );
  NOR2X0 U22595 ( .IN1(n9501), .IN2(n9498), .QN(n9522) );
  AO22X1 U22596 ( .IN1(n3909), .IN2(n9523), .IN3(n3908), .IN4(n9525), .Q(n9524) );
  INVX0 U22597 ( .IN(n9500), .QN(n3909) );
  AO221X1 U22598 ( .IN1(n9391), .IN2(n9392), .IN3(n9344), .IN4(n3919), .IN5(
        n9393), .Q(n9361) );
  NOR2X0 U22599 ( .IN1(n9341), .IN2(n9339), .QN(n9391) );
  AO22X1 U22600 ( .IN1(n3917), .IN2(n9392), .IN3(n3916), .IN4(n9394), .Q(n9393) );
  INVX0 U22601 ( .IN(n9373), .QN(n3917) );
  AND4X1 U22602 ( .IN1(n13854), .IN2(n3432), .IN3(n18163), .IN4(n13634), .Q(
        n13859) );
  AND4X1 U22603 ( .IN1(n13678), .IN2(n3430), .IN3(n18164), .IN4(n13670), .Q(
        n13728) );
  AND4X1 U22604 ( .IN1(n13545), .IN2(n3436), .IN3(n18159), .IN4(n13325), .Q(
        n13550) );
  AND4X1 U22605 ( .IN1(n13369), .IN2(n3434), .IN3(n18165), .IN4(n13361), .Q(
        n13419) );
  AND4X1 U22606 ( .IN1(n11379), .IN2(n3404), .IN3(n18160), .IN4(n11159), .Q(
        n11384) );
  AND4X1 U22607 ( .IN1(n11203), .IN2(n3402), .IN3(n18166), .IN4(n11195), .Q(
        n11253) );
  AND4X1 U22608 ( .IN1(n13236), .IN2(n3440), .IN3(n18167), .IN4(n13016), .Q(
        n13241) );
  AND4X1 U22609 ( .IN1(n13060), .IN2(n3438), .IN3(n18168), .IN4(n13052), .Q(
        n13110) );
  AND4X1 U22610 ( .IN1(n12927), .IN2(n3444), .IN3(n18169), .IN4(n12707), .Q(
        n12932) );
  AND4X1 U22611 ( .IN1(n12751), .IN2(n3442), .IN3(n18170), .IN4(n12743), .Q(
        n12801) );
  AND4X1 U22612 ( .IN1(n11070), .IN2(n3408), .IN3(n18171), .IN4(n10850), .Q(
        n11075) );
  AND4X1 U22613 ( .IN1(n10894), .IN2(n3406), .IN3(n18172), .IN4(n10886), .Q(
        n10944) );
  AND4X1 U22614 ( .IN1(n10760), .IN2(n3412), .IN3(n18173), .IN4(n10540), .Q(
        n10765) );
  AND4X1 U22615 ( .IN1(n10584), .IN2(n3410), .IN3(n18174), .IN4(n10576), .Q(
        n10634) );
  AND4X1 U22616 ( .IN1(n12618), .IN2(n3448), .IN3(n18175), .IN4(n12398), .Q(
        n12623) );
  AND4X1 U22617 ( .IN1(n12442), .IN2(n3446), .IN3(n18176), .IN4(n12434), .Q(
        n12492) );
  AND4X1 U22618 ( .IN1(n12309), .IN2(n3452), .IN3(n18161), .IN4(n12089), .Q(
        n12314) );
  AND4X1 U22619 ( .IN1(n12133), .IN2(n3450), .IN3(n18177), .IN4(n12125), .Q(
        n12183) );
  AND4X1 U22620 ( .IN1(n10451), .IN2(n3416), .IN3(n18178), .IN4(n10231), .Q(
        n10456) );
  AND4X1 U22621 ( .IN1(n10275), .IN2(n3414), .IN3(n18179), .IN4(n10267), .Q(
        n10325) );
  AND4X1 U22622 ( .IN1(n10141), .IN2(n3420), .IN3(n18180), .IN4(n9921), .Q(
        n10146) );
  AND4X1 U22623 ( .IN1(n9965), .IN2(n3418), .IN3(n18181), .IN4(n9957), .Q(
        n10015) );
  AND4X1 U22624 ( .IN1(n11999), .IN2(n3456), .IN3(n18182), .IN4(n11779), .Q(
        n12004) );
  AND4X1 U22625 ( .IN1(n11823), .IN2(n3454), .IN3(n18183), .IN4(n11815), .Q(
        n11873) );
  AND4X1 U22626 ( .IN1(n11689), .IN2(n3460), .IN3(n18184), .IN4(n11469), .Q(
        n11694) );
  AND4X1 U22627 ( .IN1(n11513), .IN2(n3458), .IN3(n18185), .IN4(n11505), .Q(
        n11563) );
  AND4X1 U22628 ( .IN1(n9831), .IN2(n3424), .IN3(n18162), .IN4(n9611), .Q(
        n9836) );
  AND4X1 U22629 ( .IN1(n9655), .IN2(n3422), .IN3(n18186), .IN4(n9647), .Q(
        n9705) );
  AND4X1 U22630 ( .IN1(n9520), .IN2(n3428), .IN3(n18187), .IN4(n9300), .Q(
        n9525) );
  AND4X1 U22631 ( .IN1(n9344), .IN2(n3426), .IN3(n18188), .IN4(n9336), .Q(
        n9394) );
  NAND3X0 U22632 ( .IN1(n13634), .IN2(n3322), .IN3(n18163), .QN(n13830) );
  NAND3X0 U22633 ( .IN1(n13670), .IN2(n3318), .IN3(n18164), .QN(n13704) );
  NAND3X0 U22634 ( .IN1(n13325), .IN2(n3330), .IN3(n18159), .QN(n13521) );
  NAND3X0 U22635 ( .IN1(n13361), .IN2(n3326), .IN3(n18165), .QN(n13395) );
  NAND3X0 U22636 ( .IN1(n11159), .IN2(n3266), .IN3(n18160), .QN(n11355) );
  NAND3X0 U22637 ( .IN1(n11195), .IN2(n3262), .IN3(n18166), .QN(n11229) );
  NAND3X0 U22638 ( .IN1(n13016), .IN2(n3338), .IN3(n18167), .QN(n13212) );
  NAND3X0 U22639 ( .IN1(n13052), .IN2(n3334), .IN3(n18168), .QN(n13086) );
  NAND3X0 U22640 ( .IN1(n12707), .IN2(n3346), .IN3(n18169), .QN(n12903) );
  NAND3X0 U22641 ( .IN1(n12743), .IN2(n3342), .IN3(n18170), .QN(n12777) );
  NAND3X0 U22642 ( .IN1(n10850), .IN2(n3274), .IN3(n18171), .QN(n11046) );
  NAND3X0 U22643 ( .IN1(n10886), .IN2(n3270), .IN3(n18172), .QN(n10920) );
  NAND3X0 U22644 ( .IN1(n10540), .IN2(n3282), .IN3(n18173), .QN(n10736) );
  NAND3X0 U22645 ( .IN1(n10576), .IN2(n3278), .IN3(n18174), .QN(n10610) );
  NAND3X0 U22646 ( .IN1(n12398), .IN2(n3354), .IN3(n18175), .QN(n12594) );
  NAND3X0 U22647 ( .IN1(n12434), .IN2(n3350), .IN3(n18176), .QN(n12468) );
  NAND3X0 U22648 ( .IN1(n12089), .IN2(n3362), .IN3(n18161), .QN(n12285) );
  NAND3X0 U22649 ( .IN1(n12125), .IN2(n3358), .IN3(n18177), .QN(n12159) );
  NAND3X0 U22650 ( .IN1(n10231), .IN2(n3290), .IN3(n18178), .QN(n10427) );
  NAND3X0 U22651 ( .IN1(n10267), .IN2(n3286), .IN3(n18179), .QN(n10301) );
  NAND3X0 U22652 ( .IN1(n9921), .IN2(n3298), .IN3(n18180), .QN(n10117) );
  NAND3X0 U22653 ( .IN1(n9957), .IN2(n3294), .IN3(n18181), .QN(n9991) );
  NAND3X0 U22654 ( .IN1(n11779), .IN2(n3370), .IN3(n18182), .QN(n11975) );
  NAND3X0 U22655 ( .IN1(n11815), .IN2(n3366), .IN3(n18183), .QN(n11849) );
  NAND3X0 U22656 ( .IN1(n11469), .IN2(n3378), .IN3(n18184), .QN(n11665) );
  NAND3X0 U22657 ( .IN1(n11505), .IN2(n3374), .IN3(n18185), .QN(n11539) );
  NAND3X0 U22658 ( .IN1(n9611), .IN2(n3306), .IN3(n18162), .QN(n9807) );
  NAND3X0 U22659 ( .IN1(n9647), .IN2(n3302), .IN3(n18186), .QN(n9681) );
  NAND3X0 U22660 ( .IN1(n9300), .IN2(n3314), .IN3(n18187), .QN(n9496) );
  NAND3X0 U22661 ( .IN1(n9336), .IN2(n3310), .IN3(n18188), .QN(n9370) );
  AO221X1 U22662 ( .IN1(n3855), .IN2(n13793), .IN3(n3856), .IN4(n13794), .IN5(
        n13795), .Q(n13747) );
  INVX0 U22663 ( .IN(n13771), .QN(n3856) );
  AO22X1 U22664 ( .IN1(n13791), .IN2(n3858), .IN3(n13796), .IN4(n13794), .Q(
        n13795) );
  NOR2X0 U22665 ( .IN1(n13772), .IN2(n13769), .QN(n13796) );
  AO221X1 U22666 ( .IN1(n3810), .IN2(n13484), .IN3(n3811), .IN4(n13485), .IN5(
        n13486), .Q(n13438) );
  INVX0 U22667 ( .IN(n13462), .QN(n3811) );
  AO22X1 U22668 ( .IN1(n13482), .IN2(n3813), .IN3(n13487), .IN4(n13485), .Q(
        n13486) );
  NOR2X0 U22669 ( .IN1(n13463), .IN2(n13460), .QN(n13487) );
  AO221X1 U22670 ( .IN1(n4170), .IN2(n11318), .IN3(n4171), .IN4(n11319), .IN5(
        n11320), .Q(n11272) );
  INVX0 U22671 ( .IN(n11296), .QN(n4171) );
  AO22X1 U22672 ( .IN1(n11316), .IN2(n4173), .IN3(n11321), .IN4(n11319), .Q(
        n11320) );
  NOR2X0 U22673 ( .IN1(n11297), .IN2(n11294), .QN(n11321) );
  AO221X1 U22674 ( .IN1(n3765), .IN2(n13175), .IN3(n3766), .IN4(n13176), .IN5(
        n13177), .Q(n13129) );
  INVX0 U22675 ( .IN(n13153), .QN(n3766) );
  AO22X1 U22676 ( .IN1(n13173), .IN2(n3768), .IN3(n13178), .IN4(n13176), .Q(
        n13177) );
  NOR2X0 U22677 ( .IN1(n13154), .IN2(n13151), .QN(n13178) );
  AO221X1 U22678 ( .IN1(n3720), .IN2(n12866), .IN3(n3721), .IN4(n12867), .IN5(
        n12868), .Q(n12820) );
  INVX0 U22679 ( .IN(n12844), .QN(n3721) );
  AO22X1 U22680 ( .IN1(n12864), .IN2(n3723), .IN3(n12869), .IN4(n12867), .Q(
        n12868) );
  NOR2X0 U22681 ( .IN1(n12845), .IN2(n12842), .QN(n12869) );
  AO221X1 U22682 ( .IN1(n4125), .IN2(n11009), .IN3(n4126), .IN4(n11010), .IN5(
        n11011), .Q(n10963) );
  INVX0 U22683 ( .IN(n10987), .QN(n4126) );
  AO22X1 U22684 ( .IN1(n11007), .IN2(n4128), .IN3(n11012), .IN4(n11010), .Q(
        n11011) );
  NOR2X0 U22685 ( .IN1(n10988), .IN2(n10985), .QN(n11012) );
  AO221X1 U22686 ( .IN1(n4080), .IN2(n10699), .IN3(n4081), .IN4(n10700), .IN5(
        n10701), .Q(n10653) );
  INVX0 U22687 ( .IN(n10677), .QN(n4081) );
  AO22X1 U22688 ( .IN1(n10697), .IN2(n4083), .IN3(n10702), .IN4(n10700), .Q(
        n10701) );
  NOR2X0 U22689 ( .IN1(n10678), .IN2(n10675), .QN(n10702) );
  AO221X1 U22690 ( .IN1(n3675), .IN2(n12557), .IN3(n3676), .IN4(n12558), .IN5(
        n12559), .Q(n12511) );
  INVX0 U22691 ( .IN(n12535), .QN(n3676) );
  AO22X1 U22692 ( .IN1(n12555), .IN2(n3678), .IN3(n12560), .IN4(n12558), .Q(
        n12559) );
  NOR2X0 U22693 ( .IN1(n12536), .IN2(n12533), .QN(n12560) );
  AO221X1 U22694 ( .IN1(n3630), .IN2(n12248), .IN3(n3631), .IN4(n12249), .IN5(
        n12250), .Q(n12202) );
  INVX0 U22695 ( .IN(n12226), .QN(n3631) );
  AO22X1 U22696 ( .IN1(n12246), .IN2(n3633), .IN3(n12251), .IN4(n12249), .Q(
        n12250) );
  NOR2X0 U22697 ( .IN1(n12227), .IN2(n12224), .QN(n12251) );
  AO221X1 U22698 ( .IN1(n4035), .IN2(n10390), .IN3(n4036), .IN4(n10391), .IN5(
        n10392), .Q(n10344) );
  INVX0 U22699 ( .IN(n10368), .QN(n4036) );
  AO22X1 U22700 ( .IN1(n10388), .IN2(n4038), .IN3(n10393), .IN4(n10391), .Q(
        n10392) );
  NOR2X0 U22701 ( .IN1(n10369), .IN2(n10366), .QN(n10393) );
  AO221X1 U22702 ( .IN1(n3990), .IN2(n10080), .IN3(n3991), .IN4(n10081), .IN5(
        n10082), .Q(n10034) );
  INVX0 U22703 ( .IN(n10058), .QN(n3991) );
  AO22X1 U22704 ( .IN1(n10078), .IN2(n3993), .IN3(n10083), .IN4(n10081), .Q(
        n10082) );
  NOR2X0 U22705 ( .IN1(n10059), .IN2(n10056), .QN(n10083) );
  AO221X1 U22706 ( .IN1(n3585), .IN2(n11938), .IN3(n3586), .IN4(n11939), .IN5(
        n11940), .Q(n11892) );
  INVX0 U22707 ( .IN(n11916), .QN(n3586) );
  AO22X1 U22708 ( .IN1(n11936), .IN2(n3588), .IN3(n11941), .IN4(n11939), .Q(
        n11940) );
  NOR2X0 U22709 ( .IN1(n11917), .IN2(n11914), .QN(n11941) );
  AO221X1 U22710 ( .IN1(n3540), .IN2(n11628), .IN3(n3541), .IN4(n11629), .IN5(
        n11630), .Q(n11582) );
  INVX0 U22711 ( .IN(n11606), .QN(n3541) );
  AO22X1 U22712 ( .IN1(n11626), .IN2(n3543), .IN3(n11631), .IN4(n11629), .Q(
        n11630) );
  NOR2X0 U22713 ( .IN1(n11607), .IN2(n11604), .QN(n11631) );
  AO221X1 U22714 ( .IN1(n3945), .IN2(n9770), .IN3(n3946), .IN4(n9771), .IN5(
        n9772), .Q(n9724) );
  INVX0 U22715 ( .IN(n9748), .QN(n3946) );
  AO22X1 U22716 ( .IN1(n9768), .IN2(n3948), .IN3(n9773), .IN4(n9771), .Q(n9772) );
  NOR2X0 U22717 ( .IN1(n9749), .IN2(n9746), .QN(n9773) );
  AO221X1 U22718 ( .IN1(n3900), .IN2(n9459), .IN3(n3901), .IN4(n9460), .IN5(
        n9461), .Q(n9413) );
  INVX0 U22719 ( .IN(n9437), .QN(n3901) );
  AO22X1 U22720 ( .IN1(n9457), .IN2(n3903), .IN3(n9462), .IN4(n9460), .Q(n9461) );
  NOR2X0 U22721 ( .IN1(n9438), .IN2(n9435), .QN(n9462) );
  AO221X1 U22722 ( .IN1(n4215), .IN2(n14057), .IN3(n4216), .IN4(n14058), .IN5(
        n14059), .Q(n14011) );
  INVX0 U22723 ( .IN(n14035), .QN(n4216) );
  AO22X1 U22724 ( .IN1(n14055), .IN2(n4218), .IN3(n14060), .IN4(n14058), .Q(
        n14059) );
  NOR2X0 U22725 ( .IN1(n14036), .IN2(n14033), .QN(n14060) );
  AO21X1 U22726 ( .IN1(n13473), .IN2(n13474), .IN3(n13471), .Q(n13431) );
  NAND3X0 U22727 ( .IN1(n13475), .IN2(n3328), .IN3(n13447), .QN(n13474) );
  AO21X1 U22728 ( .IN1(n10998), .IN2(n10999), .IN3(n10996), .Q(n10956) );
  NAND3X0 U22729 ( .IN1(n11000), .IN2(n3272), .IN3(n10972), .QN(n10999) );
  AO21X1 U22730 ( .IN1(n10379), .IN2(n10380), .IN3(n10377), .Q(n10337) );
  NAND3X0 U22731 ( .IN1(n10381), .IN2(n3288), .IN3(n10353), .QN(n10380) );
  AO21X1 U22732 ( .IN1(n9759), .IN2(n9760), .IN3(n9757), .Q(n9717) );
  NAND3X0 U22733 ( .IN1(n9761), .IN2(n3304), .IN3(n9733), .QN(n9760) );
  AO21X1 U22734 ( .IN1(n13782), .IN2(n13783), .IN3(n13780), .Q(n13740) );
  NAND3X0 U22735 ( .IN1(n13784), .IN2(n3320), .IN3(n13756), .QN(n13783) );
  AO21X1 U22736 ( .IN1(n13164), .IN2(n13165), .IN3(n13162), .Q(n13122) );
  NAND3X0 U22737 ( .IN1(n13166), .IN2(n3336), .IN3(n13138), .QN(n13165) );
  AO21X1 U22738 ( .IN1(n12855), .IN2(n12856), .IN3(n12853), .Q(n12813) );
  NAND3X0 U22739 ( .IN1(n12857), .IN2(n3344), .IN3(n12829), .QN(n12856) );
  AO21X1 U22740 ( .IN1(n12546), .IN2(n12547), .IN3(n12544), .Q(n12504) );
  NAND3X0 U22741 ( .IN1(n12548), .IN2(n3352), .IN3(n12520), .QN(n12547) );
  AO21X1 U22742 ( .IN1(n12237), .IN2(n12238), .IN3(n12235), .Q(n12195) );
  NAND3X0 U22743 ( .IN1(n12239), .IN2(n3360), .IN3(n12211), .QN(n12238) );
  AO21X1 U22744 ( .IN1(n11927), .IN2(n11928), .IN3(n11925), .Q(n11885) );
  NAND3X0 U22745 ( .IN1(n11929), .IN2(n3368), .IN3(n11901), .QN(n11928) );
  AO21X1 U22746 ( .IN1(n11617), .IN2(n11618), .IN3(n11615), .Q(n11575) );
  NAND3X0 U22747 ( .IN1(n11619), .IN2(n3376), .IN3(n11591), .QN(n11618) );
  AO21X1 U22748 ( .IN1(n11307), .IN2(n11308), .IN3(n11305), .Q(n11265) );
  NAND3X0 U22749 ( .IN1(n11309), .IN2(n3264), .IN3(n11281), .QN(n11308) );
  AO21X1 U22750 ( .IN1(n10688), .IN2(n10689), .IN3(n10686), .Q(n10646) );
  NAND3X0 U22751 ( .IN1(n10690), .IN2(n3280), .IN3(n10662), .QN(n10689) );
  AO21X1 U22752 ( .IN1(n10069), .IN2(n10070), .IN3(n10067), .Q(n10027) );
  NAND3X0 U22753 ( .IN1(n10071), .IN2(n3296), .IN3(n10043), .QN(n10070) );
  AO21X1 U22754 ( .IN1(n9448), .IN2(n9449), .IN3(n9446), .Q(n9406) );
  NAND3X0 U22755 ( .IN1(n9450), .IN2(n3312), .IN3(n9422), .QN(n9449) );
  OA21X1 U22756 ( .IN1(n13768), .IN2(n13775), .IN3(n13758), .Q(n13764) );
  OA21X1 U22757 ( .IN1(n13459), .IN2(n13466), .IN3(n13449), .Q(n13455) );
  OA21X1 U22758 ( .IN1(n11293), .IN2(n11300), .IN3(n11283), .Q(n11289) );
  OA21X1 U22759 ( .IN1(n13150), .IN2(n13157), .IN3(n13140), .Q(n13146) );
  OA21X1 U22760 ( .IN1(n12841), .IN2(n12848), .IN3(n12831), .Q(n12837) );
  OA21X1 U22761 ( .IN1(n10984), .IN2(n10991), .IN3(n10974), .Q(n10980) );
  OA21X1 U22762 ( .IN1(n10674), .IN2(n10681), .IN3(n10664), .Q(n10670) );
  OA21X1 U22763 ( .IN1(n12532), .IN2(n12539), .IN3(n12522), .Q(n12528) );
  OA21X1 U22764 ( .IN1(n12223), .IN2(n12230), .IN3(n12213), .Q(n12219) );
  OA21X1 U22765 ( .IN1(n10365), .IN2(n10372), .IN3(n10355), .Q(n10361) );
  OA21X1 U22766 ( .IN1(n10055), .IN2(n10062), .IN3(n10045), .Q(n10051) );
  OA21X1 U22767 ( .IN1(n11913), .IN2(n11920), .IN3(n11903), .Q(n11909) );
  OA21X1 U22768 ( .IN1(n11603), .IN2(n11610), .IN3(n11593), .Q(n11599) );
  OA21X1 U22769 ( .IN1(n9745), .IN2(n9752), .IN3(n9735), .Q(n9741) );
  OA21X1 U22770 ( .IN1(n9434), .IN2(n9441), .IN3(n9424), .Q(n9430) );
  OA21X1 U22771 ( .IN1(n13831), .IN2(n13838), .IN3(n13850), .Q(n13827) );
  OA21X1 U22772 ( .IN1(n13705), .IN2(n13677), .IN3(n13720), .Q(n13701) );
  OA21X1 U22773 ( .IN1(n13522), .IN2(n13529), .IN3(n13541), .Q(n13518) );
  OA21X1 U22774 ( .IN1(n13396), .IN2(n13368), .IN3(n13411), .Q(n13392) );
  OA21X1 U22775 ( .IN1(n11356), .IN2(n11363), .IN3(n11375), .Q(n11352) );
  OA21X1 U22776 ( .IN1(n11230), .IN2(n11202), .IN3(n11245), .Q(n11226) );
  OA21X1 U22777 ( .IN1(n13213), .IN2(n13220), .IN3(n13232), .Q(n13209) );
  OA21X1 U22778 ( .IN1(n13087), .IN2(n13059), .IN3(n13102), .Q(n13083) );
  OA21X1 U22779 ( .IN1(n12904), .IN2(n12911), .IN3(n12923), .Q(n12900) );
  OA21X1 U22780 ( .IN1(n12778), .IN2(n12750), .IN3(n12793), .Q(n12774) );
  OA21X1 U22781 ( .IN1(n11047), .IN2(n11054), .IN3(n11066), .Q(n11043) );
  OA21X1 U22782 ( .IN1(n10921), .IN2(n10893), .IN3(n10936), .Q(n10917) );
  OA21X1 U22783 ( .IN1(n10737), .IN2(n10744), .IN3(n10756), .Q(n10733) );
  OA21X1 U22784 ( .IN1(n10611), .IN2(n10583), .IN3(n10626), .Q(n10607) );
  OA21X1 U22785 ( .IN1(n12595), .IN2(n12602), .IN3(n12614), .Q(n12591) );
  OA21X1 U22786 ( .IN1(n12469), .IN2(n12441), .IN3(n12484), .Q(n12465) );
  OA21X1 U22787 ( .IN1(n12286), .IN2(n12293), .IN3(n12305), .Q(n12282) );
  OA21X1 U22788 ( .IN1(n12160), .IN2(n12132), .IN3(n12175), .Q(n12156) );
  OA21X1 U22789 ( .IN1(n10428), .IN2(n10435), .IN3(n10447), .Q(n10424) );
  OA21X1 U22790 ( .IN1(n10302), .IN2(n10274), .IN3(n10317), .Q(n10298) );
  OA21X1 U22791 ( .IN1(n10118), .IN2(n10125), .IN3(n10137), .Q(n10114) );
  OA21X1 U22792 ( .IN1(n9992), .IN2(n9964), .IN3(n10007), .Q(n9988) );
  OA21X1 U22793 ( .IN1(n11976), .IN2(n11983), .IN3(n11995), .Q(n11972) );
  OA21X1 U22794 ( .IN1(n11850), .IN2(n11822), .IN3(n11865), .Q(n11846) );
  OA21X1 U22795 ( .IN1(n11666), .IN2(n11673), .IN3(n11685), .Q(n11662) );
  OA21X1 U22796 ( .IN1(n11540), .IN2(n11512), .IN3(n11555), .Q(n11536) );
  OA21X1 U22797 ( .IN1(n9808), .IN2(n9815), .IN3(n9827), .Q(n9804) );
  OA21X1 U22798 ( .IN1(n9682), .IN2(n9654), .IN3(n9697), .Q(n9678) );
  OA21X1 U22799 ( .IN1(n9497), .IN2(n9504), .IN3(n9516), .Q(n9493) );
  OA21X1 U22800 ( .IN1(n9371), .IN2(n9343), .IN3(n9386), .Q(n9367) );
  AND2X1 U22801 ( .IN1(n13542), .IN2(n13543), .Q(n13522) );
  NAND3X0 U22802 ( .IN1(n18159), .IN2(n13325), .IN3(n3818), .QN(n13543) );
  AND2X1 U22803 ( .IN1(n11376), .IN2(n11377), .Q(n11356) );
  NAND3X0 U22804 ( .IN1(n18160), .IN2(n11159), .IN3(n4178), .QN(n11377) );
  AND2X1 U22805 ( .IN1(n12306), .IN2(n12307), .Q(n12286) );
  NAND3X0 U22806 ( .IN1(n18161), .IN2(n12089), .IN3(n3638), .QN(n12307) );
  AND2X1 U22807 ( .IN1(n9828), .IN2(n9829), .Q(n9808) );
  NAND3X0 U22808 ( .IN1(n18162), .IN2(n9611), .IN3(n3953), .QN(n9829) );
  ISOLANDX1 U22809 ( .D(n13728), .ISO(n13674), .Q(n13726) );
  ISOLANDX1 U22810 ( .D(n13419), .ISO(n13365), .Q(n13417) );
  ISOLANDX1 U22811 ( .D(n11253), .ISO(n11199), .Q(n11251) );
  ISOLANDX1 U22812 ( .D(n13110), .ISO(n13056), .Q(n13108) );
  ISOLANDX1 U22813 ( .D(n12801), .ISO(n12747), .Q(n12799) );
  ISOLANDX1 U22814 ( .D(n10944), .ISO(n10890), .Q(n10942) );
  ISOLANDX1 U22815 ( .D(n10634), .ISO(n10580), .Q(n10632) );
  ISOLANDX1 U22816 ( .D(n12492), .ISO(n12438), .Q(n12490) );
  ISOLANDX1 U22817 ( .D(n12183), .ISO(n12129), .Q(n12181) );
  ISOLANDX1 U22818 ( .D(n10325), .ISO(n10271), .Q(n10323) );
  ISOLANDX1 U22819 ( .D(n10015), .ISO(n9961), .Q(n10013) );
  ISOLANDX1 U22820 ( .D(n11873), .ISO(n11819), .Q(n11871) );
  ISOLANDX1 U22821 ( .D(n11563), .ISO(n11509), .Q(n11561) );
  ISOLANDX1 U22822 ( .D(n9705), .ISO(n9651), .Q(n9703) );
  ISOLANDX1 U22823 ( .D(n9394), .ISO(n9340), .Q(n9392) );
  ISOLANDX1 U22824 ( .D(n13859), .ISO(n13818), .Q(n13857) );
  ISOLANDX1 U22825 ( .D(n13550), .ISO(n13509), .Q(n13548) );
  ISOLANDX1 U22826 ( .D(n11384), .ISO(n11343), .Q(n11382) );
  ISOLANDX1 U22827 ( .D(n13241), .ISO(n13200), .Q(n13239) );
  ISOLANDX1 U22828 ( .D(n12932), .ISO(n12891), .Q(n12930) );
  ISOLANDX1 U22829 ( .D(n11075), .ISO(n11034), .Q(n11073) );
  ISOLANDX1 U22830 ( .D(n10765), .ISO(n10724), .Q(n10763) );
  ISOLANDX1 U22831 ( .D(n12623), .ISO(n12582), .Q(n12621) );
  ISOLANDX1 U22832 ( .D(n12314), .ISO(n12273), .Q(n12312) );
  ISOLANDX1 U22833 ( .D(n10456), .ISO(n10415), .Q(n10454) );
  ISOLANDX1 U22834 ( .D(n10146), .ISO(n10105), .Q(n10144) );
  ISOLANDX1 U22835 ( .D(n12004), .ISO(n11963), .Q(n12002) );
  ISOLANDX1 U22836 ( .D(n11694), .ISO(n11653), .Q(n11692) );
  ISOLANDX1 U22837 ( .D(n9836), .ISO(n9795), .Q(n9834) );
  ISOLANDX1 U22838 ( .D(n9525), .ISO(n9484), .Q(n9523) );
  ISOLANDX1 U22839 ( .D(n13793), .ISO(n13754), .Q(n13794) );
  ISOLANDX1 U22840 ( .D(n13484), .ISO(n13445), .Q(n13485) );
  ISOLANDX1 U22841 ( .D(n11318), .ISO(n11279), .Q(n11319) );
  ISOLANDX1 U22842 ( .D(n13175), .ISO(n13136), .Q(n13176) );
  ISOLANDX1 U22843 ( .D(n12866), .ISO(n12827), .Q(n12867) );
  ISOLANDX1 U22844 ( .D(n11009), .ISO(n10970), .Q(n11010) );
  ISOLANDX1 U22845 ( .D(n10699), .ISO(n10660), .Q(n10700) );
  ISOLANDX1 U22846 ( .D(n12557), .ISO(n12518), .Q(n12558) );
  ISOLANDX1 U22847 ( .D(n12248), .ISO(n12209), .Q(n12249) );
  ISOLANDX1 U22848 ( .D(n10390), .ISO(n10351), .Q(n10391) );
  ISOLANDX1 U22849 ( .D(n10080), .ISO(n10041), .Q(n10081) );
  ISOLANDX1 U22850 ( .D(n11938), .ISO(n11899), .Q(n11939) );
  ISOLANDX1 U22851 ( .D(n11628), .ISO(n11589), .Q(n11629) );
  ISOLANDX1 U22852 ( .D(n9770), .ISO(n9731), .Q(n9771) );
  ISOLANDX1 U22853 ( .D(n9459), .ISO(n9420), .Q(n9460) );
  ISOLANDX1 U22854 ( .D(n14057), .ISO(n14018), .Q(n14058) );
  OA21X1 U22855 ( .IN1(n13847), .IN2(n13848), .IN3(n13849), .Q(n13842) );
  OA21X1 U22856 ( .IN1(n13838), .IN2(n13830), .IN3(n13827), .Q(n13848) );
  OA21X1 U22857 ( .IN1(n13676), .IN2(n13718), .IN3(n13719), .Q(n13713) );
  OA21X1 U22858 ( .IN1(n13677), .IN2(n13704), .IN3(n13701), .Q(n13718) );
  OA21X1 U22859 ( .IN1(n13538), .IN2(n13539), .IN3(n13540), .Q(n13533) );
  OA21X1 U22860 ( .IN1(n13529), .IN2(n13521), .IN3(n13518), .Q(n13539) );
  OA21X1 U22861 ( .IN1(n13477), .IN2(n13478), .IN3(n13479), .Q(n13470) );
  OA21X1 U22862 ( .IN1(n13466), .IN2(n13458), .IN3(n13455), .Q(n13478) );
  OA21X1 U22863 ( .IN1(n13367), .IN2(n13409), .IN3(n13410), .Q(n13404) );
  OA21X1 U22864 ( .IN1(n13368), .IN2(n13395), .IN3(n13392), .Q(n13409) );
  OA21X1 U22865 ( .IN1(n11372), .IN2(n11373), .IN3(n11374), .Q(n11367) );
  OA21X1 U22866 ( .IN1(n11363), .IN2(n11355), .IN3(n11352), .Q(n11373) );
  OA21X1 U22867 ( .IN1(n11201), .IN2(n11243), .IN3(n11244), .Q(n11238) );
  OA21X1 U22868 ( .IN1(n11202), .IN2(n11229), .IN3(n11226), .Q(n11243) );
  OA21X1 U22869 ( .IN1(n13229), .IN2(n13230), .IN3(n13231), .Q(n13224) );
  OA21X1 U22870 ( .IN1(n13220), .IN2(n13212), .IN3(n13209), .Q(n13230) );
  OA21X1 U22871 ( .IN1(n13058), .IN2(n13100), .IN3(n13101), .Q(n13095) );
  OA21X1 U22872 ( .IN1(n13059), .IN2(n13086), .IN3(n13083), .Q(n13100) );
  OA21X1 U22873 ( .IN1(n12920), .IN2(n12921), .IN3(n12922), .Q(n12915) );
  OA21X1 U22874 ( .IN1(n12911), .IN2(n12903), .IN3(n12900), .Q(n12921) );
  OA21X1 U22875 ( .IN1(n12749), .IN2(n12791), .IN3(n12792), .Q(n12786) );
  OA21X1 U22876 ( .IN1(n12750), .IN2(n12777), .IN3(n12774), .Q(n12791) );
  OA21X1 U22877 ( .IN1(n11063), .IN2(n11064), .IN3(n11065), .Q(n11058) );
  OA21X1 U22878 ( .IN1(n11054), .IN2(n11046), .IN3(n11043), .Q(n11064) );
  OA21X1 U22879 ( .IN1(n11002), .IN2(n11003), .IN3(n11004), .Q(n10995) );
  OA21X1 U22880 ( .IN1(n10991), .IN2(n10983), .IN3(n10980), .Q(n11003) );
  OA21X1 U22881 ( .IN1(n10892), .IN2(n10934), .IN3(n10935), .Q(n10929) );
  OA21X1 U22882 ( .IN1(n10893), .IN2(n10920), .IN3(n10917), .Q(n10934) );
  OA21X1 U22883 ( .IN1(n10753), .IN2(n10754), .IN3(n10755), .Q(n10748) );
  OA21X1 U22884 ( .IN1(n10744), .IN2(n10736), .IN3(n10733), .Q(n10754) );
  OA21X1 U22885 ( .IN1(n10582), .IN2(n10624), .IN3(n10625), .Q(n10619) );
  OA21X1 U22886 ( .IN1(n10583), .IN2(n10610), .IN3(n10607), .Q(n10624) );
  OA21X1 U22887 ( .IN1(n12611), .IN2(n12612), .IN3(n12613), .Q(n12606) );
  OA21X1 U22888 ( .IN1(n12602), .IN2(n12594), .IN3(n12591), .Q(n12612) );
  OA21X1 U22889 ( .IN1(n12440), .IN2(n12482), .IN3(n12483), .Q(n12477) );
  OA21X1 U22890 ( .IN1(n12441), .IN2(n12468), .IN3(n12465), .Q(n12482) );
  OA21X1 U22891 ( .IN1(n12302), .IN2(n12303), .IN3(n12304), .Q(n12297) );
  OA21X1 U22892 ( .IN1(n12293), .IN2(n12285), .IN3(n12282), .Q(n12303) );
  OA21X1 U22893 ( .IN1(n12131), .IN2(n12173), .IN3(n12174), .Q(n12168) );
  OA21X1 U22894 ( .IN1(n12132), .IN2(n12159), .IN3(n12156), .Q(n12173) );
  OA21X1 U22895 ( .IN1(n10444), .IN2(n10445), .IN3(n10446), .Q(n10439) );
  OA21X1 U22896 ( .IN1(n10435), .IN2(n10427), .IN3(n10424), .Q(n10445) );
  OA21X1 U22897 ( .IN1(n10383), .IN2(n10384), .IN3(n10385), .Q(n10376) );
  OA21X1 U22898 ( .IN1(n10372), .IN2(n10364), .IN3(n10361), .Q(n10384) );
  OA21X1 U22899 ( .IN1(n10273), .IN2(n10315), .IN3(n10316), .Q(n10310) );
  OA21X1 U22900 ( .IN1(n10274), .IN2(n10301), .IN3(n10298), .Q(n10315) );
  OA21X1 U22901 ( .IN1(n10134), .IN2(n10135), .IN3(n10136), .Q(n10129) );
  OA21X1 U22902 ( .IN1(n10125), .IN2(n10117), .IN3(n10114), .Q(n10135) );
  OA21X1 U22903 ( .IN1(n9963), .IN2(n10005), .IN3(n10006), .Q(n10000) );
  OA21X1 U22904 ( .IN1(n9964), .IN2(n9991), .IN3(n9988), .Q(n10005) );
  OA21X1 U22905 ( .IN1(n11992), .IN2(n11993), .IN3(n11994), .Q(n11987) );
  OA21X1 U22906 ( .IN1(n11983), .IN2(n11975), .IN3(n11972), .Q(n11993) );
  OA21X1 U22907 ( .IN1(n11821), .IN2(n11863), .IN3(n11864), .Q(n11858) );
  OA21X1 U22908 ( .IN1(n11822), .IN2(n11849), .IN3(n11846), .Q(n11863) );
  OA21X1 U22909 ( .IN1(n11682), .IN2(n11683), .IN3(n11684), .Q(n11677) );
  OA21X1 U22910 ( .IN1(n11673), .IN2(n11665), .IN3(n11662), .Q(n11683) );
  OA21X1 U22911 ( .IN1(n11511), .IN2(n11553), .IN3(n11554), .Q(n11548) );
  OA21X1 U22912 ( .IN1(n11512), .IN2(n11539), .IN3(n11536), .Q(n11553) );
  OA21X1 U22913 ( .IN1(n9824), .IN2(n9825), .IN3(n9826), .Q(n9819) );
  OA21X1 U22914 ( .IN1(n9815), .IN2(n9807), .IN3(n9804), .Q(n9825) );
  OA21X1 U22915 ( .IN1(n9763), .IN2(n9764), .IN3(n9765), .Q(n9756) );
  OA21X1 U22916 ( .IN1(n9752), .IN2(n9744), .IN3(n9741), .Q(n9764) );
  OA21X1 U22917 ( .IN1(n9653), .IN2(n9695), .IN3(n9696), .Q(n9690) );
  OA21X1 U22918 ( .IN1(n9654), .IN2(n9681), .IN3(n9678), .Q(n9695) );
  OA21X1 U22919 ( .IN1(n9513), .IN2(n9514), .IN3(n9515), .Q(n9508) );
  OA21X1 U22920 ( .IN1(n9504), .IN2(n9496), .IN3(n9493), .Q(n9514) );
  OA21X1 U22921 ( .IN1(n9342), .IN2(n9384), .IN3(n9385), .Q(n9379) );
  OA21X1 U22922 ( .IN1(n9343), .IN2(n9370), .IN3(n9367), .Q(n9384) );
  NAND3X0 U22923 ( .IN1(n13775), .IN2(n13756), .IN3(n3319), .QN(n13746) );
  NAND3X0 U22924 ( .IN1(n13466), .IN2(n13447), .IN3(n3327), .QN(n13437) );
  NAND3X0 U22925 ( .IN1(n11300), .IN2(n11281), .IN3(n3263), .QN(n11271) );
  NAND3X0 U22926 ( .IN1(n13157), .IN2(n13138), .IN3(n3335), .QN(n13128) );
  NAND3X0 U22927 ( .IN1(n12848), .IN2(n12829), .IN3(n3343), .QN(n12819) );
  NAND3X0 U22928 ( .IN1(n10991), .IN2(n10972), .IN3(n3271), .QN(n10962) );
  NAND3X0 U22929 ( .IN1(n10681), .IN2(n10662), .IN3(n3279), .QN(n10652) );
  NAND3X0 U22930 ( .IN1(n12539), .IN2(n12520), .IN3(n3351), .QN(n12510) );
  NAND3X0 U22931 ( .IN1(n12230), .IN2(n12211), .IN3(n3359), .QN(n12201) );
  NAND3X0 U22932 ( .IN1(n10372), .IN2(n10353), .IN3(n3287), .QN(n10343) );
  NAND3X0 U22933 ( .IN1(n10062), .IN2(n10043), .IN3(n3295), .QN(n10033) );
  NAND3X0 U22934 ( .IN1(n11920), .IN2(n11901), .IN3(n3367), .QN(n11891) );
  NAND3X0 U22935 ( .IN1(n11610), .IN2(n11591), .IN3(n3375), .QN(n11581) );
  NAND3X0 U22936 ( .IN1(n9752), .IN2(n9733), .IN3(n3303), .QN(n9723) );
  NAND3X0 U22937 ( .IN1(n9441), .IN2(n9422), .IN3(n3311), .QN(n9412) );
  NAND3X0 U22938 ( .IN1(n14039), .IN2(n14020), .IN3(n3253), .QN(n14010) );
  OA21X1 U22939 ( .IN1(n13786), .IN2(n13787), .IN3(n13788), .Q(n13779) );
  OA21X1 U22940 ( .IN1(n13775), .IN2(n13767), .IN3(n13764), .Q(n13787) );
  OA21X1 U22941 ( .IN1(n11311), .IN2(n11312), .IN3(n11313), .Q(n11304) );
  OA21X1 U22942 ( .IN1(n11300), .IN2(n11292), .IN3(n11289), .Q(n11312) );
  OA21X1 U22943 ( .IN1(n13168), .IN2(n13169), .IN3(n13170), .Q(n13161) );
  OA21X1 U22944 ( .IN1(n13157), .IN2(n13149), .IN3(n13146), .Q(n13169) );
  OA21X1 U22945 ( .IN1(n12859), .IN2(n12860), .IN3(n12861), .Q(n12852) );
  OA21X1 U22946 ( .IN1(n12848), .IN2(n12840), .IN3(n12837), .Q(n12860) );
  OA21X1 U22947 ( .IN1(n10692), .IN2(n10693), .IN3(n10694), .Q(n10685) );
  OA21X1 U22948 ( .IN1(n10681), .IN2(n10673), .IN3(n10670), .Q(n10693) );
  OA21X1 U22949 ( .IN1(n12550), .IN2(n12551), .IN3(n12552), .Q(n12543) );
  OA21X1 U22950 ( .IN1(n12539), .IN2(n12531), .IN3(n12528), .Q(n12551) );
  OA21X1 U22951 ( .IN1(n12241), .IN2(n12242), .IN3(n12243), .Q(n12234) );
  OA21X1 U22952 ( .IN1(n12230), .IN2(n12222), .IN3(n12219), .Q(n12242) );
  OA21X1 U22953 ( .IN1(n10073), .IN2(n10074), .IN3(n10075), .Q(n10066) );
  OA21X1 U22954 ( .IN1(n10062), .IN2(n10054), .IN3(n10051), .Q(n10074) );
  OA21X1 U22955 ( .IN1(n11931), .IN2(n11932), .IN3(n11933), .Q(n11924) );
  OA21X1 U22956 ( .IN1(n11920), .IN2(n11912), .IN3(n11909), .Q(n11932) );
  OA21X1 U22957 ( .IN1(n11621), .IN2(n11622), .IN3(n11623), .Q(n11614) );
  OA21X1 U22958 ( .IN1(n11610), .IN2(n11602), .IN3(n11599), .Q(n11622) );
  OA21X1 U22959 ( .IN1(n9452), .IN2(n9453), .IN3(n9454), .Q(n9445) );
  OA21X1 U22960 ( .IN1(n9441), .IN2(n9433), .IN3(n9430), .Q(n9453) );
  OA21X1 U22961 ( .IN1(n14050), .IN2(n14051), .IN3(n14052), .Q(n14043) );
  OA21X1 U22962 ( .IN1(n14039), .IN2(n14031), .IN3(n14028), .Q(n14051) );
  AOI221X1 U22963 ( .IN1(n13853), .IN2(n13854), .IN3(n13818), .IN4(n13855), 
        .IN5(n13821), .QN(n13823) );
  NOR2X0 U22964 ( .IN1(n13838), .IN2(n13851), .QN(n13853) );
  AO221X1 U22965 ( .IN1(n13814), .IN2(n3866), .IN3(n2975), .IN4(n3223), .IN5(
        n13860), .Q(n13855) );
  INVX0 U22966 ( .IN(n13829), .QN(n2975) );
  AOI221X1 U22967 ( .IN1(n13723), .IN2(n13678), .IN3(n13674), .IN4(n13724), 
        .IN5(n13695), .QN(n13697) );
  NOR2X0 U22968 ( .IN1(n13677), .IN2(n13721), .QN(n13723) );
  AO221X1 U22969 ( .IN1(n13689), .IN2(n3874), .IN3(n2967), .IN4(n3221), .IN5(
        n13729), .Q(n13724) );
  INVX0 U22970 ( .IN(n13703), .QN(n2967) );
  AOI221X1 U22971 ( .IN1(n13544), .IN2(n13545), .IN3(n13509), .IN4(n13546), 
        .IN5(n13512), .QN(n13514) );
  NOR2X0 U22972 ( .IN1(n13529), .IN2(n13542), .QN(n13544) );
  AO221X1 U22973 ( .IN1(n13505), .IN2(n3821), .IN3(n2991), .IN4(n3227), .IN5(
        n13551), .Q(n13546) );
  INVX0 U22974 ( .IN(n13520), .QN(n2991) );
  AOI221X1 U22975 ( .IN1(n13414), .IN2(n13369), .IN3(n13365), .IN4(n13415), 
        .IN5(n13386), .QN(n13388) );
  NOR2X0 U22976 ( .IN1(n13368), .IN2(n13412), .QN(n13414) );
  AO221X1 U22977 ( .IN1(n13380), .IN2(n3829), .IN3(n2983), .IN4(n3225), .IN5(
        n13420), .Q(n13415) );
  INVX0 U22978 ( .IN(n13394), .QN(n2983) );
  AOI221X1 U22979 ( .IN1(n11378), .IN2(n11379), .IN3(n11343), .IN4(n11380), 
        .IN5(n11346), .QN(n11348) );
  NOR2X0 U22980 ( .IN1(n11363), .IN2(n11376), .QN(n11378) );
  AO221X1 U22981 ( .IN1(n11339), .IN2(n4181), .IN3(n2863), .IN4(n3195), .IN5(
        n11385), .Q(n11380) );
  INVX0 U22982 ( .IN(n11354), .QN(n2863) );
  AOI221X1 U22983 ( .IN1(n11248), .IN2(n11203), .IN3(n11199), .IN4(n11249), 
        .IN5(n11220), .QN(n11222) );
  NOR2X0 U22984 ( .IN1(n11202), .IN2(n11246), .QN(n11248) );
  AO221X1 U22985 ( .IN1(n11214), .IN2(n4189), .IN3(n2855), .IN4(n3193), .IN5(
        n11254), .Q(n11249) );
  INVX0 U22986 ( .IN(n11228), .QN(n2855) );
  AOI221X1 U22987 ( .IN1(n13235), .IN2(n13236), .IN3(n13200), .IN4(n13237), 
        .IN5(n13203), .QN(n13205) );
  NOR2X0 U22988 ( .IN1(n13220), .IN2(n13233), .QN(n13235) );
  AO221X1 U22989 ( .IN1(n13196), .IN2(n3776), .IN3(n3007), .IN4(n3231), .IN5(
        n13242), .Q(n13237) );
  INVX0 U22990 ( .IN(n13211), .QN(n3007) );
  AOI221X1 U22991 ( .IN1(n13105), .IN2(n13060), .IN3(n13056), .IN4(n13106), 
        .IN5(n13077), .QN(n13079) );
  NOR2X0 U22992 ( .IN1(n13059), .IN2(n13103), .QN(n13105) );
  AO221X1 U22993 ( .IN1(n13071), .IN2(n3784), .IN3(n2999), .IN4(n3229), .IN5(
        n13111), .Q(n13106) );
  INVX0 U22994 ( .IN(n13085), .QN(n2999) );
  AOI221X1 U22995 ( .IN1(n12926), .IN2(n12927), .IN3(n12891), .IN4(n12928), 
        .IN5(n12894), .QN(n12896) );
  NOR2X0 U22996 ( .IN1(n12911), .IN2(n12924), .QN(n12926) );
  AO221X1 U22997 ( .IN1(n12887), .IN2(n3731), .IN3(n3023), .IN4(n3235), .IN5(
        n12933), .Q(n12928) );
  INVX0 U22998 ( .IN(n12902), .QN(n3023) );
  AOI221X1 U22999 ( .IN1(n12796), .IN2(n12751), .IN3(n12747), .IN4(n12797), 
        .IN5(n12768), .QN(n12770) );
  NOR2X0 U23000 ( .IN1(n12750), .IN2(n12794), .QN(n12796) );
  AO221X1 U23001 ( .IN1(n12762), .IN2(n3739), .IN3(n3015), .IN4(n3233), .IN5(
        n12802), .Q(n12797) );
  INVX0 U23002 ( .IN(n12776), .QN(n3015) );
  AOI221X1 U23003 ( .IN1(n11069), .IN2(n11070), .IN3(n11034), .IN4(n11071), 
        .IN5(n11037), .QN(n11039) );
  NOR2X0 U23004 ( .IN1(n11054), .IN2(n11067), .QN(n11069) );
  AO221X1 U23005 ( .IN1(n11030), .IN2(n4136), .IN3(n2879), .IN4(n3199), .IN5(
        n11076), .Q(n11071) );
  INVX0 U23006 ( .IN(n11045), .QN(n2879) );
  AOI221X1 U23007 ( .IN1(n10939), .IN2(n10894), .IN3(n10890), .IN4(n10940), 
        .IN5(n10911), .QN(n10913) );
  NOR2X0 U23008 ( .IN1(n10893), .IN2(n10937), .QN(n10939) );
  AO221X1 U23009 ( .IN1(n10905), .IN2(n4144), .IN3(n2871), .IN4(n3197), .IN5(
        n10945), .Q(n10940) );
  INVX0 U23010 ( .IN(n10919), .QN(n2871) );
  AOI221X1 U23011 ( .IN1(n10759), .IN2(n10760), .IN3(n10724), .IN4(n10761), 
        .IN5(n10727), .QN(n10729) );
  NOR2X0 U23012 ( .IN1(n10744), .IN2(n10757), .QN(n10759) );
  AO221X1 U23013 ( .IN1(n10720), .IN2(n4091), .IN3(n2895), .IN4(n3203), .IN5(
        n10766), .Q(n10761) );
  INVX0 U23014 ( .IN(n10735), .QN(n2895) );
  AOI221X1 U23015 ( .IN1(n10629), .IN2(n10584), .IN3(n10580), .IN4(n10630), 
        .IN5(n10601), .QN(n10603) );
  NOR2X0 U23016 ( .IN1(n10583), .IN2(n10627), .QN(n10629) );
  AO221X1 U23017 ( .IN1(n10595), .IN2(n4099), .IN3(n2887), .IN4(n3201), .IN5(
        n10635), .Q(n10630) );
  INVX0 U23018 ( .IN(n10609), .QN(n2887) );
  AOI221X1 U23019 ( .IN1(n12617), .IN2(n12618), .IN3(n12582), .IN4(n12619), 
        .IN5(n12585), .QN(n12587) );
  NOR2X0 U23020 ( .IN1(n12602), .IN2(n12615), .QN(n12617) );
  AO221X1 U23021 ( .IN1(n12578), .IN2(n3686), .IN3(n3039), .IN4(n3239), .IN5(
        n12624), .Q(n12619) );
  INVX0 U23022 ( .IN(n12593), .QN(n3039) );
  AOI221X1 U23023 ( .IN1(n12487), .IN2(n12442), .IN3(n12438), .IN4(n12488), 
        .IN5(n12459), .QN(n12461) );
  NOR2X0 U23024 ( .IN1(n12441), .IN2(n12485), .QN(n12487) );
  AO221X1 U23025 ( .IN1(n12453), .IN2(n3694), .IN3(n3031), .IN4(n3237), .IN5(
        n12493), .Q(n12488) );
  INVX0 U23026 ( .IN(n12467), .QN(n3031) );
  AOI221X1 U23027 ( .IN1(n12308), .IN2(n12309), .IN3(n12273), .IN4(n12310), 
        .IN5(n12276), .QN(n12278) );
  NOR2X0 U23028 ( .IN1(n12293), .IN2(n12306), .QN(n12308) );
  AO221X1 U23029 ( .IN1(n12269), .IN2(n3641), .IN3(n3055), .IN4(n3243), .IN5(
        n12315), .Q(n12310) );
  INVX0 U23030 ( .IN(n12284), .QN(n3055) );
  AOI221X1 U23031 ( .IN1(n12178), .IN2(n12133), .IN3(n12129), .IN4(n12179), 
        .IN5(n12150), .QN(n12152) );
  NOR2X0 U23032 ( .IN1(n12132), .IN2(n12176), .QN(n12178) );
  AO221X1 U23033 ( .IN1(n12144), .IN2(n3649), .IN3(n3047), .IN4(n3241), .IN5(
        n12184), .Q(n12179) );
  INVX0 U23034 ( .IN(n12158), .QN(n3047) );
  AOI221X1 U23035 ( .IN1(n10450), .IN2(n10451), .IN3(n10415), .IN4(n10452), 
        .IN5(n10418), .QN(n10420) );
  NOR2X0 U23036 ( .IN1(n10435), .IN2(n10448), .QN(n10450) );
  AO221X1 U23037 ( .IN1(n10411), .IN2(n4046), .IN3(n2911), .IN4(n3207), .IN5(
        n10457), .Q(n10452) );
  INVX0 U23038 ( .IN(n10426), .QN(n2911) );
  AOI221X1 U23039 ( .IN1(n10320), .IN2(n10275), .IN3(n10271), .IN4(n10321), 
        .IN5(n10292), .QN(n10294) );
  NOR2X0 U23040 ( .IN1(n10274), .IN2(n10318), .QN(n10320) );
  AO221X1 U23041 ( .IN1(n10286), .IN2(n4054), .IN3(n2903), .IN4(n3205), .IN5(
        n10326), .Q(n10321) );
  INVX0 U23042 ( .IN(n10300), .QN(n2903) );
  AOI221X1 U23043 ( .IN1(n10140), .IN2(n10141), .IN3(n10105), .IN4(n10142), 
        .IN5(n10108), .QN(n10110) );
  NOR2X0 U23044 ( .IN1(n10125), .IN2(n10138), .QN(n10140) );
  AO221X1 U23045 ( .IN1(n10101), .IN2(n4001), .IN3(n2927), .IN4(n3211), .IN5(
        n10147), .Q(n10142) );
  INVX0 U23046 ( .IN(n10116), .QN(n2927) );
  AOI221X1 U23047 ( .IN1(n10010), .IN2(n9965), .IN3(n9961), .IN4(n10011), 
        .IN5(n9982), .QN(n9984) );
  NOR2X0 U23048 ( .IN1(n9964), .IN2(n10008), .QN(n10010) );
  AO221X1 U23049 ( .IN1(n9976), .IN2(n4009), .IN3(n2919), .IN4(n3209), .IN5(
        n10016), .Q(n10011) );
  INVX0 U23050 ( .IN(n9990), .QN(n2919) );
  AOI221X1 U23051 ( .IN1(n11998), .IN2(n11999), .IN3(n11963), .IN4(n12000), 
        .IN5(n11966), .QN(n11968) );
  NOR2X0 U23052 ( .IN1(n11983), .IN2(n11996), .QN(n11998) );
  AO221X1 U23053 ( .IN1(n11959), .IN2(n3596), .IN3(n3071), .IN4(n3247), .IN5(
        n12005), .Q(n12000) );
  INVX0 U23054 ( .IN(n11974), .QN(n3071) );
  AOI221X1 U23055 ( .IN1(n11868), .IN2(n11823), .IN3(n11819), .IN4(n11869), 
        .IN5(n11840), .QN(n11842) );
  NOR2X0 U23056 ( .IN1(n11822), .IN2(n11866), .QN(n11868) );
  AO221X1 U23057 ( .IN1(n11834), .IN2(n3604), .IN3(n3063), .IN4(n3245), .IN5(
        n11874), .Q(n11869) );
  INVX0 U23058 ( .IN(n11848), .QN(n3063) );
  AOI221X1 U23059 ( .IN1(n11688), .IN2(n11689), .IN3(n11653), .IN4(n11690), 
        .IN5(n11656), .QN(n11658) );
  NOR2X0 U23060 ( .IN1(n11673), .IN2(n11686), .QN(n11688) );
  AO221X1 U23061 ( .IN1(n11649), .IN2(n3551), .IN3(n3087), .IN4(n3251), .IN5(
        n11695), .Q(n11690) );
  INVX0 U23062 ( .IN(n11664), .QN(n3087) );
  AOI221X1 U23063 ( .IN1(n11558), .IN2(n11513), .IN3(n11509), .IN4(n11559), 
        .IN5(n11530), .QN(n11532) );
  NOR2X0 U23064 ( .IN1(n11512), .IN2(n11556), .QN(n11558) );
  AO221X1 U23065 ( .IN1(n11524), .IN2(n3559), .IN3(n3079), .IN4(n3249), .IN5(
        n11564), .Q(n11559) );
  INVX0 U23066 ( .IN(n11538), .QN(n3079) );
  AOI221X1 U23067 ( .IN1(n9830), .IN2(n9831), .IN3(n9795), .IN4(n9832), .IN5(
        n9798), .QN(n9800) );
  NOR2X0 U23068 ( .IN1(n9815), .IN2(n9828), .QN(n9830) );
  AO221X1 U23069 ( .IN1(n9791), .IN2(n3956), .IN3(n2943), .IN4(n3215), .IN5(
        n9837), .Q(n9832) );
  INVX0 U23070 ( .IN(n9806), .QN(n2943) );
  AOI221X1 U23071 ( .IN1(n9700), .IN2(n9655), .IN3(n9651), .IN4(n9701), .IN5(
        n9672), .QN(n9674) );
  NOR2X0 U23072 ( .IN1(n9654), .IN2(n9698), .QN(n9700) );
  AO221X1 U23073 ( .IN1(n9666), .IN2(n3964), .IN3(n2935), .IN4(n3213), .IN5(
        n9706), .Q(n9701) );
  INVX0 U23074 ( .IN(n9680), .QN(n2935) );
  AOI221X1 U23075 ( .IN1(n9519), .IN2(n9520), .IN3(n9484), .IN4(n9521), .IN5(
        n9487), .QN(n9489) );
  NOR2X0 U23076 ( .IN1(n9504), .IN2(n9517), .QN(n9519) );
  AO221X1 U23077 ( .IN1(n9480), .IN2(n3911), .IN3(n2959), .IN4(n3219), .IN5(
        n9526), .Q(n9521) );
  INVX0 U23078 ( .IN(n9495), .QN(n2959) );
  AOI221X1 U23079 ( .IN1(n9389), .IN2(n9344), .IN3(n9340), .IN4(n9390), .IN5(
        n9361), .QN(n9363) );
  NOR2X0 U23080 ( .IN1(n9343), .IN2(n9387), .QN(n9389) );
  AO221X1 U23081 ( .IN1(n9355), .IN2(n3919), .IN3(n2951), .IN4(n3217), .IN5(
        n9395), .Q(n9390) );
  INVX0 U23082 ( .IN(n9369), .QN(n2951) );
  AOI221X1 U23083 ( .IN1(n13790), .IN2(n13791), .IN3(n13754), .IN4(n13792), 
        .IN5(n13747), .QN(n13760) );
  ISOLANDX1 U23084 ( .D(n13789), .ISO(n13775), .Q(n13790) );
  AO221X1 U23085 ( .IN1(n13756), .IN2(n3858), .IN3(n2972), .IN4(n3222), .IN5(
        n13797), .Q(n13792) );
  INVX0 U23086 ( .IN(n13766), .QN(n2972) );
  AOI221X1 U23087 ( .IN1(n13481), .IN2(n13482), .IN3(n13445), .IN4(n13483), 
        .IN5(n13438), .QN(n13451) );
  ISOLANDX1 U23088 ( .D(n13480), .ISO(n13466), .Q(n13481) );
  AO221X1 U23089 ( .IN1(n13447), .IN2(n3813), .IN3(n2988), .IN4(n3226), .IN5(
        n13488), .Q(n13483) );
  INVX0 U23090 ( .IN(n13457), .QN(n2988) );
  AOI221X1 U23091 ( .IN1(n11315), .IN2(n11316), .IN3(n11279), .IN4(n11317), 
        .IN5(n11272), .QN(n11285) );
  ISOLANDX1 U23092 ( .D(n11314), .ISO(n11300), .Q(n11315) );
  AO221X1 U23093 ( .IN1(n11281), .IN2(n4173), .IN3(n2860), .IN4(n3194), .IN5(
        n11322), .Q(n11317) );
  INVX0 U23094 ( .IN(n11291), .QN(n2860) );
  AOI221X1 U23095 ( .IN1(n13172), .IN2(n13173), .IN3(n13136), .IN4(n13174), 
        .IN5(n13129), .QN(n13142) );
  ISOLANDX1 U23096 ( .D(n13171), .ISO(n13157), .Q(n13172) );
  AO221X1 U23097 ( .IN1(n13138), .IN2(n3768), .IN3(n3004), .IN4(n3230), .IN5(
        n13179), .Q(n13174) );
  INVX0 U23098 ( .IN(n13148), .QN(n3004) );
  AOI221X1 U23099 ( .IN1(n12863), .IN2(n12864), .IN3(n12827), .IN4(n12865), 
        .IN5(n12820), .QN(n12833) );
  ISOLANDX1 U23100 ( .D(n12862), .ISO(n12848), .Q(n12863) );
  AO221X1 U23101 ( .IN1(n12829), .IN2(n3723), .IN3(n3020), .IN4(n3234), .IN5(
        n12870), .Q(n12865) );
  INVX0 U23102 ( .IN(n12839), .QN(n3020) );
  AOI221X1 U23103 ( .IN1(n11006), .IN2(n11007), .IN3(n10970), .IN4(n11008), 
        .IN5(n10963), .QN(n10976) );
  ISOLANDX1 U23104 ( .D(n11005), .ISO(n10991), .Q(n11006) );
  AO221X1 U23105 ( .IN1(n10972), .IN2(n4128), .IN3(n2876), .IN4(n3198), .IN5(
        n11013), .Q(n11008) );
  INVX0 U23106 ( .IN(n10982), .QN(n2876) );
  AOI221X1 U23107 ( .IN1(n10696), .IN2(n10697), .IN3(n10660), .IN4(n10698), 
        .IN5(n10653), .QN(n10666) );
  ISOLANDX1 U23108 ( .D(n10695), .ISO(n10681), .Q(n10696) );
  AO221X1 U23109 ( .IN1(n10662), .IN2(n4083), .IN3(n2892), .IN4(n3202), .IN5(
        n10703), .Q(n10698) );
  INVX0 U23110 ( .IN(n10672), .QN(n2892) );
  AOI221X1 U23111 ( .IN1(n12554), .IN2(n12555), .IN3(n12518), .IN4(n12556), 
        .IN5(n12511), .QN(n12524) );
  ISOLANDX1 U23112 ( .D(n12553), .ISO(n12539), .Q(n12554) );
  AO221X1 U23113 ( .IN1(n12520), .IN2(n3678), .IN3(n3036), .IN4(n3238), .IN5(
        n12561), .Q(n12556) );
  INVX0 U23114 ( .IN(n12530), .QN(n3036) );
  AOI221X1 U23115 ( .IN1(n12245), .IN2(n12246), .IN3(n12209), .IN4(n12247), 
        .IN5(n12202), .QN(n12215) );
  ISOLANDX1 U23116 ( .D(n12244), .ISO(n12230), .Q(n12245) );
  AO221X1 U23117 ( .IN1(n12211), .IN2(n3633), .IN3(n3052), .IN4(n3242), .IN5(
        n12252), .Q(n12247) );
  INVX0 U23118 ( .IN(n12221), .QN(n3052) );
  AOI221X1 U23119 ( .IN1(n10387), .IN2(n10388), .IN3(n10351), .IN4(n10389), 
        .IN5(n10344), .QN(n10357) );
  ISOLANDX1 U23120 ( .D(n10386), .ISO(n10372), .Q(n10387) );
  AO221X1 U23121 ( .IN1(n10353), .IN2(n4038), .IN3(n2908), .IN4(n3206), .IN5(
        n10394), .Q(n10389) );
  INVX0 U23122 ( .IN(n10363), .QN(n2908) );
  AOI221X1 U23123 ( .IN1(n10077), .IN2(n10078), .IN3(n10041), .IN4(n10079), 
        .IN5(n10034), .QN(n10047) );
  ISOLANDX1 U23124 ( .D(n10076), .ISO(n10062), .Q(n10077) );
  AO221X1 U23125 ( .IN1(n10043), .IN2(n3993), .IN3(n2924), .IN4(n3210), .IN5(
        n10084), .Q(n10079) );
  INVX0 U23126 ( .IN(n10053), .QN(n2924) );
  AOI221X1 U23127 ( .IN1(n11935), .IN2(n11936), .IN3(n11899), .IN4(n11937), 
        .IN5(n11892), .QN(n11905) );
  ISOLANDX1 U23128 ( .D(n11934), .ISO(n11920), .Q(n11935) );
  AO221X1 U23129 ( .IN1(n11901), .IN2(n3588), .IN3(n3068), .IN4(n3246), .IN5(
        n11942), .Q(n11937) );
  INVX0 U23130 ( .IN(n11911), .QN(n3068) );
  AOI221X1 U23131 ( .IN1(n11625), .IN2(n11626), .IN3(n11589), .IN4(n11627), 
        .IN5(n11582), .QN(n11595) );
  ISOLANDX1 U23132 ( .D(n11624), .ISO(n11610), .Q(n11625) );
  AO221X1 U23133 ( .IN1(n11591), .IN2(n3543), .IN3(n3084), .IN4(n3250), .IN5(
        n11632), .Q(n11627) );
  INVX0 U23134 ( .IN(n11601), .QN(n3084) );
  AOI221X1 U23135 ( .IN1(n9767), .IN2(n9768), .IN3(n9731), .IN4(n9769), .IN5(
        n9724), .QN(n9737) );
  ISOLANDX1 U23136 ( .D(n9766), .ISO(n9752), .Q(n9767) );
  AO221X1 U23137 ( .IN1(n9733), .IN2(n3948), .IN3(n2940), .IN4(n3214), .IN5(
        n9774), .Q(n9769) );
  INVX0 U23138 ( .IN(n9743), .QN(n2940) );
  AOI221X1 U23139 ( .IN1(n9456), .IN2(n9457), .IN3(n9420), .IN4(n9458), .IN5(
        n9413), .QN(n9426) );
  ISOLANDX1 U23140 ( .D(n9455), .ISO(n9441), .Q(n9456) );
  AO221X1 U23141 ( .IN1(n9422), .IN2(n3903), .IN3(n2956), .IN4(n3218), .IN5(
        n9463), .Q(n9458) );
  INVX0 U23142 ( .IN(n9432), .QN(n2956) );
  NAND4X0 U23143 ( .IN1(n14064), .IN2(n14065), .IN3(n14066), .IN4(n14067), 
        .QN(n14001) );
  OA22X1 U23144 ( .IN1(n3093), .IN2(n14038), .IN3(n14037), .IN4(n2838), .Q(
        n14064) );
  OA22X1 U23145 ( .IN1(n14016), .IN2(n3254), .IN3(n14035), .IN4(n3189), .Q(
        n14065) );
  OA22X1 U23146 ( .IN1(n3462), .IN2(n14063), .IN3(n14022), .IN4(n3398), .Q(
        n14067) );
  NAND4X0 U23147 ( .IN1(n13864), .IN2(n13865), .IN3(n13866), .IN4(n13867), 
        .QN(n13804) );
  OA22X1 U23148 ( .IN1(n3144), .IN2(n13837), .IN3(n2974), .IN4(n13836), .Q(
        n13864) );
  OA22X1 U23149 ( .IN1(n3322), .IN2(n13816), .IN3(n3223), .IN4(n13834), .Q(
        n13865) );
  OA22X1 U23150 ( .IN1(n3496), .IN2(n13862), .IN3(n13850), .IN4(n3432), .Q(
        n13867) );
  NAND4X0 U23151 ( .IN1(n13733), .IN2(n13734), .IN3(n13735), .IN4(n13736), 
        .QN(n13679) );
  OA22X1 U23152 ( .IN1(n3141), .IN2(n13709), .IN3(n2966), .IN4(n13708), .Q(
        n13733) );
  OA22X1 U23153 ( .IN1(n3318), .IN2(n13691), .IN3(n3221), .IN4(n13707), .Q(
        n13734) );
  OA22X1 U23154 ( .IN1(n3494), .IN2(n13731), .IN3(n13720), .IN4(n3430), .Q(
        n13736) );
  NAND4X0 U23155 ( .IN1(n13555), .IN2(n13556), .IN3(n13557), .IN4(n13558), 
        .QN(n13495) );
  OA22X1 U23156 ( .IN1(n3150), .IN2(n13528), .IN3(n2990), .IN4(n13527), .Q(
        n13555) );
  OA22X1 U23157 ( .IN1(n3330), .IN2(n13507), .IN3(n3227), .IN4(n13525), .Q(
        n13556) );
  OA22X1 U23158 ( .IN1(n3500), .IN2(n13553), .IN3(n13541), .IN4(n3436), .Q(
        n13558) );
  NAND4X0 U23159 ( .IN1(n13424), .IN2(n13425), .IN3(n13426), .IN4(n13427), 
        .QN(n13370) );
  OA22X1 U23160 ( .IN1(n3147), .IN2(n13400), .IN3(n2982), .IN4(n13399), .Q(
        n13424) );
  OA22X1 U23161 ( .IN1(n3326), .IN2(n13382), .IN3(n3225), .IN4(n13398), .Q(
        n13425) );
  OA22X1 U23162 ( .IN1(n3498), .IN2(n13422), .IN3(n13411), .IN4(n3434), .Q(
        n13427) );
  NAND4X0 U23163 ( .IN1(n11389), .IN2(n11390), .IN3(n11391), .IN4(n11392), 
        .QN(n11329) );
  OA22X1 U23164 ( .IN1(n3102), .IN2(n11362), .IN3(n2862), .IN4(n11361), .Q(
        n11389) );
  OA22X1 U23165 ( .IN1(n3266), .IN2(n11341), .IN3(n3195), .IN4(n11359), .Q(
        n11390) );
  OA22X1 U23166 ( .IN1(n3468), .IN2(n11387), .IN3(n11375), .IN4(n3404), .Q(
        n11392) );
  NAND4X0 U23167 ( .IN1(n11258), .IN2(n11259), .IN3(n11260), .IN4(n11261), 
        .QN(n11204) );
  OA22X1 U23168 ( .IN1(n3099), .IN2(n11234), .IN3(n2854), .IN4(n11233), .Q(
        n11258) );
  OA22X1 U23169 ( .IN1(n3262), .IN2(n11216), .IN3(n3193), .IN4(n11232), .Q(
        n11259) );
  OA22X1 U23170 ( .IN1(n3466), .IN2(n11256), .IN3(n11245), .IN4(n3402), .Q(
        n11261) );
  NAND4X0 U23171 ( .IN1(n13246), .IN2(n13247), .IN3(n13248), .IN4(n13249), 
        .QN(n13186) );
  OA22X1 U23172 ( .IN1(n3156), .IN2(n13219), .IN3(n3006), .IN4(n13218), .Q(
        n13246) );
  OA22X1 U23173 ( .IN1(n3338), .IN2(n13198), .IN3(n3231), .IN4(n13216), .Q(
        n13247) );
  OA22X1 U23174 ( .IN1(n3504), .IN2(n13244), .IN3(n13232), .IN4(n3440), .Q(
        n13249) );
  NAND4X0 U23175 ( .IN1(n13115), .IN2(n13116), .IN3(n13117), .IN4(n13118), 
        .QN(n13061) );
  OA22X1 U23176 ( .IN1(n3153), .IN2(n13091), .IN3(n2998), .IN4(n13090), .Q(
        n13115) );
  OA22X1 U23177 ( .IN1(n3334), .IN2(n13073), .IN3(n3229), .IN4(n13089), .Q(
        n13116) );
  OA22X1 U23178 ( .IN1(n3502), .IN2(n13113), .IN3(n13102), .IN4(n3438), .Q(
        n13118) );
  NAND4X0 U23179 ( .IN1(n12937), .IN2(n12938), .IN3(n12939), .IN4(n12940), 
        .QN(n12877) );
  OA22X1 U23180 ( .IN1(n3162), .IN2(n12910), .IN3(n3022), .IN4(n12909), .Q(
        n12937) );
  OA22X1 U23181 ( .IN1(n3346), .IN2(n12889), .IN3(n3235), .IN4(n12907), .Q(
        n12938) );
  OA22X1 U23182 ( .IN1(n3508), .IN2(n12935), .IN3(n12923), .IN4(n3444), .Q(
        n12940) );
  NAND4X0 U23183 ( .IN1(n12806), .IN2(n12807), .IN3(n12808), .IN4(n12809), 
        .QN(n12752) );
  OA22X1 U23184 ( .IN1(n3159), .IN2(n12782), .IN3(n3014), .IN4(n12781), .Q(
        n12806) );
  OA22X1 U23185 ( .IN1(n3342), .IN2(n12764), .IN3(n3233), .IN4(n12780), .Q(
        n12807) );
  OA22X1 U23186 ( .IN1(n3506), .IN2(n12804), .IN3(n12793), .IN4(n3442), .Q(
        n12809) );
  NAND4X0 U23187 ( .IN1(n11080), .IN2(n11081), .IN3(n11082), .IN4(n11083), 
        .QN(n11020) );
  OA22X1 U23188 ( .IN1(n3108), .IN2(n11053), .IN3(n2878), .IN4(n11052), .Q(
        n11080) );
  OA22X1 U23189 ( .IN1(n3274), .IN2(n11032), .IN3(n3199), .IN4(n11050), .Q(
        n11081) );
  OA22X1 U23190 ( .IN1(n3472), .IN2(n11078), .IN3(n11066), .IN4(n3408), .Q(
        n11083) );
  NAND4X0 U23191 ( .IN1(n10949), .IN2(n10950), .IN3(n10951), .IN4(n10952), 
        .QN(n10895) );
  OA22X1 U23192 ( .IN1(n3105), .IN2(n10925), .IN3(n2870), .IN4(n10924), .Q(
        n10949) );
  OA22X1 U23193 ( .IN1(n3270), .IN2(n10907), .IN3(n3197), .IN4(n10923), .Q(
        n10950) );
  OA22X1 U23194 ( .IN1(n3470), .IN2(n10947), .IN3(n10936), .IN4(n3406), .Q(
        n10952) );
  NAND4X0 U23195 ( .IN1(n10770), .IN2(n10771), .IN3(n10772), .IN4(n10773), 
        .QN(n10710) );
  OA22X1 U23196 ( .IN1(n3114), .IN2(n10743), .IN3(n2894), .IN4(n10742), .Q(
        n10770) );
  OA22X1 U23197 ( .IN1(n3282), .IN2(n10722), .IN3(n3203), .IN4(n10740), .Q(
        n10771) );
  OA22X1 U23198 ( .IN1(n3476), .IN2(n10768), .IN3(n10756), .IN4(n3412), .Q(
        n10773) );
  NAND4X0 U23199 ( .IN1(n10639), .IN2(n10640), .IN3(n10641), .IN4(n10642), 
        .QN(n10585) );
  OA22X1 U23200 ( .IN1(n3111), .IN2(n10615), .IN3(n2886), .IN4(n10614), .Q(
        n10639) );
  OA22X1 U23201 ( .IN1(n3278), .IN2(n10597), .IN3(n3201), .IN4(n10613), .Q(
        n10640) );
  OA22X1 U23202 ( .IN1(n3474), .IN2(n10637), .IN3(n10626), .IN4(n3410), .Q(
        n10642) );
  NAND4X0 U23203 ( .IN1(n12628), .IN2(n12629), .IN3(n12630), .IN4(n12631), 
        .QN(n12568) );
  OA22X1 U23204 ( .IN1(n3168), .IN2(n12601), .IN3(n3038), .IN4(n12600), .Q(
        n12628) );
  OA22X1 U23205 ( .IN1(n3354), .IN2(n12580), .IN3(n3239), .IN4(n12598), .Q(
        n12629) );
  OA22X1 U23206 ( .IN1(n3512), .IN2(n12626), .IN3(n12614), .IN4(n3448), .Q(
        n12631) );
  NAND4X0 U23207 ( .IN1(n12497), .IN2(n12498), .IN3(n12499), .IN4(n12500), 
        .QN(n12443) );
  OA22X1 U23208 ( .IN1(n3165), .IN2(n12473), .IN3(n3030), .IN4(n12472), .Q(
        n12497) );
  OA22X1 U23209 ( .IN1(n3350), .IN2(n12455), .IN3(n3237), .IN4(n12471), .Q(
        n12498) );
  OA22X1 U23210 ( .IN1(n3510), .IN2(n12495), .IN3(n12484), .IN4(n3446), .Q(
        n12500) );
  NAND4X0 U23211 ( .IN1(n12319), .IN2(n12320), .IN3(n12321), .IN4(n12322), 
        .QN(n12259) );
  OA22X1 U23212 ( .IN1(n3174), .IN2(n12292), .IN3(n3054), .IN4(n12291), .Q(
        n12319) );
  OA22X1 U23213 ( .IN1(n3362), .IN2(n12271), .IN3(n3243), .IN4(n12289), .Q(
        n12320) );
  OA22X1 U23214 ( .IN1(n3516), .IN2(n12317), .IN3(n12305), .IN4(n3452), .Q(
        n12322) );
  NAND4X0 U23215 ( .IN1(n12188), .IN2(n12189), .IN3(n12190), .IN4(n12191), 
        .QN(n12134) );
  OA22X1 U23216 ( .IN1(n3171), .IN2(n12164), .IN3(n3046), .IN4(n12163), .Q(
        n12188) );
  OA22X1 U23217 ( .IN1(n3358), .IN2(n12146), .IN3(n3241), .IN4(n12162), .Q(
        n12189) );
  OA22X1 U23218 ( .IN1(n3514), .IN2(n12186), .IN3(n12175), .IN4(n3450), .Q(
        n12191) );
  NAND4X0 U23219 ( .IN1(n10461), .IN2(n10462), .IN3(n10463), .IN4(n10464), 
        .QN(n10401) );
  OA22X1 U23220 ( .IN1(n3120), .IN2(n10434), .IN3(n2910), .IN4(n10433), .Q(
        n10461) );
  OA22X1 U23221 ( .IN1(n3290), .IN2(n10413), .IN3(n3207), .IN4(n10431), .Q(
        n10462) );
  OA22X1 U23222 ( .IN1(n3480), .IN2(n10459), .IN3(n10447), .IN4(n3416), .Q(
        n10464) );
  NAND4X0 U23223 ( .IN1(n10330), .IN2(n10331), .IN3(n10332), .IN4(n10333), 
        .QN(n10276) );
  OA22X1 U23224 ( .IN1(n3117), .IN2(n10306), .IN3(n2902), .IN4(n10305), .Q(
        n10330) );
  OA22X1 U23225 ( .IN1(n3286), .IN2(n10288), .IN3(n3205), .IN4(n10304), .Q(
        n10331) );
  OA22X1 U23226 ( .IN1(n3478), .IN2(n10328), .IN3(n10317), .IN4(n3414), .Q(
        n10333) );
  NAND4X0 U23227 ( .IN1(n10151), .IN2(n10152), .IN3(n10153), .IN4(n10154), 
        .QN(n10091) );
  OA22X1 U23228 ( .IN1(n3126), .IN2(n10124), .IN3(n2926), .IN4(n10123), .Q(
        n10151) );
  OA22X1 U23229 ( .IN1(n3298), .IN2(n10103), .IN3(n3211), .IN4(n10121), .Q(
        n10152) );
  OA22X1 U23230 ( .IN1(n3484), .IN2(n10149), .IN3(n10137), .IN4(n3420), .Q(
        n10154) );
  NAND4X0 U23231 ( .IN1(n10020), .IN2(n10021), .IN3(n10022), .IN4(n10023), 
        .QN(n9966) );
  OA22X1 U23232 ( .IN1(n3123), .IN2(n9996), .IN3(n2918), .IN4(n9995), .Q(
        n10020) );
  OA22X1 U23233 ( .IN1(n3294), .IN2(n9978), .IN3(n3209), .IN4(n9994), .Q(
        n10021) );
  OA22X1 U23234 ( .IN1(n3482), .IN2(n10018), .IN3(n10007), .IN4(n3418), .Q(
        n10023) );
  NAND4X0 U23235 ( .IN1(n12009), .IN2(n12010), .IN3(n12011), .IN4(n12012), 
        .QN(n11949) );
  OA22X1 U23236 ( .IN1(n3180), .IN2(n11982), .IN3(n3070), .IN4(n11981), .Q(
        n12009) );
  OA22X1 U23237 ( .IN1(n3370), .IN2(n11961), .IN3(n3247), .IN4(n11979), .Q(
        n12010) );
  OA22X1 U23238 ( .IN1(n3520), .IN2(n12007), .IN3(n11995), .IN4(n3456), .Q(
        n12012) );
  NAND4X0 U23239 ( .IN1(n11878), .IN2(n11879), .IN3(n11880), .IN4(n11881), 
        .QN(n11824) );
  OA22X1 U23240 ( .IN1(n3177), .IN2(n11854), .IN3(n3062), .IN4(n11853), .Q(
        n11878) );
  OA22X1 U23241 ( .IN1(n3366), .IN2(n11836), .IN3(n3245), .IN4(n11852), .Q(
        n11879) );
  OA22X1 U23242 ( .IN1(n3518), .IN2(n11876), .IN3(n11865), .IN4(n3454), .Q(
        n11881) );
  NAND4X0 U23243 ( .IN1(n11699), .IN2(n11700), .IN3(n11701), .IN4(n11702), 
        .QN(n11639) );
  OA22X1 U23244 ( .IN1(n3186), .IN2(n11672), .IN3(n3086), .IN4(n11671), .Q(
        n11699) );
  OA22X1 U23245 ( .IN1(n3378), .IN2(n11651), .IN3(n3251), .IN4(n11669), .Q(
        n11700) );
  OA22X1 U23246 ( .IN1(n3524), .IN2(n11697), .IN3(n11685), .IN4(n3460), .Q(
        n11702) );
  NAND4X0 U23247 ( .IN1(n11568), .IN2(n11569), .IN3(n11570), .IN4(n11571), 
        .QN(n11514) );
  OA22X1 U23248 ( .IN1(n3183), .IN2(n11544), .IN3(n3078), .IN4(n11543), .Q(
        n11568) );
  OA22X1 U23249 ( .IN1(n3374), .IN2(n11526), .IN3(n3249), .IN4(n11542), .Q(
        n11569) );
  OA22X1 U23250 ( .IN1(n3522), .IN2(n11566), .IN3(n11555), .IN4(n3458), .Q(
        n11571) );
  NAND4X0 U23251 ( .IN1(n9841), .IN2(n9842), .IN3(n9843), .IN4(n9844), .QN(
        n9781) );
  OA22X1 U23252 ( .IN1(n3132), .IN2(n9814), .IN3(n2942), .IN4(n9813), .Q(n9841) );
  OA22X1 U23253 ( .IN1(n3306), .IN2(n9793), .IN3(n3215), .IN4(n9811), .Q(n9842) );
  OA22X1 U23254 ( .IN1(n3488), .IN2(n9839), .IN3(n9827), .IN4(n3424), .Q(n9844) );
  NAND4X0 U23255 ( .IN1(n9710), .IN2(n9711), .IN3(n9712), .IN4(n9713), .QN(
        n9656) );
  OA22X1 U23256 ( .IN1(n3129), .IN2(n9686), .IN3(n2934), .IN4(n9685), .Q(n9710) );
  OA22X1 U23257 ( .IN1(n3302), .IN2(n9668), .IN3(n3213), .IN4(n9684), .Q(n9711) );
  OA22X1 U23258 ( .IN1(n3486), .IN2(n9708), .IN3(n9697), .IN4(n3422), .Q(n9713) );
  NAND4X0 U23259 ( .IN1(n9530), .IN2(n9531), .IN3(n9532), .IN4(n9533), .QN(
        n9470) );
  OA22X1 U23260 ( .IN1(n3138), .IN2(n9503), .IN3(n2958), .IN4(n9502), .Q(n9530) );
  OA22X1 U23261 ( .IN1(n3314), .IN2(n9482), .IN3(n3219), .IN4(n9500), .Q(n9531) );
  OA22X1 U23262 ( .IN1(n3492), .IN2(n9528), .IN3(n9516), .IN4(n3428), .Q(n9533) );
  NAND4X0 U23263 ( .IN1(n9399), .IN2(n9400), .IN3(n9401), .IN4(n9402), .QN(
        n9345) );
  OA22X1 U23264 ( .IN1(n3135), .IN2(n9375), .IN3(n2950), .IN4(n9374), .Q(n9399) );
  OA22X1 U23265 ( .IN1(n3310), .IN2(n9357), .IN3(n3217), .IN4(n9373), .Q(n9400) );
  OA22X1 U23266 ( .IN1(n3490), .IN2(n9397), .IN3(n9386), .IN4(n3426), .Q(n9402) );
  NAND4X0 U23267 ( .IN1(n14490), .IN2(n14491), .IN3(n14492), .IN4(n14493), 
        .QN(m7_rty_o) );
  OA221X1 U23268 ( .IN1(n8847), .IN2(n2346), .IN3(n8551), .IN4(n2696), .IN5(
        n14499), .Q(n14490) );
  OA221X1 U23269 ( .IN1(n6591), .IN2(n2416), .IN3(n6295), .IN4(n2451), .IN5(
        n14495), .Q(n14492) );
  OA221X1 U23270 ( .IN1(n4815), .IN2(n2626), .IN3(n4519), .IN4(n2661), .IN5(
        n14494), .Q(n14493) );
  NAND4X0 U23271 ( .IN1(n14500), .IN2(n14501), .IN3(n14502), .IN4(n14503), 
        .QN(m7_err_o) );
  OA221X1 U23272 ( .IN1(n8847), .IN2(n2345), .IN3(n8551), .IN4(n2695), .IN5(
        n14508), .Q(n14500) );
  OA221X1 U23273 ( .IN1(n6591), .IN2(n2415), .IN3(n6295), .IN4(n2450), .IN5(
        n14505), .Q(n14502) );
  OA221X1 U23274 ( .IN1(n4815), .IN2(n2625), .IN3(n4519), .IN4(n2660), .IN5(
        n14504), .Q(n14503) );
  NAND4X0 U23275 ( .IN1(n14813), .IN2(n14814), .IN3(n14815), .IN4(n14816), 
        .QN(m7_ack_o) );
  OA221X1 U23276 ( .IN1(n8847), .IN2(n2344), .IN3(n8551), .IN4(n2694), .IN5(
        n14862), .Q(n14813) );
  OA221X1 U23277 ( .IN1(n6591), .IN2(n2414), .IN3(n6295), .IN4(n2449), .IN5(
        n14836), .Q(n14815) );
  OA221X1 U23278 ( .IN1(n4815), .IN2(n2624), .IN3(n4519), .IN4(n2659), .IN5(
        n14817), .Q(n14816) );
  NAND4X0 U23279 ( .IN1(n14804), .IN2(n14805), .IN3(n14806), .IN4(n14807), 
        .QN(m7_data_o[0]) );
  OA221X1 U23280 ( .IN1(n18776), .IN2(n2413), .IN3(n18773), .IN4(n2448), .IN5(
        n14812), .Q(n14804) );
  OA221X1 U23281 ( .IN1(n18789), .IN2(n2483), .IN3(n18785), .IN4(n2518), .IN5(
        n14811), .Q(n14805) );
  OA221X1 U23282 ( .IN1(n18800), .IN2(n2623), .IN3(n18797), .IN4(n2658), .IN5(
        n14810), .Q(n14806) );
  NAND4X0 U23283 ( .IN1(n14705), .IN2(n14706), .IN3(n14707), .IN4(n14708), 
        .QN(m7_data_o[1]) );
  OA221X1 U23284 ( .IN1(n18778), .IN2(n2412), .IN3(n18774), .IN4(n2447), .IN5(
        n14713), .Q(n14705) );
  OA221X1 U23285 ( .IN1(n18788), .IN2(n2482), .IN3(n18785), .IN4(n2517), .IN5(
        n14712), .Q(n14706) );
  OA221X1 U23286 ( .IN1(n18800), .IN2(n2622), .IN3(n18797), .IN4(n2657), .IN5(
        n14711), .Q(n14707) );
  NAND4X0 U23287 ( .IN1(n14606), .IN2(n14607), .IN3(n14608), .IN4(n14609), 
        .QN(m7_data_o[2]) );
  OA221X1 U23288 ( .IN1(n18776), .IN2(n2411), .IN3(n18773), .IN4(n2446), .IN5(
        n14614), .Q(n14606) );
  OA221X1 U23289 ( .IN1(n18788), .IN2(n2481), .IN3(n18787), .IN4(n2516), .IN5(
        n14613), .Q(n14607) );
  OA221X1 U23290 ( .IN1(n18802), .IN2(n2621), .IN3(n18798), .IN4(n2656), .IN5(
        n14612), .Q(n14608) );
  NAND4X0 U23291 ( .IN1(n14579), .IN2(n14580), .IN3(n14581), .IN4(n14582), 
        .QN(m7_data_o[3]) );
  OA221X1 U23292 ( .IN1(n18777), .IN2(n2410), .IN3(n18775), .IN4(n2445), .IN5(
        n14587), .Q(n14579) );
  OA221X1 U23293 ( .IN1(n18790), .IN2(n2480), .IN3(n18786), .IN4(n2515), .IN5(
        n14586), .Q(n14580) );
  OA221X1 U23294 ( .IN1(n18802), .IN2(n2620), .IN3(n18798), .IN4(n2655), .IN5(
        n14585), .Q(n14581) );
  NAND4X0 U23295 ( .IN1(n14570), .IN2(n14571), .IN3(n14572), .IN4(n14573), 
        .QN(m7_data_o[4]) );
  OA221X1 U23296 ( .IN1(n18777), .IN2(n2409), .IN3(n18773), .IN4(n2444), .IN5(
        n14578), .Q(n14570) );
  OA221X1 U23297 ( .IN1(n18789), .IN2(n2479), .IN3(n18786), .IN4(n2514), .IN5(
        n14577), .Q(n14571) );
  OA221X1 U23298 ( .IN1(n18801), .IN2(n2619), .IN3(n18799), .IN4(n2654), .IN5(
        n14576), .Q(n14572) );
  NAND4X0 U23299 ( .IN1(n14561), .IN2(n14562), .IN3(n14563), .IN4(n14564), 
        .QN(m7_data_o[5]) );
  OA221X1 U23300 ( .IN1(n18776), .IN2(n2408), .IN3(n18774), .IN4(n2443), .IN5(
        n14569), .Q(n14561) );
  OA221X1 U23301 ( .IN1(n18790), .IN2(n2478), .IN3(n18786), .IN4(n2513), .IN5(
        n14568), .Q(n14562) );
  OA221X1 U23302 ( .IN1(n18802), .IN2(n2618), .IN3(n18798), .IN4(n2653), .IN5(
        n14567), .Q(n14563) );
  NAND4X0 U23303 ( .IN1(n14552), .IN2(n14553), .IN3(n14554), .IN4(n14555), 
        .QN(m7_data_o[6]) );
  OA221X1 U23304 ( .IN1(n18778), .IN2(n2407), .IN3(n18775), .IN4(n2442), .IN5(
        n14560), .Q(n14552) );
  OA221X1 U23305 ( .IN1(n18790), .IN2(n2477), .IN3(n18787), .IN4(n2512), .IN5(
        n14559), .Q(n14553) );
  OA221X1 U23306 ( .IN1(n18802), .IN2(n2617), .IN3(n18799), .IN4(n2652), .IN5(
        n14558), .Q(n14554) );
  NAND4X0 U23307 ( .IN1(n14543), .IN2(n14544), .IN3(n14545), .IN4(n14546), 
        .QN(m7_data_o[7]) );
  OA221X1 U23308 ( .IN1(n18778), .IN2(n2406), .IN3(n18775), .IN4(n2441), .IN5(
        n14551), .Q(n14543) );
  OA221X1 U23309 ( .IN1(n18790), .IN2(n2476), .IN3(n18787), .IN4(n2511), .IN5(
        n14550), .Q(n14544) );
  OA221X1 U23310 ( .IN1(n18802), .IN2(n2616), .IN3(n18799), .IN4(n2651), .IN5(
        n14549), .Q(n14545) );
  NAND4X0 U23311 ( .IN1(n14534), .IN2(n14535), .IN3(n14536), .IN4(n14537), 
        .QN(m7_data_o[8]) );
  OA221X1 U23312 ( .IN1(n18778), .IN2(n2405), .IN3(n18775), .IN4(n2440), .IN5(
        n14542), .Q(n14534) );
  OA221X1 U23313 ( .IN1(n18790), .IN2(n2475), .IN3(n18787), .IN4(n2510), .IN5(
        n14541), .Q(n14535) );
  OA221X1 U23314 ( .IN1(n18802), .IN2(n2615), .IN3(n18799), .IN4(n2650), .IN5(
        n14540), .Q(n14536) );
  NAND4X0 U23315 ( .IN1(n14509), .IN2(n14510), .IN3(n14511), .IN4(n14512), 
        .QN(m7_data_o[9]) );
  OA221X1 U23316 ( .IN1(n18778), .IN2(n2404), .IN3(n18775), .IN4(n2439), .IN5(
        n14531), .Q(n14509) );
  OA221X1 U23317 ( .IN1(n18790), .IN2(n2474), .IN3(n18787), .IN4(n2509), .IN5(
        n14526), .Q(n14510) );
  OA221X1 U23318 ( .IN1(n18802), .IN2(n2614), .IN3(n18799), .IN4(n2649), .IN5(
        n14521), .Q(n14511) );
  NAND4X0 U23319 ( .IN1(n14795), .IN2(n14796), .IN3(n14797), .IN4(n14798), 
        .QN(m7_data_o[10]) );
  OA221X1 U23320 ( .IN1(n18778), .IN2(n2403), .IN3(n18773), .IN4(n2438), .IN5(
        n14803), .Q(n14795) );
  OA221X1 U23321 ( .IN1(n18790), .IN2(n2473), .IN3(n18785), .IN4(n2508), .IN5(
        n14802), .Q(n14796) );
  OA221X1 U23322 ( .IN1(n18800), .IN2(n2613), .IN3(n18797), .IN4(n2648), .IN5(
        n14801), .Q(n14797) );
  NAND4X0 U23323 ( .IN1(n14786), .IN2(n14787), .IN3(n14788), .IN4(n14789), 
        .QN(m7_data_o[11]) );
  OA221X1 U23324 ( .IN1(n18777), .IN2(n2402), .IN3(n18773), .IN4(n2437), .IN5(
        n14794), .Q(n14786) );
  OA221X1 U23325 ( .IN1(n18788), .IN2(n2472), .IN3(n18785), .IN4(n2507), .IN5(
        n14793), .Q(n14787) );
  OA221X1 U23326 ( .IN1(n18800), .IN2(n2612), .IN3(n18797), .IN4(n2647), .IN5(
        n14792), .Q(n14788) );
  NAND4X0 U23327 ( .IN1(n14777), .IN2(n14778), .IN3(n14779), .IN4(n14780), 
        .QN(m7_data_o[12]) );
  OA221X1 U23328 ( .IN1(n18776), .IN2(n2401), .IN3(n18773), .IN4(n2436), .IN5(
        n14785), .Q(n14777) );
  OA221X1 U23329 ( .IN1(n18789), .IN2(n2471), .IN3(n18785), .IN4(n2506), .IN5(
        n14784), .Q(n14778) );
  OA221X1 U23330 ( .IN1(n18800), .IN2(n2611), .IN3(n18797), .IN4(n2646), .IN5(
        n14783), .Q(n14779) );
  NAND4X0 U23331 ( .IN1(n14768), .IN2(n14769), .IN3(n14770), .IN4(n14771), 
        .QN(m7_data_o[13]) );
  OA221X1 U23332 ( .IN1(n18776), .IN2(n2400), .IN3(n18774), .IN4(n2435), .IN5(
        n14776), .Q(n14768) );
  OA221X1 U23333 ( .IN1(n18790), .IN2(n2470), .IN3(n18787), .IN4(n2505), .IN5(
        n14775), .Q(n14769) );
  OA221X1 U23334 ( .IN1(n18800), .IN2(n2610), .IN3(n18799), .IN4(n2645), .IN5(
        n14774), .Q(n14770) );
  NAND4X0 U23335 ( .IN1(n14759), .IN2(n14760), .IN3(n14761), .IN4(n14762), 
        .QN(m7_data_o[14]) );
  OA221X1 U23336 ( .IN1(n18778), .IN2(n2399), .IN3(n18774), .IN4(n2434), .IN5(
        n14767), .Q(n14759) );
  OA221X1 U23337 ( .IN1(n18788), .IN2(n2469), .IN3(n18785), .IN4(n2504), .IN5(
        n14766), .Q(n14760) );
  OA221X1 U23338 ( .IN1(n18800), .IN2(n2609), .IN3(n18797), .IN4(n2644), .IN5(
        n14765), .Q(n14761) );
  NAND4X0 U23339 ( .IN1(n14750), .IN2(n14751), .IN3(n14752), .IN4(n14753), 
        .QN(m7_data_o[15]) );
  OA221X1 U23340 ( .IN1(n18777), .IN2(n2398), .IN3(n18774), .IN4(n2433), .IN5(
        n14758), .Q(n14750) );
  OA221X1 U23341 ( .IN1(n18788), .IN2(n2468), .IN3(n18786), .IN4(n2503), .IN5(
        n14757), .Q(n14751) );
  OA221X1 U23342 ( .IN1(n18800), .IN2(n2608), .IN3(n18798), .IN4(n2643), .IN5(
        n14756), .Q(n14752) );
  NAND4X0 U23343 ( .IN1(n14741), .IN2(n14742), .IN3(n14743), .IN4(n14744), 
        .QN(m7_data_o[16]) );
  OA221X1 U23344 ( .IN1(n18776), .IN2(n2397), .IN3(n18774), .IN4(n2432), .IN5(
        n14749), .Q(n14741) );
  OA221X1 U23345 ( .IN1(n18789), .IN2(n2467), .IN3(n18786), .IN4(n2502), .IN5(
        n14748), .Q(n14742) );
  OA221X1 U23346 ( .IN1(n18801), .IN2(n2607), .IN3(n18798), .IN4(n2642), .IN5(
        n14747), .Q(n14743) );
  NAND4X0 U23347 ( .IN1(n14732), .IN2(n14733), .IN3(n14734), .IN4(n14735), 
        .QN(m7_data_o[17]) );
  OA221X1 U23348 ( .IN1(n18777), .IN2(n2396), .IN3(n18775), .IN4(n2431), .IN5(
        n14740), .Q(n14732) );
  OA221X1 U23349 ( .IN1(n18790), .IN2(n2466), .IN3(n18787), .IN4(n2501), .IN5(
        n14739), .Q(n14733) );
  OA221X1 U23350 ( .IN1(n18802), .IN2(n2606), .IN3(n18799), .IN4(n2641), .IN5(
        n14738), .Q(n14734) );
  NAND4X0 U23351 ( .IN1(n14723), .IN2(n14724), .IN3(n14725), .IN4(n14726), 
        .QN(m7_data_o[18]) );
  OA221X1 U23352 ( .IN1(n18777), .IN2(n2395), .IN3(n18773), .IN4(n2430), .IN5(
        n14731), .Q(n14723) );
  OA221X1 U23353 ( .IN1(n18789), .IN2(n2465), .IN3(n18785), .IN4(n2500), .IN5(
        n14730), .Q(n14724) );
  OA221X1 U23354 ( .IN1(n18800), .IN2(n2605), .IN3(n18797), .IN4(n2640), .IN5(
        n14729), .Q(n14725) );
  NAND4X0 U23355 ( .IN1(n14714), .IN2(n14715), .IN3(n14716), .IN4(n14717), 
        .QN(m7_data_o[19]) );
  OA221X1 U23356 ( .IN1(n18778), .IN2(n2394), .IN3(n18774), .IN4(n2429), .IN5(
        n14722), .Q(n14714) );
  OA221X1 U23357 ( .IN1(n18788), .IN2(n2464), .IN3(n18785), .IN4(n2499), .IN5(
        n14721), .Q(n14715) );
  OA221X1 U23358 ( .IN1(n18801), .IN2(n2604), .IN3(n18797), .IN4(n2639), .IN5(
        n14720), .Q(n14716) );
  NAND4X0 U23359 ( .IN1(n14696), .IN2(n14697), .IN3(n14698), .IN4(n14699), 
        .QN(m7_data_o[20]) );
  OA221X1 U23360 ( .IN1(n18776), .IN2(n2393), .IN3(n18773), .IN4(n2428), .IN5(
        n14704), .Q(n14696) );
  OA221X1 U23361 ( .IN1(n18788), .IN2(n2463), .IN3(n18786), .IN4(n2498), .IN5(
        n14703), .Q(n14697) );
  OA221X1 U23362 ( .IN1(n18801), .IN2(n2603), .IN3(n18798), .IN4(n2638), .IN5(
        n14702), .Q(n14698) );
  NAND4X0 U23363 ( .IN1(n14687), .IN2(n14688), .IN3(n14689), .IN4(n14690), 
        .QN(m7_data_o[21]) );
  OA221X1 U23364 ( .IN1(n18776), .IN2(n2392), .IN3(n18774), .IN4(n2427), .IN5(
        n14695), .Q(n14687) );
  OA221X1 U23365 ( .IN1(n18788), .IN2(n2462), .IN3(n18786), .IN4(n2497), .IN5(
        n14694), .Q(n14688) );
  OA221X1 U23366 ( .IN1(n18801), .IN2(n2602), .IN3(n18798), .IN4(n2637), .IN5(
        n14693), .Q(n14689) );
  NAND4X0 U23367 ( .IN1(n14678), .IN2(n14679), .IN3(n14680), .IN4(n14681), 
        .QN(m7_data_o[22]) );
  OA221X1 U23368 ( .IN1(n18776), .IN2(n2391), .IN3(n18775), .IN4(n2426), .IN5(
        n14686), .Q(n14678) );
  OA221X1 U23369 ( .IN1(n18788), .IN2(n2461), .IN3(n18786), .IN4(n2496), .IN5(
        n14685), .Q(n14679) );
  OA221X1 U23370 ( .IN1(n18801), .IN2(n2601), .IN3(n18798), .IN4(n2636), .IN5(
        n14684), .Q(n14680) );
  NAND4X0 U23371 ( .IN1(n14669), .IN2(n14670), .IN3(n14671), .IN4(n14672), 
        .QN(m7_data_o[23]) );
  OA221X1 U23372 ( .IN1(n18776), .IN2(n2390), .IN3(n18773), .IN4(n2425), .IN5(
        n14677), .Q(n14669) );
  OA221X1 U23373 ( .IN1(n18788), .IN2(n2460), .IN3(n18786), .IN4(n2495), .IN5(
        n14676), .Q(n14670) );
  OA221X1 U23374 ( .IN1(n18801), .IN2(n2600), .IN3(n18798), .IN4(n2635), .IN5(
        n14675), .Q(n14671) );
  NAND4X0 U23375 ( .IN1(n14660), .IN2(n14661), .IN3(n14662), .IN4(n14663), 
        .QN(m7_data_o[24]) );
  OA221X1 U23376 ( .IN1(n18777), .IN2(n2389), .IN3(n18775), .IN4(n2424), .IN5(
        n14668), .Q(n14660) );
  OA221X1 U23377 ( .IN1(n18789), .IN2(n2459), .IN3(n18787), .IN4(n2494), .IN5(
        n14667), .Q(n14661) );
  OA221X1 U23378 ( .IN1(n18800), .IN2(n2599), .IN3(n18799), .IN4(n2634), .IN5(
        n14666), .Q(n14662) );
  NAND4X0 U23379 ( .IN1(n14651), .IN2(n14652), .IN3(n14653), .IN4(n14654), 
        .QN(m7_data_o[25]) );
  OA221X1 U23380 ( .IN1(n18777), .IN2(n2388), .IN3(n18775), .IN4(n2423), .IN5(
        n14659), .Q(n14651) );
  OA221X1 U23381 ( .IN1(n18789), .IN2(n2458), .IN3(n18785), .IN4(n2493), .IN5(
        n14658), .Q(n14652) );
  OA221X1 U23382 ( .IN1(n18802), .IN2(n2598), .IN3(n18797), .IN4(n2633), .IN5(
        n14657), .Q(n14653) );
  NAND4X0 U23383 ( .IN1(n14642), .IN2(n14643), .IN3(n14644), .IN4(n14645), 
        .QN(m7_data_o[26]) );
  OA221X1 U23384 ( .IN1(n18777), .IN2(n2387), .IN3(n18773), .IN4(n2422), .IN5(
        n14650), .Q(n14642) );
  OA221X1 U23385 ( .IN1(n18789), .IN2(n2457), .IN3(n18786), .IN4(n2492), .IN5(
        n14649), .Q(n14643) );
  OA221X1 U23386 ( .IN1(n18801), .IN2(n2597), .IN3(n18798), .IN4(n2632), .IN5(
        n14648), .Q(n14644) );
  NAND4X0 U23387 ( .IN1(n14633), .IN2(n14634), .IN3(n14635), .IN4(n14636), 
        .QN(m7_data_o[27]) );
  OA221X1 U23388 ( .IN1(n18777), .IN2(n2386), .IN3(n18774), .IN4(n2421), .IN5(
        n14641), .Q(n14633) );
  OA221X1 U23389 ( .IN1(n18789), .IN2(n2456), .IN3(n18787), .IN4(n2491), .IN5(
        n14640), .Q(n14634) );
  OA221X1 U23390 ( .IN1(n18802), .IN2(n2596), .IN3(n18799), .IN4(n2631), .IN5(
        n14639), .Q(n14635) );
  NAND4X0 U23391 ( .IN1(n14624), .IN2(n14625), .IN3(n14626), .IN4(n14627), 
        .QN(m7_data_o[28]) );
  OA221X1 U23392 ( .IN1(n18778), .IN2(n2385), .IN3(n18774), .IN4(n2420), .IN5(
        n14632), .Q(n14624) );
  OA221X1 U23393 ( .IN1(n18789), .IN2(n2455), .IN3(n18787), .IN4(n2490), .IN5(
        n14631), .Q(n14625) );
  OA221X1 U23394 ( .IN1(n18801), .IN2(n2595), .IN3(n18799), .IN4(n2630), .IN5(
        n14630), .Q(n14626) );
  NAND4X0 U23395 ( .IN1(n14615), .IN2(n14616), .IN3(n14617), .IN4(n14618), 
        .QN(m7_data_o[29]) );
  OA221X1 U23396 ( .IN1(n18777), .IN2(n2384), .IN3(n18775), .IN4(n2419), .IN5(
        n14623), .Q(n14615) );
  OA221X1 U23397 ( .IN1(n18789), .IN2(n2454), .IN3(n18786), .IN4(n2489), .IN5(
        n14622), .Q(n14616) );
  OA221X1 U23398 ( .IN1(n18801), .IN2(n2594), .IN3(n18797), .IN4(n2629), .IN5(
        n14621), .Q(n14617) );
  NAND4X0 U23399 ( .IN1(n14597), .IN2(n14598), .IN3(n14599), .IN4(n14600), 
        .QN(m7_data_o[30]) );
  OA221X1 U23400 ( .IN1(n18776), .IN2(n2383), .IN3(n18773), .IN4(n2418), .IN5(
        n14605), .Q(n14597) );
  OA221X1 U23401 ( .IN1(n18790), .IN2(n2453), .IN3(n18785), .IN4(n2488), .IN5(
        n14604), .Q(n14598) );
  OA221X1 U23402 ( .IN1(n18802), .IN2(n2593), .IN3(n18798), .IN4(n2628), .IN5(
        n14603), .Q(n14599) );
  NAND4X0 U23403 ( .IN1(n14588), .IN2(n14589), .IN3(n14590), .IN4(n14591), 
        .QN(m7_data_o[31]) );
  OA221X1 U23404 ( .IN1(n18778), .IN2(n2382), .IN3(n18775), .IN4(n2417), .IN5(
        n14596), .Q(n14588) );
  OA221X1 U23405 ( .IN1(n18788), .IN2(n2452), .IN3(n18787), .IN4(n2487), .IN5(
        n14595), .Q(n14589) );
  OA221X1 U23406 ( .IN1(n18801), .IN2(n2592), .IN3(n18799), .IN4(n2627), .IN5(
        n14594), .Q(n14590) );
  NAND4X0 U23407 ( .IN1(n14875), .IN2(n14876), .IN3(n14877), .IN4(n14878), 
        .QN(m6_rty_o) );
  OA221X1 U23408 ( .IN1(n8848), .IN2(n2346), .IN3(n8552), .IN4(n2696), .IN5(
        n14883), .Q(n14875) );
  OA221X1 U23409 ( .IN1(n6592), .IN2(n2416), .IN3(n6296), .IN4(n2451), .IN5(
        n14880), .Q(n14877) );
  OA221X1 U23410 ( .IN1(n4816), .IN2(n2626), .IN3(n4520), .IN4(n2661), .IN5(
        n14879), .Q(n14878) );
  NAND4X0 U23411 ( .IN1(n14884), .IN2(n14885), .IN3(n14886), .IN4(n14887), 
        .QN(m6_err_o) );
  OA221X1 U23412 ( .IN1(n8848), .IN2(n2345), .IN3(n8552), .IN4(n2695), .IN5(
        n14891), .Q(n14884) );
  OA221X1 U23413 ( .IN1(n6592), .IN2(n2415), .IN3(n6296), .IN4(n2450), .IN5(
        n14889), .Q(n14886) );
  OA221X1 U23414 ( .IN1(n4816), .IN2(n2625), .IN3(n4520), .IN4(n2660), .IN5(
        n14888), .Q(n14887) );
  NAND4X0 U23415 ( .IN1(n15164), .IN2(n15165), .IN3(n15166), .IN4(n15167), 
        .QN(m6_ack_o) );
  OA221X1 U23416 ( .IN1(n8848), .IN2(n2344), .IN3(n8552), .IN4(n2694), .IN5(
        n15179), .Q(n15164) );
  OA221X1 U23417 ( .IN1(n6592), .IN2(n2414), .IN3(n6296), .IN4(n2449), .IN5(
        n15175), .Q(n15166) );
  OA221X1 U23418 ( .IN1(n4816), .IN2(n2624), .IN3(n4520), .IN4(n2659), .IN5(
        n15168), .Q(n15167) );
  NAND4X0 U23419 ( .IN1(n15156), .IN2(n15157), .IN3(n15158), .IN4(n15159), 
        .QN(m6_data_o[0]) );
  OA221X1 U23420 ( .IN1(n18728), .IN2(n2413), .IN3(n14912), .IN4(n2448), .IN5(
        n15163), .Q(n15156) );
  OA221X1 U23421 ( .IN1(n18740), .IN2(n2483), .IN3(n18737), .IN4(n2518), .IN5(
        n15162), .Q(n15157) );
  OA221X1 U23422 ( .IN1(n18752), .IN2(n2623), .IN3(n18749), .IN4(n2658), .IN5(
        n15161), .Q(n15158) );
  NAND4X0 U23423 ( .IN1(n15068), .IN2(n15069), .IN3(n15070), .IN4(n15071), 
        .QN(m6_data_o[1]) );
  OA221X1 U23424 ( .IN1(n18730), .IN2(n2412), .IN3(n18726), .IN4(n2447), .IN5(
        n15075), .Q(n15068) );
  OA221X1 U23425 ( .IN1(n18742), .IN2(n2482), .IN3(n18737), .IN4(n2517), .IN5(
        n15074), .Q(n15069) );
  OA221X1 U23426 ( .IN1(n18754), .IN2(n2622), .IN3(n18749), .IN4(n2657), .IN5(
        n15073), .Q(n15070) );
  NAND4X0 U23427 ( .IN1(n14980), .IN2(n14981), .IN3(n14982), .IN4(n14983), 
        .QN(m6_data_o[2]) );
  OA221X1 U23428 ( .IN1(n18728), .IN2(n2411), .IN3(n18726), .IN4(n2446), .IN5(
        n14987), .Q(n14980) );
  OA221X1 U23429 ( .IN1(n18742), .IN2(n2481), .IN3(n18739), .IN4(n2516), .IN5(
        n14986), .Q(n14981) );
  OA221X1 U23430 ( .IN1(n18754), .IN2(n2621), .IN3(n18751), .IN4(n2656), .IN5(
        n14985), .Q(n14982) );
  NAND4X0 U23431 ( .IN1(n14956), .IN2(n14957), .IN3(n14958), .IN4(n14959), 
        .QN(m6_data_o[3]) );
  OA221X1 U23432 ( .IN1(n18730), .IN2(n2410), .IN3(n18726), .IN4(n2445), .IN5(
        n14963), .Q(n14956) );
  OA221X1 U23433 ( .IN1(n18742), .IN2(n2480), .IN3(n18738), .IN4(n2515), .IN5(
        n14962), .Q(n14957) );
  OA221X1 U23434 ( .IN1(n18754), .IN2(n2620), .IN3(n18750), .IN4(n2655), .IN5(
        n14961), .Q(n14958) );
  NAND4X0 U23435 ( .IN1(n14948), .IN2(n14949), .IN3(n14950), .IN4(n14951), 
        .QN(m6_data_o[4]) );
  OA221X1 U23436 ( .IN1(n18728), .IN2(n2409), .IN3(n18725), .IN4(n2444), .IN5(
        n14955), .Q(n14948) );
  OA221X1 U23437 ( .IN1(n18740), .IN2(n2479), .IN3(n18739), .IN4(n2514), .IN5(
        n14954), .Q(n14949) );
  OA221X1 U23438 ( .IN1(n18752), .IN2(n2619), .IN3(n18751), .IN4(n2654), .IN5(
        n14953), .Q(n14950) );
  NAND4X0 U23439 ( .IN1(n14940), .IN2(n14941), .IN3(n14942), .IN4(n14943), 
        .QN(m6_data_o[5]) );
  OA221X1 U23440 ( .IN1(n18729), .IN2(n2408), .IN3(n14912), .IN4(n2443), .IN5(
        n14947), .Q(n14940) );
  OA221X1 U23441 ( .IN1(n18741), .IN2(n2478), .IN3(n18739), .IN4(n2513), .IN5(
        n14946), .Q(n14941) );
  OA221X1 U23442 ( .IN1(n18753), .IN2(n2618), .IN3(n18751), .IN4(n2653), .IN5(
        n14945), .Q(n14942) );
  NAND4X0 U23443 ( .IN1(n14932), .IN2(n14933), .IN3(n14934), .IN4(n14935), 
        .QN(m6_data_o[6]) );
  OA221X1 U23444 ( .IN1(n18730), .IN2(n2407), .IN3(n18726), .IN4(n2442), .IN5(
        n14939), .Q(n14932) );
  OA221X1 U23445 ( .IN1(n18742), .IN2(n2477), .IN3(n18739), .IN4(n2512), .IN5(
        n14938), .Q(n14933) );
  OA221X1 U23446 ( .IN1(n18754), .IN2(n2617), .IN3(n18751), .IN4(n2652), .IN5(
        n14937), .Q(n14934) );
  NAND4X0 U23447 ( .IN1(n14924), .IN2(n14925), .IN3(n14926), .IN4(n14927), 
        .QN(m6_data_o[7]) );
  OA221X1 U23448 ( .IN1(n18730), .IN2(n2406), .IN3(n18726), .IN4(n2441), .IN5(
        n14931), .Q(n14924) );
  OA221X1 U23449 ( .IN1(n18742), .IN2(n2476), .IN3(n18739), .IN4(n2511), .IN5(
        n14930), .Q(n14925) );
  OA221X1 U23450 ( .IN1(n18754), .IN2(n2616), .IN3(n18751), .IN4(n2651), .IN5(
        n14929), .Q(n14926) );
  NAND4X0 U23451 ( .IN1(n14916), .IN2(n14917), .IN3(n14918), .IN4(n14919), 
        .QN(m6_data_o[8]) );
  OA221X1 U23452 ( .IN1(n18730), .IN2(n2405), .IN3(n18726), .IN4(n2440), .IN5(
        n14923), .Q(n14916) );
  OA221X1 U23453 ( .IN1(n18742), .IN2(n2475), .IN3(n18739), .IN4(n2510), .IN5(
        n14922), .Q(n14917) );
  OA221X1 U23454 ( .IN1(n18754), .IN2(n2615), .IN3(n18751), .IN4(n2650), .IN5(
        n14921), .Q(n14918) );
  NAND4X0 U23455 ( .IN1(n14892), .IN2(n14893), .IN3(n14894), .IN4(n14895), 
        .QN(m6_data_o[9]) );
  OA221X1 U23456 ( .IN1(n18730), .IN2(n2404), .IN3(n18726), .IN4(n2439), .IN5(
        n14913), .Q(n14892) );
  OA221X1 U23457 ( .IN1(n18742), .IN2(n2474), .IN3(n18739), .IN4(n2509), .IN5(
        n14908), .Q(n14893) );
  OA221X1 U23458 ( .IN1(n18754), .IN2(n2614), .IN3(n18751), .IN4(n2649), .IN5(
        n14903), .Q(n14894) );
  NAND4X0 U23459 ( .IN1(n15148), .IN2(n15149), .IN3(n15150), .IN4(n15151), 
        .QN(m6_data_o[10]) );
  OA221X1 U23460 ( .IN1(n18729), .IN2(n2403), .IN3(n14912), .IN4(n2438), .IN5(
        n15155), .Q(n15148) );
  OA221X1 U23461 ( .IN1(n18742), .IN2(n2473), .IN3(n18737), .IN4(n2508), .IN5(
        n15154), .Q(n15149) );
  OA221X1 U23462 ( .IN1(n18754), .IN2(n2613), .IN3(n18749), .IN4(n2648), .IN5(
        n15153), .Q(n15150) );
  NAND4X0 U23463 ( .IN1(n15140), .IN2(n15141), .IN3(n15142), .IN4(n15143), 
        .QN(m6_data_o[11]) );
  OA221X1 U23464 ( .IN1(n18728), .IN2(n2402), .IN3(n14912), .IN4(n2437), .IN5(
        n15147), .Q(n15140) );
  OA221X1 U23465 ( .IN1(n18740), .IN2(n2472), .IN3(n18737), .IN4(n2507), .IN5(
        n15146), .Q(n15141) );
  OA221X1 U23466 ( .IN1(n18752), .IN2(n2612), .IN3(n18749), .IN4(n2647), .IN5(
        n15145), .Q(n15142) );
  NAND4X0 U23467 ( .IN1(n15132), .IN2(n15133), .IN3(n15134), .IN4(n15135), 
        .QN(m6_data_o[12]) );
  OA221X1 U23468 ( .IN1(n18729), .IN2(n2401), .IN3(n14912), .IN4(n2436), .IN5(
        n15139), .Q(n15132) );
  OA221X1 U23469 ( .IN1(n18741), .IN2(n2471), .IN3(n18737), .IN4(n2506), .IN5(
        n15138), .Q(n15133) );
  OA221X1 U23470 ( .IN1(n18753), .IN2(n2611), .IN3(n18749), .IN4(n2646), .IN5(
        n15137), .Q(n15134) );
  NAND4X0 U23471 ( .IN1(n15124), .IN2(n15125), .IN3(n15126), .IN4(n15127), 
        .QN(m6_data_o[13]) );
  OA221X1 U23472 ( .IN1(n18728), .IN2(n2400), .IN3(n18725), .IN4(n2435), .IN5(
        n15131), .Q(n15124) );
  OA221X1 U23473 ( .IN1(n18740), .IN2(n2470), .IN3(n18738), .IN4(n2505), .IN5(
        n15130), .Q(n15125) );
  OA221X1 U23474 ( .IN1(n18752), .IN2(n2610), .IN3(n18750), .IN4(n2645), .IN5(
        n15129), .Q(n15126) );
  NAND4X0 U23475 ( .IN1(n15116), .IN2(n15117), .IN3(n15118), .IN4(n15119), 
        .QN(m6_data_o[14]) );
  OA221X1 U23476 ( .IN1(n18728), .IN2(n2399), .IN3(n18725), .IN4(n2434), .IN5(
        n15123), .Q(n15116) );
  OA221X1 U23477 ( .IN1(n18740), .IN2(n2469), .IN3(n18738), .IN4(n2504), .IN5(
        n15122), .Q(n15117) );
  OA221X1 U23478 ( .IN1(n18752), .IN2(n2609), .IN3(n18750), .IN4(n2644), .IN5(
        n15121), .Q(n15118) );
  NAND4X0 U23479 ( .IN1(n15108), .IN2(n15109), .IN3(n15110), .IN4(n15111), 
        .QN(m6_data_o[15]) );
  OA221X1 U23480 ( .IN1(n18728), .IN2(n2398), .IN3(n18725), .IN4(n2433), .IN5(
        n15115), .Q(n15108) );
  OA221X1 U23481 ( .IN1(n18740), .IN2(n2468), .IN3(n18738), .IN4(n2503), .IN5(
        n15114), .Q(n15109) );
  OA221X1 U23482 ( .IN1(n18752), .IN2(n2608), .IN3(n18750), .IN4(n2643), .IN5(
        n15113), .Q(n15110) );
  NAND4X0 U23483 ( .IN1(n15100), .IN2(n15101), .IN3(n15102), .IN4(n15103), 
        .QN(m6_data_o[16]) );
  OA221X1 U23484 ( .IN1(n18728), .IN2(n2397), .IN3(n18725), .IN4(n2432), .IN5(
        n15107), .Q(n15100) );
  OA221X1 U23485 ( .IN1(n18740), .IN2(n2467), .IN3(n18738), .IN4(n2502), .IN5(
        n15106), .Q(n15101) );
  OA221X1 U23486 ( .IN1(n18752), .IN2(n2607), .IN3(n18750), .IN4(n2642), .IN5(
        n15105), .Q(n15102) );
  NAND4X0 U23487 ( .IN1(n15092), .IN2(n15093), .IN3(n15094), .IN4(n15095), 
        .QN(m6_data_o[17]) );
  OA221X1 U23488 ( .IN1(n18729), .IN2(n2396), .IN3(n18725), .IN4(n2431), .IN5(
        n15099), .Q(n15092) );
  OA221X1 U23489 ( .IN1(n18741), .IN2(n2466), .IN3(n18738), .IN4(n2501), .IN5(
        n15098), .Q(n15093) );
  OA221X1 U23490 ( .IN1(n18753), .IN2(n2606), .IN3(n18750), .IN4(n2641), .IN5(
        n15097), .Q(n15094) );
  NAND4X0 U23491 ( .IN1(n15084), .IN2(n15085), .IN3(n15086), .IN4(n15087), 
        .QN(m6_data_o[18]) );
  OA221X1 U23492 ( .IN1(n18729), .IN2(n2395), .IN3(n18726), .IN4(n2430), .IN5(
        n15091), .Q(n15084) );
  OA221X1 U23493 ( .IN1(n18741), .IN2(n2465), .IN3(n18739), .IN4(n2500), .IN5(
        n15090), .Q(n15085) );
  OA221X1 U23494 ( .IN1(n18753), .IN2(n2605), .IN3(n18751), .IN4(n2640), .IN5(
        n15089), .Q(n15086) );
  NAND4X0 U23495 ( .IN1(n15076), .IN2(n15077), .IN3(n15078), .IN4(n15079), 
        .QN(m6_data_o[19]) );
  OA221X1 U23496 ( .IN1(n18728), .IN2(n2394), .IN3(n18726), .IN4(n2429), .IN5(
        n15083), .Q(n15076) );
  OA221X1 U23497 ( .IN1(n18740), .IN2(n2464), .IN3(n18737), .IN4(n2499), .IN5(
        n15082), .Q(n15077) );
  OA221X1 U23498 ( .IN1(n18752), .IN2(n2604), .IN3(n18749), .IN4(n2639), .IN5(
        n15081), .Q(n15078) );
  NAND4X0 U23499 ( .IN1(n15060), .IN2(n15061), .IN3(n15062), .IN4(n15063), 
        .QN(m6_data_o[20]) );
  OA221X1 U23500 ( .IN1(n18729), .IN2(n2393), .IN3(n14912), .IN4(n2428), .IN5(
        n15067), .Q(n15060) );
  OA221X1 U23501 ( .IN1(n18741), .IN2(n2463), .IN3(n18737), .IN4(n2498), .IN5(
        n15066), .Q(n15061) );
  OA221X1 U23502 ( .IN1(n18753), .IN2(n2603), .IN3(n18749), .IN4(n2638), .IN5(
        n15065), .Q(n15062) );
  NAND4X0 U23503 ( .IN1(n15052), .IN2(n15053), .IN3(n15054), .IN4(n15055), 
        .QN(m6_data_o[21]) );
  OA221X1 U23504 ( .IN1(n18729), .IN2(n2392), .IN3(n14912), .IN4(n2427), .IN5(
        n15059), .Q(n15052) );
  OA221X1 U23505 ( .IN1(n18741), .IN2(n2462), .IN3(n18738), .IN4(n2497), .IN5(
        n15058), .Q(n15053) );
  OA221X1 U23506 ( .IN1(n18753), .IN2(n2602), .IN3(n18750), .IN4(n2637), .IN5(
        n15057), .Q(n15054) );
  NAND4X0 U23507 ( .IN1(n15044), .IN2(n15045), .IN3(n15046), .IN4(n15047), 
        .QN(m6_data_o[22]) );
  OA221X1 U23508 ( .IN1(n18729), .IN2(n2391), .IN3(n14912), .IN4(n2426), .IN5(
        n15051), .Q(n15044) );
  OA221X1 U23509 ( .IN1(n18741), .IN2(n2461), .IN3(n18739), .IN4(n2496), .IN5(
        n15050), .Q(n15045) );
  OA221X1 U23510 ( .IN1(n18753), .IN2(n2601), .IN3(n18751), .IN4(n2636), .IN5(
        n15049), .Q(n15046) );
  NAND4X0 U23511 ( .IN1(n15036), .IN2(n15037), .IN3(n15038), .IN4(n15039), 
        .QN(m6_data_o[23]) );
  OA221X1 U23512 ( .IN1(n18729), .IN2(n2390), .IN3(n14912), .IN4(n2425), .IN5(
        n15043), .Q(n15036) );
  OA221X1 U23513 ( .IN1(n18741), .IN2(n2460), .IN3(n18737), .IN4(n2495), .IN5(
        n15042), .Q(n15037) );
  OA221X1 U23514 ( .IN1(n18753), .IN2(n2600), .IN3(n18749), .IN4(n2635), .IN5(
        n15041), .Q(n15038) );
  NAND4X0 U23515 ( .IN1(n15028), .IN2(n15029), .IN3(n15030), .IN4(n15031), 
        .QN(m6_data_o[24]) );
  OA221X1 U23516 ( .IN1(n18729), .IN2(n2389), .IN3(n18725), .IN4(n2424), .IN5(
        n15035), .Q(n15028) );
  OA221X1 U23517 ( .IN1(n18741), .IN2(n2459), .IN3(n18737), .IN4(n2494), .IN5(
        n15034), .Q(n15029) );
  OA221X1 U23518 ( .IN1(n18753), .IN2(n2599), .IN3(n18749), .IN4(n2634), .IN5(
        n15033), .Q(n15030) );
  NAND4X0 U23519 ( .IN1(n15020), .IN2(n15021), .IN3(n15022), .IN4(n15023), 
        .QN(m6_data_o[25]) );
  OA221X1 U23520 ( .IN1(n18730), .IN2(n2388), .IN3(n18725), .IN4(n2423), .IN5(
        n15027), .Q(n15020) );
  OA221X1 U23521 ( .IN1(n18742), .IN2(n2458), .IN3(n18738), .IN4(n2493), .IN5(
        n15026), .Q(n15021) );
  OA221X1 U23522 ( .IN1(n18754), .IN2(n2598), .IN3(n18750), .IN4(n2633), .IN5(
        n15025), .Q(n15022) );
  NAND4X0 U23523 ( .IN1(n15012), .IN2(n15013), .IN3(n15014), .IN4(n15015), 
        .QN(m6_data_o[26]) );
  OA221X1 U23524 ( .IN1(n18729), .IN2(n2387), .IN3(n14912), .IN4(n2422), .IN5(
        n15019), .Q(n15012) );
  OA221X1 U23525 ( .IN1(n18741), .IN2(n2457), .IN3(n18739), .IN4(n2492), .IN5(
        n15018), .Q(n15013) );
  OA221X1 U23526 ( .IN1(n18753), .IN2(n2597), .IN3(n18751), .IN4(n2632), .IN5(
        n15017), .Q(n15014) );
  NAND4X0 U23527 ( .IN1(n15004), .IN2(n15005), .IN3(n15006), .IN4(n15007), 
        .QN(m6_data_o[27]) );
  OA221X1 U23528 ( .IN1(n18728), .IN2(n2386), .IN3(n14912), .IN4(n2421), .IN5(
        n15011), .Q(n15004) );
  OA221X1 U23529 ( .IN1(n18740), .IN2(n2456), .IN3(n18737), .IN4(n2491), .IN5(
        n15010), .Q(n15005) );
  OA221X1 U23530 ( .IN1(n18752), .IN2(n2596), .IN3(n18749), .IN4(n2631), .IN5(
        n15009), .Q(n15006) );
  NAND4X0 U23531 ( .IN1(n14996), .IN2(n14997), .IN3(n14998), .IN4(n14999), 
        .QN(m6_data_o[28]) );
  OA221X1 U23532 ( .IN1(n18730), .IN2(n2385), .IN3(n14912), .IN4(n2420), .IN5(
        n15003), .Q(n14996) );
  OA221X1 U23533 ( .IN1(n18740), .IN2(n2455), .IN3(n18737), .IN4(n2490), .IN5(
        n15002), .Q(n14997) );
  OA221X1 U23534 ( .IN1(n18752), .IN2(n2595), .IN3(n18749), .IN4(n2630), .IN5(
        n15001), .Q(n14998) );
  NAND4X0 U23535 ( .IN1(n14988), .IN2(n14989), .IN3(n14990), .IN4(n14991), 
        .QN(m6_data_o[29]) );
  OA221X1 U23536 ( .IN1(n18728), .IN2(n2384), .IN3(n18725), .IN4(n2419), .IN5(
        n14995), .Q(n14988) );
  OA221X1 U23537 ( .IN1(n18741), .IN2(n2454), .IN3(n18738), .IN4(n2489), .IN5(
        n14994), .Q(n14989) );
  OA221X1 U23538 ( .IN1(n18753), .IN2(n2594), .IN3(n18750), .IN4(n2629), .IN5(
        n14993), .Q(n14990) );
  NAND4X0 U23539 ( .IN1(n14972), .IN2(n14973), .IN3(n14974), .IN4(n14975), 
        .QN(m6_data_o[30]) );
  OA221X1 U23540 ( .IN1(n18730), .IN2(n2383), .IN3(n18726), .IN4(n2418), .IN5(
        n14979), .Q(n14972) );
  OA221X1 U23541 ( .IN1(n18742), .IN2(n2453), .IN3(n18739), .IN4(n2488), .IN5(
        n14978), .Q(n14973) );
  OA221X1 U23542 ( .IN1(n18754), .IN2(n2593), .IN3(n18751), .IN4(n2628), .IN5(
        n14977), .Q(n14974) );
  NAND4X0 U23543 ( .IN1(n14964), .IN2(n14965), .IN3(n14966), .IN4(n14967), 
        .QN(m6_data_o[31]) );
  OA221X1 U23544 ( .IN1(n18730), .IN2(n2382), .IN3(n18725), .IN4(n2417), .IN5(
        n14971), .Q(n14964) );
  OA221X1 U23545 ( .IN1(n18742), .IN2(n2452), .IN3(n18738), .IN4(n2487), .IN5(
        n14970), .Q(n14965) );
  OA221X1 U23546 ( .IN1(n18754), .IN2(n2592), .IN3(n18750), .IN4(n2627), .IN5(
        n14969), .Q(n14966) );
  NAND4X0 U23547 ( .IN1(n15180), .IN2(n15181), .IN3(n15182), .IN4(n15183), 
        .QN(m5_rty_o) );
  OA221X1 U23548 ( .IN1(n8849), .IN2(n2346), .IN3(n8553), .IN4(n2696), .IN5(
        n15188), .Q(n15180) );
  OA221X1 U23549 ( .IN1(n6593), .IN2(n2416), .IN3(n6297), .IN4(n2451), .IN5(
        n15185), .Q(n15182) );
  OA221X1 U23550 ( .IN1(n4817), .IN2(n2626), .IN3(n4521), .IN4(n2661), .IN5(
        n15184), .Q(n15183) );
  NAND4X0 U23551 ( .IN1(n15189), .IN2(n15190), .IN3(n15191), .IN4(n15192), 
        .QN(m5_err_o) );
  OA221X1 U23552 ( .IN1(n8849), .IN2(n2345), .IN3(n8553), .IN4(n2695), .IN5(
        n15196), .Q(n15189) );
  OA221X1 U23553 ( .IN1(n6593), .IN2(n2415), .IN3(n6297), .IN4(n2450), .IN5(
        n15194), .Q(n15191) );
  OA221X1 U23554 ( .IN1(n4817), .IN2(n2625), .IN3(n4521), .IN4(n2660), .IN5(
        n15193), .Q(n15192) );
  NAND4X0 U23555 ( .IN1(n15469), .IN2(n15470), .IN3(n15471), .IN4(n15472), 
        .QN(m5_ack_o) );
  OA221X1 U23556 ( .IN1(n8849), .IN2(n2344), .IN3(n8553), .IN4(n2694), .IN5(
        n15484), .Q(n15469) );
  OA221X1 U23557 ( .IN1(n6593), .IN2(n2414), .IN3(n6297), .IN4(n2449), .IN5(
        n15480), .Q(n15471) );
  OA221X1 U23558 ( .IN1(n4817), .IN2(n2624), .IN3(n4521), .IN4(n2659), .IN5(
        n15473), .Q(n15472) );
  NAND4X0 U23559 ( .IN1(n15461), .IN2(n15462), .IN3(n15463), .IN4(n15464), 
        .QN(m5_data_o[0]) );
  OA221X1 U23560 ( .IN1(n18680), .IN2(n2413), .IN3(n18677), .IN4(n2448), .IN5(
        n15468), .Q(n15461) );
  OA221X1 U23561 ( .IN1(n18693), .IN2(n2483), .IN3(n18689), .IN4(n2518), .IN5(
        n15467), .Q(n15462) );
  OA221X1 U23562 ( .IN1(n18704), .IN2(n2623), .IN3(n18701), .IN4(n2658), .IN5(
        n15466), .Q(n15463) );
  NAND4X0 U23563 ( .IN1(n15373), .IN2(n15374), .IN3(n15375), .IN4(n15376), 
        .QN(m5_data_o[1]) );
  OA221X1 U23564 ( .IN1(n18682), .IN2(n2412), .IN3(n18678), .IN4(n2447), .IN5(
        n15380), .Q(n15373) );
  OA221X1 U23565 ( .IN1(n18692), .IN2(n2482), .IN3(n18689), .IN4(n2517), .IN5(
        n15379), .Q(n15374) );
  OA221X1 U23566 ( .IN1(n18706), .IN2(n2622), .IN3(n18701), .IN4(n2657), .IN5(
        n15378), .Q(n15375) );
  NAND4X0 U23567 ( .IN1(n15285), .IN2(n15286), .IN3(n15287), .IN4(n15288), 
        .QN(m5_data_o[2]) );
  OA221X1 U23568 ( .IN1(n18680), .IN2(n2411), .IN3(n18677), .IN4(n2446), .IN5(
        n15292), .Q(n15285) );
  OA221X1 U23569 ( .IN1(n18692), .IN2(n2481), .IN3(n18691), .IN4(n2516), .IN5(
        n15291), .Q(n15286) );
  OA221X1 U23570 ( .IN1(n18705), .IN2(n2621), .IN3(n18703), .IN4(n2656), .IN5(
        n15290), .Q(n15287) );
  NAND4X0 U23571 ( .IN1(n15261), .IN2(n15262), .IN3(n15263), .IN4(n15264), 
        .QN(m5_data_o[3]) );
  OA221X1 U23572 ( .IN1(n18681), .IN2(n2410), .IN3(n18679), .IN4(n2445), .IN5(
        n15268), .Q(n15261) );
  OA221X1 U23573 ( .IN1(n18694), .IN2(n2480), .IN3(n18690), .IN4(n2515), .IN5(
        n15267), .Q(n15262) );
  OA221X1 U23574 ( .IN1(n18705), .IN2(n2620), .IN3(n18702), .IN4(n2655), .IN5(
        n15266), .Q(n15263) );
  NAND4X0 U23575 ( .IN1(n15253), .IN2(n15254), .IN3(n15255), .IN4(n15256), 
        .QN(m5_data_o[4]) );
  OA221X1 U23576 ( .IN1(n18681), .IN2(n2409), .IN3(n18677), .IN4(n2444), .IN5(
        n15260), .Q(n15253) );
  OA221X1 U23577 ( .IN1(n18693), .IN2(n2479), .IN3(n18690), .IN4(n2514), .IN5(
        n15259), .Q(n15254) );
  OA221X1 U23578 ( .IN1(n18705), .IN2(n2619), .IN3(n18703), .IN4(n2654), .IN5(
        n15258), .Q(n15255) );
  NAND4X0 U23579 ( .IN1(n15245), .IN2(n15246), .IN3(n15247), .IN4(n15248), 
        .QN(m5_data_o[5]) );
  OA221X1 U23580 ( .IN1(n18680), .IN2(n2408), .IN3(n18678), .IN4(n2443), .IN5(
        n15252), .Q(n15245) );
  OA221X1 U23581 ( .IN1(n18694), .IN2(n2478), .IN3(n18690), .IN4(n2513), .IN5(
        n15251), .Q(n15246) );
  OA221X1 U23582 ( .IN1(n18704), .IN2(n2618), .IN3(n18703), .IN4(n2653), .IN5(
        n15250), .Q(n15247) );
  NAND4X0 U23583 ( .IN1(n15237), .IN2(n15238), .IN3(n15239), .IN4(n15240), 
        .QN(m5_data_o[6]) );
  OA221X1 U23584 ( .IN1(n18682), .IN2(n2407), .IN3(n18679), .IN4(n2442), .IN5(
        n15244), .Q(n15237) );
  OA221X1 U23585 ( .IN1(n18694), .IN2(n2477), .IN3(n18691), .IN4(n2512), .IN5(
        n15243), .Q(n15238) );
  OA221X1 U23586 ( .IN1(n18706), .IN2(n2617), .IN3(n18703), .IN4(n2652), .IN5(
        n15242), .Q(n15239) );
  NAND4X0 U23587 ( .IN1(n15229), .IN2(n15230), .IN3(n15231), .IN4(n15232), 
        .QN(m5_data_o[7]) );
  OA221X1 U23588 ( .IN1(n18682), .IN2(n2406), .IN3(n18679), .IN4(n2441), .IN5(
        n15236), .Q(n15229) );
  OA221X1 U23589 ( .IN1(n18694), .IN2(n2476), .IN3(n18691), .IN4(n2511), .IN5(
        n15235), .Q(n15230) );
  OA221X1 U23590 ( .IN1(n18706), .IN2(n2616), .IN3(n18703), .IN4(n2651), .IN5(
        n15234), .Q(n15231) );
  NAND4X0 U23591 ( .IN1(n15221), .IN2(n15222), .IN3(n15223), .IN4(n15224), 
        .QN(m5_data_o[8]) );
  OA221X1 U23592 ( .IN1(n18682), .IN2(n2405), .IN3(n18679), .IN4(n2440), .IN5(
        n15228), .Q(n15221) );
  OA221X1 U23593 ( .IN1(n18694), .IN2(n2475), .IN3(n18691), .IN4(n2510), .IN5(
        n15227), .Q(n15222) );
  OA221X1 U23594 ( .IN1(n18706), .IN2(n2615), .IN3(n18703), .IN4(n2650), .IN5(
        n15226), .Q(n15223) );
  NAND4X0 U23595 ( .IN1(n15197), .IN2(n15198), .IN3(n15199), .IN4(n15200), 
        .QN(m5_data_o[9]) );
  OA221X1 U23596 ( .IN1(n18682), .IN2(n2404), .IN3(n18679), .IN4(n2439), .IN5(
        n15218), .Q(n15197) );
  OA221X1 U23597 ( .IN1(n18694), .IN2(n2474), .IN3(n18691), .IN4(n2509), .IN5(
        n15213), .Q(n15198) );
  OA221X1 U23598 ( .IN1(n18706), .IN2(n2614), .IN3(n18703), .IN4(n2649), .IN5(
        n15208), .Q(n15199) );
  NAND4X0 U23599 ( .IN1(n15453), .IN2(n15454), .IN3(n15455), .IN4(n15456), 
        .QN(m5_data_o[10]) );
  OA221X1 U23600 ( .IN1(n18682), .IN2(n2403), .IN3(n18677), .IN4(n2438), .IN5(
        n15460), .Q(n15453) );
  OA221X1 U23601 ( .IN1(n18694), .IN2(n2473), .IN3(n18689), .IN4(n2508), .IN5(
        n15459), .Q(n15454) );
  OA221X1 U23602 ( .IN1(n18706), .IN2(n2613), .IN3(n18701), .IN4(n2648), .IN5(
        n15458), .Q(n15455) );
  NAND4X0 U23603 ( .IN1(n15445), .IN2(n15446), .IN3(n15447), .IN4(n15448), 
        .QN(m5_data_o[11]) );
  OA221X1 U23604 ( .IN1(n18681), .IN2(n2402), .IN3(n18677), .IN4(n2437), .IN5(
        n15452), .Q(n15445) );
  OA221X1 U23605 ( .IN1(n18692), .IN2(n2472), .IN3(n18689), .IN4(n2507), .IN5(
        n15451), .Q(n15446) );
  OA221X1 U23606 ( .IN1(n18705), .IN2(n2612), .IN3(n18701), .IN4(n2647), .IN5(
        n15450), .Q(n15447) );
  NAND4X0 U23607 ( .IN1(n15437), .IN2(n15438), .IN3(n15439), .IN4(n15440), 
        .QN(m5_data_o[12]) );
  OA221X1 U23608 ( .IN1(n18680), .IN2(n2401), .IN3(n18677), .IN4(n2436), .IN5(
        n15444), .Q(n15437) );
  OA221X1 U23609 ( .IN1(n18693), .IN2(n2471), .IN3(n18689), .IN4(n2506), .IN5(
        n15443), .Q(n15438) );
  OA221X1 U23610 ( .IN1(n18704), .IN2(n2611), .IN3(n18701), .IN4(n2646), .IN5(
        n15442), .Q(n15439) );
  NAND4X0 U23611 ( .IN1(n15429), .IN2(n15430), .IN3(n15431), .IN4(n15432), 
        .QN(m5_data_o[13]) );
  OA221X1 U23612 ( .IN1(n18680), .IN2(n2400), .IN3(n18678), .IN4(n2435), .IN5(
        n15436), .Q(n15429) );
  OA221X1 U23613 ( .IN1(n18694), .IN2(n2470), .IN3(n18691), .IN4(n2505), .IN5(
        n15435), .Q(n15430) );
  OA221X1 U23614 ( .IN1(n18706), .IN2(n2610), .IN3(n18702), .IN4(n2645), .IN5(
        n15434), .Q(n15431) );
  NAND4X0 U23615 ( .IN1(n15421), .IN2(n15422), .IN3(n15423), .IN4(n15424), 
        .QN(m5_data_o[14]) );
  OA221X1 U23616 ( .IN1(n18682), .IN2(n2399), .IN3(n18678), .IN4(n2434), .IN5(
        n15428), .Q(n15421) );
  OA221X1 U23617 ( .IN1(n18692), .IN2(n2469), .IN3(n18689), .IN4(n2504), .IN5(
        n15427), .Q(n15422) );
  OA221X1 U23618 ( .IN1(n18704), .IN2(n2609), .IN3(n18702), .IN4(n2644), .IN5(
        n15426), .Q(n15423) );
  NAND4X0 U23619 ( .IN1(n15413), .IN2(n15414), .IN3(n15415), .IN4(n15416), 
        .QN(m5_data_o[15]) );
  OA221X1 U23620 ( .IN1(n18681), .IN2(n2398), .IN3(n18678), .IN4(n2433), .IN5(
        n15420), .Q(n15413) );
  OA221X1 U23621 ( .IN1(n18692), .IN2(n2468), .IN3(n18690), .IN4(n2503), .IN5(
        n15419), .Q(n15414) );
  OA221X1 U23622 ( .IN1(n18704), .IN2(n2608), .IN3(n18702), .IN4(n2643), .IN5(
        n15418), .Q(n15415) );
  NAND4X0 U23623 ( .IN1(n15405), .IN2(n15406), .IN3(n15407), .IN4(n15408), 
        .QN(m5_data_o[16]) );
  OA221X1 U23624 ( .IN1(n18680), .IN2(n2397), .IN3(n18678), .IN4(n2432), .IN5(
        n15412), .Q(n15405) );
  OA221X1 U23625 ( .IN1(n18693), .IN2(n2467), .IN3(n18690), .IN4(n2502), .IN5(
        n15411), .Q(n15406) );
  OA221X1 U23626 ( .IN1(n18705), .IN2(n2607), .IN3(n18702), .IN4(n2642), .IN5(
        n15410), .Q(n15407) );
  NAND4X0 U23627 ( .IN1(n15397), .IN2(n15398), .IN3(n15399), .IN4(n15400), 
        .QN(m5_data_o[17]) );
  OA221X1 U23628 ( .IN1(n18681), .IN2(n2396), .IN3(n18679), .IN4(n2431), .IN5(
        n15404), .Q(n15397) );
  OA221X1 U23629 ( .IN1(n18694), .IN2(n2466), .IN3(n18691), .IN4(n2501), .IN5(
        n15403), .Q(n15398) );
  OA221X1 U23630 ( .IN1(n18705), .IN2(n2606), .IN3(n18702), .IN4(n2641), .IN5(
        n15402), .Q(n15399) );
  NAND4X0 U23631 ( .IN1(n15389), .IN2(n15390), .IN3(n15391), .IN4(n15392), 
        .QN(m5_data_o[18]) );
  OA221X1 U23632 ( .IN1(n18681), .IN2(n2395), .IN3(n18677), .IN4(n2430), .IN5(
        n15396), .Q(n15389) );
  OA221X1 U23633 ( .IN1(n18693), .IN2(n2465), .IN3(n18689), .IN4(n2500), .IN5(
        n15395), .Q(n15390) );
  OA221X1 U23634 ( .IN1(n18705), .IN2(n2605), .IN3(n18703), .IN4(n2640), .IN5(
        n15394), .Q(n15391) );
  NAND4X0 U23635 ( .IN1(n15381), .IN2(n15382), .IN3(n15383), .IN4(n15384), 
        .QN(m5_data_o[19]) );
  OA221X1 U23636 ( .IN1(n18682), .IN2(n2394), .IN3(n18678), .IN4(n2429), .IN5(
        n15388), .Q(n15381) );
  OA221X1 U23637 ( .IN1(n18692), .IN2(n2464), .IN3(n18689), .IN4(n2499), .IN5(
        n15387), .Q(n15382) );
  OA221X1 U23638 ( .IN1(n18706), .IN2(n2604), .IN3(n18701), .IN4(n2639), .IN5(
        n15386), .Q(n15383) );
  NAND4X0 U23639 ( .IN1(n15365), .IN2(n15366), .IN3(n15367), .IN4(n15368), 
        .QN(m5_data_o[20]) );
  OA221X1 U23640 ( .IN1(n18680), .IN2(n2393), .IN3(n18677), .IN4(n2428), .IN5(
        n15372), .Q(n15365) );
  OA221X1 U23641 ( .IN1(n18692), .IN2(n2463), .IN3(n18690), .IN4(n2498), .IN5(
        n15371), .Q(n15366) );
  OA221X1 U23642 ( .IN1(n18704), .IN2(n2603), .IN3(n18701), .IN4(n2638), .IN5(
        n15370), .Q(n15367) );
  NAND4X0 U23643 ( .IN1(n15357), .IN2(n15358), .IN3(n15359), .IN4(n15360), 
        .QN(m5_data_o[21]) );
  OA221X1 U23644 ( .IN1(n18680), .IN2(n2392), .IN3(n18678), .IN4(n2427), .IN5(
        n15364), .Q(n15357) );
  OA221X1 U23645 ( .IN1(n18692), .IN2(n2462), .IN3(n18690), .IN4(n2497), .IN5(
        n15363), .Q(n15358) );
  OA221X1 U23646 ( .IN1(n18704), .IN2(n2602), .IN3(n18702), .IN4(n2637), .IN5(
        n15362), .Q(n15359) );
  NAND4X0 U23647 ( .IN1(n15349), .IN2(n15350), .IN3(n15351), .IN4(n15352), 
        .QN(m5_data_o[22]) );
  OA221X1 U23648 ( .IN1(n18680), .IN2(n2391), .IN3(n18679), .IN4(n2426), .IN5(
        n15356), .Q(n15349) );
  OA221X1 U23649 ( .IN1(n18692), .IN2(n2461), .IN3(n18690), .IN4(n2496), .IN5(
        n15355), .Q(n15350) );
  OA221X1 U23650 ( .IN1(n18704), .IN2(n2601), .IN3(n18703), .IN4(n2636), .IN5(
        n15354), .Q(n15351) );
  NAND4X0 U23651 ( .IN1(n15341), .IN2(n15342), .IN3(n15343), .IN4(n15344), 
        .QN(m5_data_o[23]) );
  OA221X1 U23652 ( .IN1(n18680), .IN2(n2390), .IN3(n18677), .IN4(n2425), .IN5(
        n15348), .Q(n15341) );
  OA221X1 U23653 ( .IN1(n18692), .IN2(n2460), .IN3(n18690), .IN4(n2495), .IN5(
        n15347), .Q(n15342) );
  OA221X1 U23654 ( .IN1(n18704), .IN2(n2600), .IN3(n18701), .IN4(n2635), .IN5(
        n15346), .Q(n15343) );
  NAND4X0 U23655 ( .IN1(n15333), .IN2(n15334), .IN3(n15335), .IN4(n15336), 
        .QN(m5_data_o[24]) );
  OA221X1 U23656 ( .IN1(n18681), .IN2(n2389), .IN3(n18679), .IN4(n2424), .IN5(
        n15340), .Q(n15333) );
  OA221X1 U23657 ( .IN1(n18693), .IN2(n2459), .IN3(n18691), .IN4(n2494), .IN5(
        n15339), .Q(n15334) );
  OA221X1 U23658 ( .IN1(n18704), .IN2(n2599), .IN3(n18701), .IN4(n2634), .IN5(
        n15338), .Q(n15335) );
  NAND4X0 U23659 ( .IN1(n15325), .IN2(n15326), .IN3(n15327), .IN4(n15328), 
        .QN(m5_data_o[25]) );
  OA221X1 U23660 ( .IN1(n18681), .IN2(n2388), .IN3(n18679), .IN4(n2423), .IN5(
        n15332), .Q(n15325) );
  OA221X1 U23661 ( .IN1(n18693), .IN2(n2458), .IN3(n18689), .IN4(n2493), .IN5(
        n15331), .Q(n15326) );
  OA221X1 U23662 ( .IN1(n18706), .IN2(n2598), .IN3(n18702), .IN4(n2633), .IN5(
        n15330), .Q(n15327) );
  NAND4X0 U23663 ( .IN1(n15317), .IN2(n15318), .IN3(n15319), .IN4(n15320), 
        .QN(m5_data_o[26]) );
  OA221X1 U23664 ( .IN1(n18681), .IN2(n2387), .IN3(n18677), .IN4(n2422), .IN5(
        n15324), .Q(n15317) );
  OA221X1 U23665 ( .IN1(n18693), .IN2(n2457), .IN3(n18690), .IN4(n2492), .IN5(
        n15323), .Q(n15318) );
  OA221X1 U23666 ( .IN1(n18705), .IN2(n2597), .IN3(n18703), .IN4(n2632), .IN5(
        n15322), .Q(n15319) );
  NAND4X0 U23667 ( .IN1(n15309), .IN2(n15310), .IN3(n15311), .IN4(n15312), 
        .QN(m5_data_o[27]) );
  OA221X1 U23668 ( .IN1(n18681), .IN2(n2386), .IN3(n18678), .IN4(n2421), .IN5(
        n15316), .Q(n15309) );
  OA221X1 U23669 ( .IN1(n18693), .IN2(n2456), .IN3(n18691), .IN4(n2491), .IN5(
        n15315), .Q(n15310) );
  OA221X1 U23670 ( .IN1(n18704), .IN2(n2596), .IN3(n18701), .IN4(n2631), .IN5(
        n15314), .Q(n15311) );
  NAND4X0 U23671 ( .IN1(n15301), .IN2(n15302), .IN3(n15303), .IN4(n15304), 
        .QN(m5_data_o[28]) );
  OA221X1 U23672 ( .IN1(n18682), .IN2(n2385), .IN3(n18678), .IN4(n2420), .IN5(
        n15308), .Q(n15301) );
  OA221X1 U23673 ( .IN1(n18693), .IN2(n2455), .IN3(n18691), .IN4(n2490), .IN5(
        n15307), .Q(n15302) );
  OA221X1 U23674 ( .IN1(n18705), .IN2(n2595), .IN3(n18701), .IN4(n2630), .IN5(
        n15306), .Q(n15303) );
  NAND4X0 U23675 ( .IN1(n15293), .IN2(n15294), .IN3(n15295), .IN4(n15296), 
        .QN(m5_data_o[29]) );
  OA221X1 U23676 ( .IN1(n18681), .IN2(n2384), .IN3(n18679), .IN4(n2419), .IN5(
        n15300), .Q(n15293) );
  OA221X1 U23677 ( .IN1(n18693), .IN2(n2454), .IN3(n18690), .IN4(n2489), .IN5(
        n15299), .Q(n15294) );
  OA221X1 U23678 ( .IN1(n18705), .IN2(n2594), .IN3(n18702), .IN4(n2629), .IN5(
        n15298), .Q(n15295) );
  NAND4X0 U23679 ( .IN1(n15277), .IN2(n15278), .IN3(n15279), .IN4(n15280), 
        .QN(m5_data_o[30]) );
  OA221X1 U23680 ( .IN1(n18680), .IN2(n2383), .IN3(n18677), .IN4(n2418), .IN5(
        n15284), .Q(n15277) );
  OA221X1 U23681 ( .IN1(n18694), .IN2(n2453), .IN3(n18689), .IN4(n2488), .IN5(
        n15283), .Q(n15278) );
  OA221X1 U23682 ( .IN1(n18705), .IN2(n2593), .IN3(n18703), .IN4(n2628), .IN5(
        n15282), .Q(n15279) );
  NAND4X0 U23683 ( .IN1(n15269), .IN2(n15270), .IN3(n15271), .IN4(n15272), 
        .QN(m5_data_o[31]) );
  OA221X1 U23684 ( .IN1(n18682), .IN2(n2382), .IN3(n18679), .IN4(n2417), .IN5(
        n15276), .Q(n15269) );
  OA221X1 U23685 ( .IN1(n18692), .IN2(n2452), .IN3(n18691), .IN4(n2487), .IN5(
        n15275), .Q(n15270) );
  OA221X1 U23686 ( .IN1(n18706), .IN2(n2592), .IN3(n18702), .IN4(n2627), .IN5(
        n15274), .Q(n15271) );
  NAND4X0 U23687 ( .IN1(n15485), .IN2(n15486), .IN3(n15487), .IN4(n15488), 
        .QN(m4_rty_o) );
  OA221X1 U23688 ( .IN1(n8850), .IN2(n2346), .IN3(n8554), .IN4(n2696), .IN5(
        n15493), .Q(n15485) );
  OA221X1 U23689 ( .IN1(n6594), .IN2(n2416), .IN3(n6298), .IN4(n2451), .IN5(
        n15490), .Q(n15487) );
  OA221X1 U23690 ( .IN1(n4818), .IN2(n2626), .IN3(n4522), .IN4(n2661), .IN5(
        n15489), .Q(n15488) );
  NAND4X0 U23691 ( .IN1(n15494), .IN2(n15495), .IN3(n15496), .IN4(n15497), 
        .QN(m4_err_o) );
  OA221X1 U23692 ( .IN1(n8850), .IN2(n2345), .IN3(n8554), .IN4(n2695), .IN5(
        n15501), .Q(n15494) );
  OA221X1 U23693 ( .IN1(n6594), .IN2(n2415), .IN3(n6298), .IN4(n2450), .IN5(
        n15499), .Q(n15496) );
  OA221X1 U23694 ( .IN1(n4818), .IN2(n2625), .IN3(n4522), .IN4(n2660), .IN5(
        n15498), .Q(n15497) );
  NAND4X0 U23695 ( .IN1(n15774), .IN2(n15775), .IN3(n15776), .IN4(n15777), 
        .QN(m4_ack_o) );
  OA221X1 U23696 ( .IN1(n8850), .IN2(n2344), .IN3(n8554), .IN4(n2694), .IN5(
        n15789), .Q(n15774) );
  OA221X1 U23697 ( .IN1(n6594), .IN2(n2414), .IN3(n6298), .IN4(n2449), .IN5(
        n15785), .Q(n15776) );
  OA221X1 U23698 ( .IN1(n4818), .IN2(n2624), .IN3(n4522), .IN4(n2659), .IN5(
        n15778), .Q(n15777) );
  NAND4X0 U23699 ( .IN1(n15766), .IN2(n15767), .IN3(n15768), .IN4(n15769), 
        .QN(m4_data_o[0]) );
  OA221X1 U23700 ( .IN1(n18632), .IN2(n2413), .IN3(n15522), .IN4(n2448), .IN5(
        n15773), .Q(n15766) );
  OA221X1 U23701 ( .IN1(n18644), .IN2(n2483), .IN3(n18641), .IN4(n2518), .IN5(
        n15772), .Q(n15767) );
  OA221X1 U23702 ( .IN1(n18657), .IN2(n2623), .IN3(n18653), .IN4(n2658), .IN5(
        n15771), .Q(n15768) );
  NAND4X0 U23703 ( .IN1(n15678), .IN2(n15679), .IN3(n15680), .IN4(n15681), 
        .QN(m4_data_o[1]) );
  OA221X1 U23704 ( .IN1(n18634), .IN2(n2412), .IN3(n18630), .IN4(n2447), .IN5(
        n15685), .Q(n15678) );
  OA221X1 U23705 ( .IN1(n18646), .IN2(n2482), .IN3(n18641), .IN4(n2517), .IN5(
        n15684), .Q(n15679) );
  OA221X1 U23706 ( .IN1(n18658), .IN2(n2622), .IN3(n18653), .IN4(n2657), .IN5(
        n15683), .Q(n15680) );
  NAND4X0 U23707 ( .IN1(n15590), .IN2(n15591), .IN3(n15592), .IN4(n15593), 
        .QN(m4_data_o[2]) );
  OA221X1 U23708 ( .IN1(n18632), .IN2(n2411), .IN3(n18630), .IN4(n2446), .IN5(
        n15597), .Q(n15590) );
  OA221X1 U23709 ( .IN1(n18646), .IN2(n2481), .IN3(n18643), .IN4(n2516), .IN5(
        n15596), .Q(n15591) );
  OA221X1 U23710 ( .IN1(n18658), .IN2(n2621), .IN3(n18654), .IN4(n2656), .IN5(
        n15595), .Q(n15592) );
  NAND4X0 U23711 ( .IN1(n15566), .IN2(n15567), .IN3(n15568), .IN4(n15569), 
        .QN(m4_data_o[3]) );
  OA221X1 U23712 ( .IN1(n18634), .IN2(n2410), .IN3(n18630), .IN4(n2445), .IN5(
        n15573), .Q(n15566) );
  OA221X1 U23713 ( .IN1(n18646), .IN2(n2480), .IN3(n18642), .IN4(n2515), .IN5(
        n15572), .Q(n15567) );
  OA221X1 U23714 ( .IN1(n18658), .IN2(n2620), .IN3(n18654), .IN4(n2655), .IN5(
        n15571), .Q(n15568) );
  NAND4X0 U23715 ( .IN1(n15558), .IN2(n15559), .IN3(n15560), .IN4(n15561), 
        .QN(m4_data_o[4]) );
  OA221X1 U23716 ( .IN1(n18632), .IN2(n2409), .IN3(n18629), .IN4(n2444), .IN5(
        n15565), .Q(n15558) );
  OA221X1 U23717 ( .IN1(n18644), .IN2(n2479), .IN3(n18643), .IN4(n2514), .IN5(
        n15564), .Q(n15559) );
  OA221X1 U23718 ( .IN1(n18657), .IN2(n2619), .IN3(n18655), .IN4(n2654), .IN5(
        n15563), .Q(n15560) );
  NAND4X0 U23719 ( .IN1(n15550), .IN2(n15551), .IN3(n15552), .IN4(n15553), 
        .QN(m4_data_o[5]) );
  OA221X1 U23720 ( .IN1(n18633), .IN2(n2408), .IN3(n15522), .IN4(n2443), .IN5(
        n15557), .Q(n15550) );
  OA221X1 U23721 ( .IN1(n18645), .IN2(n2478), .IN3(n18643), .IN4(n2513), .IN5(
        n15556), .Q(n15551) );
  OA221X1 U23722 ( .IN1(n18656), .IN2(n2618), .IN3(n18654), .IN4(n2653), .IN5(
        n15555), .Q(n15552) );
  NAND4X0 U23723 ( .IN1(n15542), .IN2(n15543), .IN3(n15544), .IN4(n15545), 
        .QN(m4_data_o[6]) );
  OA221X1 U23724 ( .IN1(n18634), .IN2(n2407), .IN3(n18630), .IN4(n2442), .IN5(
        n15549), .Q(n15542) );
  OA221X1 U23725 ( .IN1(n18646), .IN2(n2477), .IN3(n18643), .IN4(n2512), .IN5(
        n15548), .Q(n15543) );
  OA221X1 U23726 ( .IN1(n18658), .IN2(n2617), .IN3(n18655), .IN4(n2652), .IN5(
        n15547), .Q(n15544) );
  NAND4X0 U23727 ( .IN1(n15534), .IN2(n15535), .IN3(n15536), .IN4(n15537), 
        .QN(m4_data_o[7]) );
  OA221X1 U23728 ( .IN1(n18634), .IN2(n2406), .IN3(n18630), .IN4(n2441), .IN5(
        n15541), .Q(n15534) );
  OA221X1 U23729 ( .IN1(n18646), .IN2(n2476), .IN3(n18643), .IN4(n2511), .IN5(
        n15540), .Q(n15535) );
  OA221X1 U23730 ( .IN1(n18658), .IN2(n2616), .IN3(n18655), .IN4(n2651), .IN5(
        n15539), .Q(n15536) );
  NAND4X0 U23731 ( .IN1(n15526), .IN2(n15527), .IN3(n15528), .IN4(n15529), 
        .QN(m4_data_o[8]) );
  OA221X1 U23732 ( .IN1(n18634), .IN2(n2405), .IN3(n18630), .IN4(n2440), .IN5(
        n15533), .Q(n15526) );
  OA221X1 U23733 ( .IN1(n18646), .IN2(n2475), .IN3(n18643), .IN4(n2510), .IN5(
        n15532), .Q(n15527) );
  OA221X1 U23734 ( .IN1(n18658), .IN2(n2615), .IN3(n18655), .IN4(n2650), .IN5(
        n15531), .Q(n15528) );
  NAND4X0 U23735 ( .IN1(n15502), .IN2(n15503), .IN3(n15504), .IN4(n15505), 
        .QN(m4_data_o[9]) );
  OA221X1 U23736 ( .IN1(n18634), .IN2(n2404), .IN3(n18630), .IN4(n2439), .IN5(
        n15523), .Q(n15502) );
  OA221X1 U23737 ( .IN1(n18646), .IN2(n2474), .IN3(n18643), .IN4(n2509), .IN5(
        n15518), .Q(n15503) );
  OA221X1 U23738 ( .IN1(n18658), .IN2(n2614), .IN3(n18655), .IN4(n2649), .IN5(
        n15513), .Q(n15504) );
  NAND4X0 U23739 ( .IN1(n15758), .IN2(n15759), .IN3(n15760), .IN4(n15761), 
        .QN(m4_data_o[10]) );
  OA221X1 U23740 ( .IN1(n18633), .IN2(n2403), .IN3(n15522), .IN4(n2438), .IN5(
        n15765), .Q(n15758) );
  OA221X1 U23741 ( .IN1(n18646), .IN2(n2473), .IN3(n18641), .IN4(n2508), .IN5(
        n15764), .Q(n15759) );
  OA221X1 U23742 ( .IN1(n18656), .IN2(n2613), .IN3(n18653), .IN4(n2648), .IN5(
        n15763), .Q(n15760) );
  NAND4X0 U23743 ( .IN1(n15750), .IN2(n15751), .IN3(n15752), .IN4(n15753), 
        .QN(m4_data_o[11]) );
  OA221X1 U23744 ( .IN1(n18632), .IN2(n2402), .IN3(n15522), .IN4(n2437), .IN5(
        n15757), .Q(n15750) );
  OA221X1 U23745 ( .IN1(n18644), .IN2(n2472), .IN3(n18641), .IN4(n2507), .IN5(
        n15756), .Q(n15751) );
  OA221X1 U23746 ( .IN1(n18658), .IN2(n2612), .IN3(n18653), .IN4(n2647), .IN5(
        n15755), .Q(n15752) );
  NAND4X0 U23747 ( .IN1(n15742), .IN2(n15743), .IN3(n15744), .IN4(n15745), 
        .QN(m4_data_o[12]) );
  OA221X1 U23748 ( .IN1(n18633), .IN2(n2401), .IN3(n15522), .IN4(n2436), .IN5(
        n15749), .Q(n15742) );
  OA221X1 U23749 ( .IN1(n18645), .IN2(n2471), .IN3(n18641), .IN4(n2506), .IN5(
        n15748), .Q(n15743) );
  OA221X1 U23750 ( .IN1(n18657), .IN2(n2611), .IN3(n18653), .IN4(n2646), .IN5(
        n15747), .Q(n15744) );
  NAND4X0 U23751 ( .IN1(n15734), .IN2(n15735), .IN3(n15736), .IN4(n15737), 
        .QN(m4_data_o[13]) );
  OA221X1 U23752 ( .IN1(n18632), .IN2(n2400), .IN3(n18629), .IN4(n2435), .IN5(
        n15741), .Q(n15734) );
  OA221X1 U23753 ( .IN1(n18644), .IN2(n2470), .IN3(n18642), .IN4(n2505), .IN5(
        n15740), .Q(n15735) );
  OA221X1 U23754 ( .IN1(n18656), .IN2(n2610), .IN3(n18655), .IN4(n2645), .IN5(
        n15739), .Q(n15736) );
  NAND4X0 U23755 ( .IN1(n15726), .IN2(n15727), .IN3(n15728), .IN4(n15729), 
        .QN(m4_data_o[14]) );
  OA221X1 U23756 ( .IN1(n18632), .IN2(n2399), .IN3(n18629), .IN4(n2434), .IN5(
        n15733), .Q(n15726) );
  OA221X1 U23757 ( .IN1(n18644), .IN2(n2469), .IN3(n18642), .IN4(n2504), .IN5(
        n15732), .Q(n15727) );
  OA221X1 U23758 ( .IN1(n18656), .IN2(n2609), .IN3(n18653), .IN4(n2644), .IN5(
        n15731), .Q(n15728) );
  NAND4X0 U23759 ( .IN1(n15718), .IN2(n15719), .IN3(n15720), .IN4(n15721), 
        .QN(m4_data_o[15]) );
  OA221X1 U23760 ( .IN1(n18632), .IN2(n2398), .IN3(n18629), .IN4(n2433), .IN5(
        n15725), .Q(n15718) );
  OA221X1 U23761 ( .IN1(n18644), .IN2(n2468), .IN3(n18642), .IN4(n2503), .IN5(
        n15724), .Q(n15719) );
  OA221X1 U23762 ( .IN1(n18656), .IN2(n2608), .IN3(n18654), .IN4(n2643), .IN5(
        n15723), .Q(n15720) );
  NAND4X0 U23763 ( .IN1(n15710), .IN2(n15711), .IN3(n15712), .IN4(n15713), 
        .QN(m4_data_o[16]) );
  OA221X1 U23764 ( .IN1(n18632), .IN2(n2397), .IN3(n18629), .IN4(n2432), .IN5(
        n15717), .Q(n15710) );
  OA221X1 U23765 ( .IN1(n18644), .IN2(n2467), .IN3(n18642), .IN4(n2502), .IN5(
        n15716), .Q(n15711) );
  OA221X1 U23766 ( .IN1(n18656), .IN2(n2607), .IN3(n18654), .IN4(n2642), .IN5(
        n15715), .Q(n15712) );
  NAND4X0 U23767 ( .IN1(n15702), .IN2(n15703), .IN3(n15704), .IN4(n15705), 
        .QN(m4_data_o[17]) );
  OA221X1 U23768 ( .IN1(n18633), .IN2(n2396), .IN3(n18629), .IN4(n2431), .IN5(
        n15709), .Q(n15702) );
  OA221X1 U23769 ( .IN1(n18645), .IN2(n2466), .IN3(n18642), .IN4(n2501), .IN5(
        n15708), .Q(n15703) );
  OA221X1 U23770 ( .IN1(n18656), .IN2(n2606), .IN3(n18655), .IN4(n2641), .IN5(
        n15707), .Q(n15704) );
  NAND4X0 U23771 ( .IN1(n15694), .IN2(n15695), .IN3(n15696), .IN4(n15697), 
        .QN(m4_data_o[18]) );
  OA221X1 U23772 ( .IN1(n18633), .IN2(n2395), .IN3(n18630), .IN4(n2430), .IN5(
        n15701), .Q(n15694) );
  OA221X1 U23773 ( .IN1(n18645), .IN2(n2465), .IN3(n18643), .IN4(n2500), .IN5(
        n15700), .Q(n15695) );
  OA221X1 U23774 ( .IN1(n18657), .IN2(n2605), .IN3(n18653), .IN4(n2640), .IN5(
        n15699), .Q(n15696) );
  NAND4X0 U23775 ( .IN1(n15686), .IN2(n15687), .IN3(n15688), .IN4(n15689), 
        .QN(m4_data_o[19]) );
  OA221X1 U23776 ( .IN1(n18632), .IN2(n2394), .IN3(n18630), .IN4(n2429), .IN5(
        n15693), .Q(n15686) );
  OA221X1 U23777 ( .IN1(n18644), .IN2(n2464), .IN3(n18641), .IN4(n2499), .IN5(
        n15692), .Q(n15687) );
  OA221X1 U23778 ( .IN1(n18658), .IN2(n2604), .IN3(n18653), .IN4(n2639), .IN5(
        n15691), .Q(n15688) );
  NAND4X0 U23779 ( .IN1(n15670), .IN2(n15671), .IN3(n15672), .IN4(n15673), 
        .QN(m4_data_o[20]) );
  OA221X1 U23780 ( .IN1(n18633), .IN2(n2393), .IN3(n15522), .IN4(n2428), .IN5(
        n15677), .Q(n15670) );
  OA221X1 U23781 ( .IN1(n18645), .IN2(n2463), .IN3(n18641), .IN4(n2498), .IN5(
        n15676), .Q(n15671) );
  OA221X1 U23782 ( .IN1(n18656), .IN2(n2603), .IN3(n18654), .IN4(n2638), .IN5(
        n15675), .Q(n15672) );
  NAND4X0 U23783 ( .IN1(n15662), .IN2(n15663), .IN3(n15664), .IN4(n15665), 
        .QN(m4_data_o[21]) );
  OA221X1 U23784 ( .IN1(n18633), .IN2(n2392), .IN3(n15522), .IN4(n2427), .IN5(
        n15669), .Q(n15662) );
  OA221X1 U23785 ( .IN1(n18645), .IN2(n2462), .IN3(n18642), .IN4(n2497), .IN5(
        n15668), .Q(n15663) );
  OA221X1 U23786 ( .IN1(n18656), .IN2(n2602), .IN3(n18654), .IN4(n2637), .IN5(
        n15667), .Q(n15664) );
  NAND4X0 U23787 ( .IN1(n15654), .IN2(n15655), .IN3(n15656), .IN4(n15657), 
        .QN(m4_data_o[22]) );
  OA221X1 U23788 ( .IN1(n18633), .IN2(n2391), .IN3(n15522), .IN4(n2426), .IN5(
        n15661), .Q(n15654) );
  OA221X1 U23789 ( .IN1(n18645), .IN2(n2461), .IN3(n18643), .IN4(n2496), .IN5(
        n15660), .Q(n15655) );
  OA221X1 U23790 ( .IN1(n18657), .IN2(n2601), .IN3(n18654), .IN4(n2636), .IN5(
        n15659), .Q(n15656) );
  NAND4X0 U23791 ( .IN1(n15646), .IN2(n15647), .IN3(n15648), .IN4(n15649), 
        .QN(m4_data_o[23]) );
  OA221X1 U23792 ( .IN1(n18633), .IN2(n2390), .IN3(n15522), .IN4(n2425), .IN5(
        n15653), .Q(n15646) );
  OA221X1 U23793 ( .IN1(n18645), .IN2(n2460), .IN3(n18641), .IN4(n2495), .IN5(
        n15652), .Q(n15647) );
  OA221X1 U23794 ( .IN1(n18658), .IN2(n2600), .IN3(n18654), .IN4(n2635), .IN5(
        n15651), .Q(n15648) );
  NAND4X0 U23795 ( .IN1(n15638), .IN2(n15639), .IN3(n15640), .IN4(n15641), 
        .QN(m4_data_o[24]) );
  OA221X1 U23796 ( .IN1(n18633), .IN2(n2389), .IN3(n18629), .IN4(n2424), .IN5(
        n15645), .Q(n15638) );
  OA221X1 U23797 ( .IN1(n18645), .IN2(n2459), .IN3(n18641), .IN4(n2494), .IN5(
        n15644), .Q(n15639) );
  OA221X1 U23798 ( .IN1(n18657), .IN2(n2599), .IN3(n18655), .IN4(n2634), .IN5(
        n15643), .Q(n15640) );
  NAND4X0 U23799 ( .IN1(n15630), .IN2(n15631), .IN3(n15632), .IN4(n15633), 
        .QN(m4_data_o[25]) );
  OA221X1 U23800 ( .IN1(n18634), .IN2(n2388), .IN3(n18629), .IN4(n2423), .IN5(
        n15637), .Q(n15630) );
  OA221X1 U23801 ( .IN1(n18646), .IN2(n2458), .IN3(n18642), .IN4(n2493), .IN5(
        n15636), .Q(n15631) );
  OA221X1 U23802 ( .IN1(n18657), .IN2(n2598), .IN3(n18653), .IN4(n2633), .IN5(
        n15635), .Q(n15632) );
  NAND4X0 U23803 ( .IN1(n15622), .IN2(n15623), .IN3(n15624), .IN4(n15625), 
        .QN(m4_data_o[26]) );
  OA221X1 U23804 ( .IN1(n18633), .IN2(n2387), .IN3(n15522), .IN4(n2422), .IN5(
        n15629), .Q(n15622) );
  OA221X1 U23805 ( .IN1(n18645), .IN2(n2457), .IN3(n18643), .IN4(n2492), .IN5(
        n15628), .Q(n15623) );
  OA221X1 U23806 ( .IN1(n18657), .IN2(n2597), .IN3(n18654), .IN4(n2632), .IN5(
        n15627), .Q(n15624) );
  NAND4X0 U23807 ( .IN1(n15614), .IN2(n15615), .IN3(n15616), .IN4(n15617), 
        .QN(m4_data_o[27]) );
  OA221X1 U23808 ( .IN1(n18632), .IN2(n2386), .IN3(n15522), .IN4(n2421), .IN5(
        n15621), .Q(n15614) );
  OA221X1 U23809 ( .IN1(n18644), .IN2(n2456), .IN3(n18641), .IN4(n2491), .IN5(
        n15620), .Q(n15615) );
  OA221X1 U23810 ( .IN1(n18657), .IN2(n2596), .IN3(n18655), .IN4(n2631), .IN5(
        n15619), .Q(n15616) );
  NAND4X0 U23811 ( .IN1(n15606), .IN2(n15607), .IN3(n15608), .IN4(n15609), 
        .QN(m4_data_o[28]) );
  OA221X1 U23812 ( .IN1(n18634), .IN2(n2385), .IN3(n15522), .IN4(n2420), .IN5(
        n15613), .Q(n15606) );
  OA221X1 U23813 ( .IN1(n18644), .IN2(n2455), .IN3(n18641), .IN4(n2490), .IN5(
        n15612), .Q(n15607) );
  OA221X1 U23814 ( .IN1(n18658), .IN2(n2595), .IN3(n18655), .IN4(n2630), .IN5(
        n15611), .Q(n15608) );
  NAND4X0 U23815 ( .IN1(n15598), .IN2(n15599), .IN3(n15600), .IN4(n15601), 
        .QN(m4_data_o[29]) );
  OA221X1 U23816 ( .IN1(n18632), .IN2(n2384), .IN3(n18629), .IN4(n2419), .IN5(
        n15605), .Q(n15598) );
  OA221X1 U23817 ( .IN1(n18645), .IN2(n2454), .IN3(n18642), .IN4(n2489), .IN5(
        n15604), .Q(n15599) );
  OA221X1 U23818 ( .IN1(n18656), .IN2(n2594), .IN3(n18653), .IN4(n2629), .IN5(
        n15603), .Q(n15600) );
  NAND4X0 U23819 ( .IN1(n15582), .IN2(n15583), .IN3(n15584), .IN4(n15585), 
        .QN(m4_data_o[30]) );
  OA221X1 U23820 ( .IN1(n18634), .IN2(n2383), .IN3(n18630), .IN4(n2418), .IN5(
        n15589), .Q(n15582) );
  OA221X1 U23821 ( .IN1(n18646), .IN2(n2453), .IN3(n18643), .IN4(n2488), .IN5(
        n15588), .Q(n15583) );
  OA221X1 U23822 ( .IN1(n18657), .IN2(n2593), .IN3(n18654), .IN4(n2628), .IN5(
        n15587), .Q(n15584) );
  NAND4X0 U23823 ( .IN1(n15574), .IN2(n15575), .IN3(n15576), .IN4(n15577), 
        .QN(m4_data_o[31]) );
  OA221X1 U23824 ( .IN1(n18634), .IN2(n2382), .IN3(n18629), .IN4(n2417), .IN5(
        n15581), .Q(n15574) );
  OA221X1 U23825 ( .IN1(n18646), .IN2(n2452), .IN3(n18642), .IN4(n2487), .IN5(
        n15580), .Q(n15575) );
  OA221X1 U23826 ( .IN1(n18657), .IN2(n2592), .IN3(n18655), .IN4(n2627), .IN5(
        n15579), .Q(n15576) );
  NAND4X0 U23827 ( .IN1(n15790), .IN2(n15791), .IN3(n15792), .IN4(n15793), 
        .QN(m3_rty_o) );
  OA221X1 U23828 ( .IN1(n8851), .IN2(n2346), .IN3(n8555), .IN4(n2696), .IN5(
        n15798), .Q(n15790) );
  OA221X1 U23829 ( .IN1(n6595), .IN2(n2416), .IN3(n6299), .IN4(n2451), .IN5(
        n15795), .Q(n15792) );
  OA221X1 U23830 ( .IN1(n4819), .IN2(n2626), .IN3(n4523), .IN4(n2661), .IN5(
        n15794), .Q(n15793) );
  NAND4X0 U23831 ( .IN1(n15799), .IN2(n15800), .IN3(n15801), .IN4(n15802), 
        .QN(m3_err_o) );
  OA221X1 U23832 ( .IN1(n8851), .IN2(n2345), .IN3(n8555), .IN4(n2695), .IN5(
        n15806), .Q(n15799) );
  OA221X1 U23833 ( .IN1(n6595), .IN2(n2415), .IN3(n6299), .IN4(n2450), .IN5(
        n15804), .Q(n15801) );
  OA221X1 U23834 ( .IN1(n4819), .IN2(n2625), .IN3(n4523), .IN4(n2660), .IN5(
        n15803), .Q(n15802) );
  NAND4X0 U23835 ( .IN1(n16079), .IN2(n16080), .IN3(n16081), .IN4(n16082), 
        .QN(m3_ack_o) );
  OA221X1 U23836 ( .IN1(n8851), .IN2(n2344), .IN3(n8555), .IN4(n2694), .IN5(
        n16094), .Q(n16079) );
  OA221X1 U23837 ( .IN1(n6595), .IN2(n2414), .IN3(n6299), .IN4(n2449), .IN5(
        n16090), .Q(n16081) );
  OA221X1 U23838 ( .IN1(n4819), .IN2(n2624), .IN3(n4523), .IN4(n2659), .IN5(
        n16083), .Q(n16082) );
  NAND4X0 U23839 ( .IN1(n16071), .IN2(n16072), .IN3(n16073), .IN4(n16074), 
        .QN(m3_data_o[0]) );
  OA221X1 U23840 ( .IN1(n18584), .IN2(n2413), .IN3(n18581), .IN4(n2448), .IN5(
        n16078), .Q(n16071) );
  OA221X1 U23841 ( .IN1(n18597), .IN2(n2483), .IN3(n18593), .IN4(n2518), .IN5(
        n16077), .Q(n16072) );
  OA221X1 U23842 ( .IN1(n18608), .IN2(n2623), .IN3(n18605), .IN4(n2658), .IN5(
        n16076), .Q(n16073) );
  NAND4X0 U23843 ( .IN1(n15983), .IN2(n15984), .IN3(n15985), .IN4(n15986), 
        .QN(m3_data_o[1]) );
  OA221X1 U23844 ( .IN1(n18586), .IN2(n2412), .IN3(n18582), .IN4(n2447), .IN5(
        n15990), .Q(n15983) );
  OA221X1 U23845 ( .IN1(n18596), .IN2(n2482), .IN3(n18593), .IN4(n2517), .IN5(
        n15989), .Q(n15984) );
  OA221X1 U23846 ( .IN1(n18609), .IN2(n2622), .IN3(n18605), .IN4(n2657), .IN5(
        n15988), .Q(n15985) );
  NAND4X0 U23847 ( .IN1(n15895), .IN2(n15896), .IN3(n15897), .IN4(n15898), 
        .QN(m3_data_o[2]) );
  OA221X1 U23848 ( .IN1(n18584), .IN2(n2411), .IN3(n18581), .IN4(n2446), .IN5(
        n15902), .Q(n15895) );
  OA221X1 U23849 ( .IN1(n18596), .IN2(n2481), .IN3(n18595), .IN4(n2516), .IN5(
        n15901), .Q(n15896) );
  OA221X1 U23850 ( .IN1(n18608), .IN2(n2621), .IN3(n18607), .IN4(n2656), .IN5(
        n15900), .Q(n15897) );
  NAND4X0 U23851 ( .IN1(n15871), .IN2(n15872), .IN3(n15873), .IN4(n15874), 
        .QN(m3_data_o[3]) );
  OA221X1 U23852 ( .IN1(n18585), .IN2(n2410), .IN3(n18583), .IN4(n2445), .IN5(
        n15878), .Q(n15871) );
  OA221X1 U23853 ( .IN1(n18598), .IN2(n2480), .IN3(n18594), .IN4(n2515), .IN5(
        n15877), .Q(n15872) );
  OA221X1 U23854 ( .IN1(n18610), .IN2(n2620), .IN3(n18606), .IN4(n2655), .IN5(
        n15876), .Q(n15873) );
  NAND4X0 U23855 ( .IN1(n15863), .IN2(n15864), .IN3(n15865), .IN4(n15866), 
        .QN(m3_data_o[4]) );
  OA221X1 U23856 ( .IN1(n18585), .IN2(n2409), .IN3(n18581), .IN4(n2444), .IN5(
        n15870), .Q(n15863) );
  OA221X1 U23857 ( .IN1(n18597), .IN2(n2479), .IN3(n18594), .IN4(n2514), .IN5(
        n15869), .Q(n15864) );
  OA221X1 U23858 ( .IN1(n18610), .IN2(n2619), .IN3(n18607), .IN4(n2654), .IN5(
        n15868), .Q(n15865) );
  NAND4X0 U23859 ( .IN1(n15855), .IN2(n15856), .IN3(n15857), .IN4(n15858), 
        .QN(m3_data_o[5]) );
  OA221X1 U23860 ( .IN1(n18584), .IN2(n2408), .IN3(n18582), .IN4(n2443), .IN5(
        n15862), .Q(n15855) );
  OA221X1 U23861 ( .IN1(n18598), .IN2(n2478), .IN3(n18594), .IN4(n2513), .IN5(
        n15861), .Q(n15856) );
  OA221X1 U23862 ( .IN1(n18609), .IN2(n2618), .IN3(n18607), .IN4(n2653), .IN5(
        n15860), .Q(n15857) );
  NAND4X0 U23863 ( .IN1(n15847), .IN2(n15848), .IN3(n15849), .IN4(n15850), 
        .QN(m3_data_o[6]) );
  OA221X1 U23864 ( .IN1(n18586), .IN2(n2407), .IN3(n18583), .IN4(n2442), .IN5(
        n15854), .Q(n15847) );
  OA221X1 U23865 ( .IN1(n18598), .IN2(n2477), .IN3(n18595), .IN4(n2512), .IN5(
        n15853), .Q(n15848) );
  OA221X1 U23866 ( .IN1(n18608), .IN2(n2617), .IN3(n18607), .IN4(n2652), .IN5(
        n15852), .Q(n15849) );
  NAND4X0 U23867 ( .IN1(n15839), .IN2(n15840), .IN3(n15841), .IN4(n15842), 
        .QN(m3_data_o[7]) );
  OA221X1 U23868 ( .IN1(n18586), .IN2(n2406), .IN3(n18583), .IN4(n2441), .IN5(
        n15846), .Q(n15839) );
  OA221X1 U23869 ( .IN1(n18598), .IN2(n2476), .IN3(n18595), .IN4(n2511), .IN5(
        n15845), .Q(n15840) );
  OA221X1 U23870 ( .IN1(n18608), .IN2(n2616), .IN3(n18607), .IN4(n2651), .IN5(
        n15844), .Q(n15841) );
  NAND4X0 U23871 ( .IN1(n15831), .IN2(n15832), .IN3(n15833), .IN4(n15834), 
        .QN(m3_data_o[8]) );
  OA221X1 U23872 ( .IN1(n18586), .IN2(n2405), .IN3(n18583), .IN4(n2440), .IN5(
        n15838), .Q(n15831) );
  OA221X1 U23873 ( .IN1(n18598), .IN2(n2475), .IN3(n18595), .IN4(n2510), .IN5(
        n15837), .Q(n15832) );
  OA221X1 U23874 ( .IN1(n18610), .IN2(n2615), .IN3(n18607), .IN4(n2650), .IN5(
        n15836), .Q(n15833) );
  NAND4X0 U23875 ( .IN1(n15807), .IN2(n15808), .IN3(n15809), .IN4(n15810), 
        .QN(m3_data_o[9]) );
  OA221X1 U23876 ( .IN1(n18586), .IN2(n2404), .IN3(n18583), .IN4(n2439), .IN5(
        n15828), .Q(n15807) );
  OA221X1 U23877 ( .IN1(n18598), .IN2(n2474), .IN3(n18595), .IN4(n2509), .IN5(
        n15823), .Q(n15808) );
  OA221X1 U23878 ( .IN1(n18609), .IN2(n2614), .IN3(n18607), .IN4(n2649), .IN5(
        n15818), .Q(n15809) );
  NAND4X0 U23879 ( .IN1(n16063), .IN2(n16064), .IN3(n16065), .IN4(n16066), 
        .QN(m3_data_o[10]) );
  OA221X1 U23880 ( .IN1(n18586), .IN2(n2403), .IN3(n18581), .IN4(n2438), .IN5(
        n16070), .Q(n16063) );
  OA221X1 U23881 ( .IN1(n18598), .IN2(n2473), .IN3(n18593), .IN4(n2508), .IN5(
        n16069), .Q(n16064) );
  OA221X1 U23882 ( .IN1(n18608), .IN2(n2613), .IN3(n18605), .IN4(n2648), .IN5(
        n16068), .Q(n16065) );
  NAND4X0 U23883 ( .IN1(n16055), .IN2(n16056), .IN3(n16057), .IN4(n16058), 
        .QN(m3_data_o[11]) );
  OA221X1 U23884 ( .IN1(n18585), .IN2(n2402), .IN3(n18581), .IN4(n2437), .IN5(
        n16062), .Q(n16055) );
  OA221X1 U23885 ( .IN1(n18596), .IN2(n2472), .IN3(n18593), .IN4(n2507), .IN5(
        n16061), .Q(n16056) );
  OA221X1 U23886 ( .IN1(n18608), .IN2(n2612), .IN3(n18605), .IN4(n2647), .IN5(
        n16060), .Q(n16057) );
  NAND4X0 U23887 ( .IN1(n16047), .IN2(n16048), .IN3(n16049), .IN4(n16050), 
        .QN(m3_data_o[12]) );
  OA221X1 U23888 ( .IN1(n18584), .IN2(n2401), .IN3(n18581), .IN4(n2436), .IN5(
        n16054), .Q(n16047) );
  OA221X1 U23889 ( .IN1(n18597), .IN2(n2471), .IN3(n18593), .IN4(n2506), .IN5(
        n16053), .Q(n16048) );
  OA221X1 U23890 ( .IN1(n18608), .IN2(n2611), .IN3(n18605), .IN4(n2646), .IN5(
        n16052), .Q(n16049) );
  NAND4X0 U23891 ( .IN1(n16039), .IN2(n16040), .IN3(n16041), .IN4(n16042), 
        .QN(m3_data_o[13]) );
  OA221X1 U23892 ( .IN1(n18584), .IN2(n2400), .IN3(n18582), .IN4(n2435), .IN5(
        n16046), .Q(n16039) );
  OA221X1 U23893 ( .IN1(n18598), .IN2(n2470), .IN3(n18595), .IN4(n2505), .IN5(
        n16045), .Q(n16040) );
  OA221X1 U23894 ( .IN1(n18608), .IN2(n2610), .IN3(n18606), .IN4(n2645), .IN5(
        n16044), .Q(n16041) );
  NAND4X0 U23895 ( .IN1(n16031), .IN2(n16032), .IN3(n16033), .IN4(n16034), 
        .QN(m3_data_o[14]) );
  OA221X1 U23896 ( .IN1(n18586), .IN2(n2399), .IN3(n18582), .IN4(n2434), .IN5(
        n16038), .Q(n16031) );
  OA221X1 U23897 ( .IN1(n18596), .IN2(n2469), .IN3(n18593), .IN4(n2504), .IN5(
        n16037), .Q(n16032) );
  OA221X1 U23898 ( .IN1(n18609), .IN2(n2609), .IN3(n18606), .IN4(n2644), .IN5(
        n16036), .Q(n16033) );
  NAND4X0 U23899 ( .IN1(n16023), .IN2(n16024), .IN3(n16025), .IN4(n16026), 
        .QN(m3_data_o[15]) );
  OA221X1 U23900 ( .IN1(n18585), .IN2(n2398), .IN3(n18582), .IN4(n2433), .IN5(
        n16030), .Q(n16023) );
  OA221X1 U23901 ( .IN1(n18596), .IN2(n2468), .IN3(n18594), .IN4(n2503), .IN5(
        n16029), .Q(n16024) );
  OA221X1 U23902 ( .IN1(n18608), .IN2(n2608), .IN3(n18606), .IN4(n2643), .IN5(
        n16028), .Q(n16025) );
  NAND4X0 U23903 ( .IN1(n16015), .IN2(n16016), .IN3(n16017), .IN4(n16018), 
        .QN(m3_data_o[16]) );
  OA221X1 U23904 ( .IN1(n18584), .IN2(n2397), .IN3(n18582), .IN4(n2432), .IN5(
        n16022), .Q(n16015) );
  OA221X1 U23905 ( .IN1(n18597), .IN2(n2467), .IN3(n18594), .IN4(n2502), .IN5(
        n16021), .Q(n16016) );
  OA221X1 U23906 ( .IN1(n18609), .IN2(n2607), .IN3(n18606), .IN4(n2642), .IN5(
        n16020), .Q(n16017) );
  NAND4X0 U23907 ( .IN1(n16007), .IN2(n16008), .IN3(n16009), .IN4(n16010), 
        .QN(m3_data_o[17]) );
  OA221X1 U23908 ( .IN1(n18585), .IN2(n2396), .IN3(n18583), .IN4(n2431), .IN5(
        n16014), .Q(n16007) );
  OA221X1 U23909 ( .IN1(n18598), .IN2(n2466), .IN3(n18595), .IN4(n2501), .IN5(
        n16013), .Q(n16008) );
  OA221X1 U23910 ( .IN1(n18609), .IN2(n2606), .IN3(n18606), .IN4(n2641), .IN5(
        n16012), .Q(n16009) );
  NAND4X0 U23911 ( .IN1(n15999), .IN2(n16000), .IN3(n16001), .IN4(n16002), 
        .QN(m3_data_o[18]) );
  OA221X1 U23912 ( .IN1(n18585), .IN2(n2395), .IN3(n18581), .IN4(n2430), .IN5(
        n16006), .Q(n15999) );
  OA221X1 U23913 ( .IN1(n18597), .IN2(n2465), .IN3(n18593), .IN4(n2500), .IN5(
        n16005), .Q(n16000) );
  OA221X1 U23914 ( .IN1(n18609), .IN2(n2605), .IN3(n18607), .IN4(n2640), .IN5(
        n16004), .Q(n16001) );
  NAND4X0 U23915 ( .IN1(n15991), .IN2(n15992), .IN3(n15993), .IN4(n15994), 
        .QN(m3_data_o[19]) );
  OA221X1 U23916 ( .IN1(n18586), .IN2(n2394), .IN3(n18582), .IN4(n2429), .IN5(
        n15998), .Q(n15991) );
  OA221X1 U23917 ( .IN1(n18596), .IN2(n2464), .IN3(n18593), .IN4(n2499), .IN5(
        n15997), .Q(n15992) );
  OA221X1 U23918 ( .IN1(n18609), .IN2(n2604), .IN3(n18605), .IN4(n2639), .IN5(
        n15996), .Q(n15993) );
  NAND4X0 U23919 ( .IN1(n15975), .IN2(n15976), .IN3(n15977), .IN4(n15978), 
        .QN(m3_data_o[20]) );
  OA221X1 U23920 ( .IN1(n18584), .IN2(n2393), .IN3(n18581), .IN4(n2428), .IN5(
        n15982), .Q(n15975) );
  OA221X1 U23921 ( .IN1(n18596), .IN2(n2463), .IN3(n18594), .IN4(n2498), .IN5(
        n15981), .Q(n15976) );
  OA221X1 U23922 ( .IN1(n18608), .IN2(n2603), .IN3(n18605), .IN4(n2638), .IN5(
        n15980), .Q(n15977) );
  NAND4X0 U23923 ( .IN1(n15967), .IN2(n15968), .IN3(n15969), .IN4(n15970), 
        .QN(m3_data_o[21]) );
  OA221X1 U23924 ( .IN1(n18584), .IN2(n2392), .IN3(n18582), .IN4(n2427), .IN5(
        n15974), .Q(n15967) );
  OA221X1 U23925 ( .IN1(n18596), .IN2(n2462), .IN3(n18594), .IN4(n2497), .IN5(
        n15973), .Q(n15968) );
  OA221X1 U23926 ( .IN1(n18609), .IN2(n2602), .IN3(n18606), .IN4(n2637), .IN5(
        n15972), .Q(n15969) );
  NAND4X0 U23927 ( .IN1(n15959), .IN2(n15960), .IN3(n15961), .IN4(n15962), 
        .QN(m3_data_o[22]) );
  OA221X1 U23928 ( .IN1(n18584), .IN2(n2391), .IN3(n18583), .IN4(n2426), .IN5(
        n15966), .Q(n15959) );
  OA221X1 U23929 ( .IN1(n18596), .IN2(n2461), .IN3(n18594), .IN4(n2496), .IN5(
        n15965), .Q(n15960) );
  OA221X1 U23930 ( .IN1(n18610), .IN2(n2601), .IN3(n18607), .IN4(n2636), .IN5(
        n15964), .Q(n15961) );
  NAND4X0 U23931 ( .IN1(n15951), .IN2(n15952), .IN3(n15953), .IN4(n15954), 
        .QN(m3_data_o[23]) );
  OA221X1 U23932 ( .IN1(n18584), .IN2(n2390), .IN3(n18581), .IN4(n2425), .IN5(
        n15958), .Q(n15951) );
  OA221X1 U23933 ( .IN1(n18596), .IN2(n2460), .IN3(n18594), .IN4(n2495), .IN5(
        n15957), .Q(n15952) );
  OA221X1 U23934 ( .IN1(n18610), .IN2(n2600), .IN3(n18605), .IN4(n2635), .IN5(
        n15956), .Q(n15953) );
  NAND4X0 U23935 ( .IN1(n15943), .IN2(n15944), .IN3(n15945), .IN4(n15946), 
        .QN(m3_data_o[24]) );
  OA221X1 U23936 ( .IN1(n18585), .IN2(n2389), .IN3(n18583), .IN4(n2424), .IN5(
        n15950), .Q(n15943) );
  OA221X1 U23937 ( .IN1(n18597), .IN2(n2459), .IN3(n18595), .IN4(n2494), .IN5(
        n15949), .Q(n15944) );
  OA221X1 U23938 ( .IN1(n18610), .IN2(n2599), .IN3(n18605), .IN4(n2634), .IN5(
        n15948), .Q(n15945) );
  NAND4X0 U23939 ( .IN1(n15935), .IN2(n15936), .IN3(n15937), .IN4(n15938), 
        .QN(m3_data_o[25]) );
  OA221X1 U23940 ( .IN1(n18585), .IN2(n2388), .IN3(n18583), .IN4(n2423), .IN5(
        n15942), .Q(n15935) );
  OA221X1 U23941 ( .IN1(n18597), .IN2(n2458), .IN3(n18593), .IN4(n2493), .IN5(
        n15941), .Q(n15936) );
  OA221X1 U23942 ( .IN1(n18610), .IN2(n2598), .IN3(n18606), .IN4(n2633), .IN5(
        n15940), .Q(n15937) );
  NAND4X0 U23943 ( .IN1(n15927), .IN2(n15928), .IN3(n15929), .IN4(n15930), 
        .QN(m3_data_o[26]) );
  OA221X1 U23944 ( .IN1(n18585), .IN2(n2387), .IN3(n18581), .IN4(n2422), .IN5(
        n15934), .Q(n15927) );
  OA221X1 U23945 ( .IN1(n18597), .IN2(n2457), .IN3(n18594), .IN4(n2492), .IN5(
        n15933), .Q(n15928) );
  OA221X1 U23946 ( .IN1(n18610), .IN2(n2597), .IN3(n18607), .IN4(n2632), .IN5(
        n15932), .Q(n15929) );
  NAND4X0 U23947 ( .IN1(n15919), .IN2(n15920), .IN3(n15921), .IN4(n15922), 
        .QN(m3_data_o[27]) );
  OA221X1 U23948 ( .IN1(n18585), .IN2(n2386), .IN3(n18582), .IN4(n2421), .IN5(
        n15926), .Q(n15919) );
  OA221X1 U23949 ( .IN1(n18597), .IN2(n2456), .IN3(n18595), .IN4(n2491), .IN5(
        n15925), .Q(n15920) );
  OA221X1 U23950 ( .IN1(n18610), .IN2(n2596), .IN3(n18605), .IN4(n2631), .IN5(
        n15924), .Q(n15921) );
  NAND4X0 U23951 ( .IN1(n15911), .IN2(n15912), .IN3(n15913), .IN4(n15914), 
        .QN(m3_data_o[28]) );
  OA221X1 U23952 ( .IN1(n18586), .IN2(n2385), .IN3(n18582), .IN4(n2420), .IN5(
        n15918), .Q(n15911) );
  OA221X1 U23953 ( .IN1(n18597), .IN2(n2455), .IN3(n18595), .IN4(n2490), .IN5(
        n15917), .Q(n15912) );
  OA221X1 U23954 ( .IN1(n18609), .IN2(n2595), .IN3(n18605), .IN4(n2630), .IN5(
        n15916), .Q(n15913) );
  NAND4X0 U23955 ( .IN1(n15903), .IN2(n15904), .IN3(n15905), .IN4(n15906), 
        .QN(m3_data_o[29]) );
  OA221X1 U23956 ( .IN1(n18585), .IN2(n2384), .IN3(n18583), .IN4(n2419), .IN5(
        n15910), .Q(n15903) );
  OA221X1 U23957 ( .IN1(n18597), .IN2(n2454), .IN3(n18594), .IN4(n2489), .IN5(
        n15909), .Q(n15904) );
  OA221X1 U23958 ( .IN1(n18608), .IN2(n2594), .IN3(n18606), .IN4(n2629), .IN5(
        n15908), .Q(n15905) );
  NAND4X0 U23959 ( .IN1(n15887), .IN2(n15888), .IN3(n15889), .IN4(n15890), 
        .QN(m3_data_o[30]) );
  OA221X1 U23960 ( .IN1(n18584), .IN2(n2383), .IN3(n18581), .IN4(n2418), .IN5(
        n15894), .Q(n15887) );
  OA221X1 U23961 ( .IN1(n18598), .IN2(n2453), .IN3(n18593), .IN4(n2488), .IN5(
        n15893), .Q(n15888) );
  OA221X1 U23962 ( .IN1(n18610), .IN2(n2593), .IN3(n18607), .IN4(n2628), .IN5(
        n15892), .Q(n15889) );
  NAND4X0 U23963 ( .IN1(n15879), .IN2(n15880), .IN3(n15881), .IN4(n15882), 
        .QN(m3_data_o[31]) );
  OA221X1 U23964 ( .IN1(n18586), .IN2(n2382), .IN3(n18583), .IN4(n2417), .IN5(
        n15886), .Q(n15879) );
  OA221X1 U23965 ( .IN1(n18596), .IN2(n2452), .IN3(n18595), .IN4(n2487), .IN5(
        n15885), .Q(n15880) );
  OA221X1 U23966 ( .IN1(n18610), .IN2(n2592), .IN3(n18606), .IN4(n2627), .IN5(
        n15884), .Q(n15881) );
  NAND4X0 U23967 ( .IN1(n16095), .IN2(n16096), .IN3(n16097), .IN4(n16098), 
        .QN(m2_rty_o) );
  OA221X1 U23968 ( .IN1(n8852), .IN2(n2346), .IN3(n8556), .IN4(n2696), .IN5(
        n16103), .Q(n16095) );
  OA221X1 U23969 ( .IN1(n6596), .IN2(n2416), .IN3(n6300), .IN4(n2451), .IN5(
        n16100), .Q(n16097) );
  OA221X1 U23970 ( .IN1(n4820), .IN2(n2626), .IN3(n4524), .IN4(n2661), .IN5(
        n16099), .Q(n16098) );
  NAND4X0 U23971 ( .IN1(n16104), .IN2(n16105), .IN3(n16106), .IN4(n16107), 
        .QN(m2_err_o) );
  OA221X1 U23972 ( .IN1(n8852), .IN2(n2345), .IN3(n8556), .IN4(n2695), .IN5(
        n16111), .Q(n16104) );
  OA221X1 U23973 ( .IN1(n6596), .IN2(n2415), .IN3(n6300), .IN4(n2450), .IN5(
        n16109), .Q(n16106) );
  OA221X1 U23974 ( .IN1(n4820), .IN2(n2625), .IN3(n4524), .IN4(n2660), .IN5(
        n16108), .Q(n16107) );
  NAND4X0 U23975 ( .IN1(n16384), .IN2(n16385), .IN3(n16386), .IN4(n16387), 
        .QN(m2_ack_o) );
  OA221X1 U23976 ( .IN1(n8852), .IN2(n2344), .IN3(n8556), .IN4(n2694), .IN5(
        n16399), .Q(n16384) );
  OA221X1 U23977 ( .IN1(n6596), .IN2(n2414), .IN3(n6300), .IN4(n2449), .IN5(
        n16395), .Q(n16386) );
  OA221X1 U23978 ( .IN1(n4820), .IN2(n2624), .IN3(n4524), .IN4(n2659), .IN5(
        n16388), .Q(n16387) );
  NAND4X0 U23979 ( .IN1(n16376), .IN2(n16377), .IN3(n16378), .IN4(n16379), 
        .QN(m2_data_o[0]) );
  OA221X1 U23980 ( .IN1(n18536), .IN2(n2413), .IN3(n16132), .IN4(n2448), .IN5(
        n16383), .Q(n16376) );
  OA221X1 U23981 ( .IN1(n18548), .IN2(n2483), .IN3(n18545), .IN4(n2518), .IN5(
        n16382), .Q(n16377) );
  OA221X1 U23982 ( .IN1(n18561), .IN2(n2623), .IN3(n18557), .IN4(n2658), .IN5(
        n16381), .Q(n16378) );
  NAND4X0 U23983 ( .IN1(n16288), .IN2(n16289), .IN3(n16290), .IN4(n16291), 
        .QN(m2_data_o[1]) );
  OA221X1 U23984 ( .IN1(n18538), .IN2(n2412), .IN3(n18534), .IN4(n2447), .IN5(
        n16295), .Q(n16288) );
  OA221X1 U23985 ( .IN1(n18550), .IN2(n2482), .IN3(n18545), .IN4(n2517), .IN5(
        n16294), .Q(n16289) );
  OA221X1 U23986 ( .IN1(n18562), .IN2(n2622), .IN3(n18557), .IN4(n2657), .IN5(
        n16293), .Q(n16290) );
  NAND4X0 U23987 ( .IN1(n16200), .IN2(n16201), .IN3(n16202), .IN4(n16203), 
        .QN(m2_data_o[2]) );
  OA221X1 U23988 ( .IN1(n18536), .IN2(n2411), .IN3(n18534), .IN4(n2446), .IN5(
        n16207), .Q(n16200) );
  OA221X1 U23989 ( .IN1(n18550), .IN2(n2481), .IN3(n18547), .IN4(n2516), .IN5(
        n16206), .Q(n16201) );
  OA221X1 U23990 ( .IN1(n18562), .IN2(n2621), .IN3(n18558), .IN4(n2656), .IN5(
        n16205), .Q(n16202) );
  NAND4X0 U23991 ( .IN1(n16176), .IN2(n16177), .IN3(n16178), .IN4(n16179), 
        .QN(m2_data_o[3]) );
  OA221X1 U23992 ( .IN1(n18538), .IN2(n2410), .IN3(n18534), .IN4(n2445), .IN5(
        n16183), .Q(n16176) );
  OA221X1 U23993 ( .IN1(n18550), .IN2(n2480), .IN3(n18546), .IN4(n2515), .IN5(
        n16182), .Q(n16177) );
  OA221X1 U23994 ( .IN1(n18562), .IN2(n2620), .IN3(n18558), .IN4(n2655), .IN5(
        n16181), .Q(n16178) );
  NAND4X0 U23995 ( .IN1(n16168), .IN2(n16169), .IN3(n16170), .IN4(n16171), 
        .QN(m2_data_o[4]) );
  OA221X1 U23996 ( .IN1(n18536), .IN2(n2409), .IN3(n18533), .IN4(n2444), .IN5(
        n16175), .Q(n16168) );
  OA221X1 U23997 ( .IN1(n18548), .IN2(n2479), .IN3(n18547), .IN4(n2514), .IN5(
        n16174), .Q(n16169) );
  OA221X1 U23998 ( .IN1(n18561), .IN2(n2619), .IN3(n18559), .IN4(n2654), .IN5(
        n16173), .Q(n16170) );
  NAND4X0 U23999 ( .IN1(n16160), .IN2(n16161), .IN3(n16162), .IN4(n16163), 
        .QN(m2_data_o[5]) );
  OA221X1 U24000 ( .IN1(n18537), .IN2(n2408), .IN3(n16132), .IN4(n2443), .IN5(
        n16167), .Q(n16160) );
  OA221X1 U24001 ( .IN1(n18549), .IN2(n2478), .IN3(n18547), .IN4(n2513), .IN5(
        n16166), .Q(n16161) );
  OA221X1 U24002 ( .IN1(n18560), .IN2(n2618), .IN3(n18558), .IN4(n2653), .IN5(
        n16165), .Q(n16162) );
  NAND4X0 U24003 ( .IN1(n16152), .IN2(n16153), .IN3(n16154), .IN4(n16155), 
        .QN(m2_data_o[6]) );
  OA221X1 U24004 ( .IN1(n18538), .IN2(n2407), .IN3(n18534), .IN4(n2442), .IN5(
        n16159), .Q(n16152) );
  OA221X1 U24005 ( .IN1(n18550), .IN2(n2477), .IN3(n18547), .IN4(n2512), .IN5(
        n16158), .Q(n16153) );
  OA221X1 U24006 ( .IN1(n18562), .IN2(n2617), .IN3(n18559), .IN4(n2652), .IN5(
        n16157), .Q(n16154) );
  NAND4X0 U24007 ( .IN1(n16144), .IN2(n16145), .IN3(n16146), .IN4(n16147), 
        .QN(m2_data_o[7]) );
  OA221X1 U24008 ( .IN1(n18538), .IN2(n2406), .IN3(n18534), .IN4(n2441), .IN5(
        n16151), .Q(n16144) );
  OA221X1 U24009 ( .IN1(n18550), .IN2(n2476), .IN3(n18547), .IN4(n2511), .IN5(
        n16150), .Q(n16145) );
  OA221X1 U24010 ( .IN1(n18562), .IN2(n2616), .IN3(n18559), .IN4(n2651), .IN5(
        n16149), .Q(n16146) );
  NAND4X0 U24011 ( .IN1(n16136), .IN2(n16137), .IN3(n16138), .IN4(n16139), 
        .QN(m2_data_o[8]) );
  OA221X1 U24012 ( .IN1(n18538), .IN2(n2405), .IN3(n18534), .IN4(n2440), .IN5(
        n16143), .Q(n16136) );
  OA221X1 U24013 ( .IN1(n18550), .IN2(n2475), .IN3(n18547), .IN4(n2510), .IN5(
        n16142), .Q(n16137) );
  OA221X1 U24014 ( .IN1(n18562), .IN2(n2615), .IN3(n18559), .IN4(n2650), .IN5(
        n16141), .Q(n16138) );
  NAND4X0 U24015 ( .IN1(n16112), .IN2(n16113), .IN3(n16114), .IN4(n16115), 
        .QN(m2_data_o[9]) );
  OA221X1 U24016 ( .IN1(n18538), .IN2(n2404), .IN3(n18534), .IN4(n2439), .IN5(
        n16133), .Q(n16112) );
  OA221X1 U24017 ( .IN1(n18550), .IN2(n2474), .IN3(n18547), .IN4(n2509), .IN5(
        n16128), .Q(n16113) );
  OA221X1 U24018 ( .IN1(n18562), .IN2(n2614), .IN3(n18559), .IN4(n2649), .IN5(
        n16123), .Q(n16114) );
  NAND4X0 U24019 ( .IN1(n16368), .IN2(n16369), .IN3(n16370), .IN4(n16371), 
        .QN(m2_data_o[10]) );
  OA221X1 U24020 ( .IN1(n18537), .IN2(n2403), .IN3(n16132), .IN4(n2438), .IN5(
        n16375), .Q(n16368) );
  OA221X1 U24021 ( .IN1(n18550), .IN2(n2473), .IN3(n18545), .IN4(n2508), .IN5(
        n16374), .Q(n16369) );
  OA221X1 U24022 ( .IN1(n18560), .IN2(n2613), .IN3(n18557), .IN4(n2648), .IN5(
        n16373), .Q(n16370) );
  NAND4X0 U24023 ( .IN1(n16360), .IN2(n16361), .IN3(n16362), .IN4(n16363), 
        .QN(m2_data_o[11]) );
  OA221X1 U24024 ( .IN1(n18536), .IN2(n2402), .IN3(n16132), .IN4(n2437), .IN5(
        n16367), .Q(n16360) );
  OA221X1 U24025 ( .IN1(n18548), .IN2(n2472), .IN3(n18545), .IN4(n2507), .IN5(
        n16366), .Q(n16361) );
  OA221X1 U24026 ( .IN1(n18562), .IN2(n2612), .IN3(n18557), .IN4(n2647), .IN5(
        n16365), .Q(n16362) );
  NAND4X0 U24027 ( .IN1(n16352), .IN2(n16353), .IN3(n16354), .IN4(n16355), 
        .QN(m2_data_o[12]) );
  OA221X1 U24028 ( .IN1(n18537), .IN2(n2401), .IN3(n16132), .IN4(n2436), .IN5(
        n16359), .Q(n16352) );
  OA221X1 U24029 ( .IN1(n18549), .IN2(n2471), .IN3(n18545), .IN4(n2506), .IN5(
        n16358), .Q(n16353) );
  OA221X1 U24030 ( .IN1(n18561), .IN2(n2611), .IN3(n18557), .IN4(n2646), .IN5(
        n16357), .Q(n16354) );
  NAND4X0 U24031 ( .IN1(n16344), .IN2(n16345), .IN3(n16346), .IN4(n16347), 
        .QN(m2_data_o[13]) );
  OA221X1 U24032 ( .IN1(n18536), .IN2(n2400), .IN3(n18533), .IN4(n2435), .IN5(
        n16351), .Q(n16344) );
  OA221X1 U24033 ( .IN1(n18548), .IN2(n2470), .IN3(n18546), .IN4(n2505), .IN5(
        n16350), .Q(n16345) );
  OA221X1 U24034 ( .IN1(n18560), .IN2(n2610), .IN3(n18559), .IN4(n2645), .IN5(
        n16349), .Q(n16346) );
  NAND4X0 U24035 ( .IN1(n16336), .IN2(n16337), .IN3(n16338), .IN4(n16339), 
        .QN(m2_data_o[14]) );
  OA221X1 U24036 ( .IN1(n18536), .IN2(n2399), .IN3(n18533), .IN4(n2434), .IN5(
        n16343), .Q(n16336) );
  OA221X1 U24037 ( .IN1(n18548), .IN2(n2469), .IN3(n18546), .IN4(n2504), .IN5(
        n16342), .Q(n16337) );
  OA221X1 U24038 ( .IN1(n18560), .IN2(n2609), .IN3(n18557), .IN4(n2644), .IN5(
        n16341), .Q(n16338) );
  NAND4X0 U24039 ( .IN1(n16328), .IN2(n16329), .IN3(n16330), .IN4(n16331), 
        .QN(m2_data_o[15]) );
  OA221X1 U24040 ( .IN1(n18536), .IN2(n2398), .IN3(n18533), .IN4(n2433), .IN5(
        n16335), .Q(n16328) );
  OA221X1 U24041 ( .IN1(n18548), .IN2(n2468), .IN3(n18546), .IN4(n2503), .IN5(
        n16334), .Q(n16329) );
  OA221X1 U24042 ( .IN1(n18560), .IN2(n2608), .IN3(n18558), .IN4(n2643), .IN5(
        n16333), .Q(n16330) );
  NAND4X0 U24043 ( .IN1(n16320), .IN2(n16321), .IN3(n16322), .IN4(n16323), 
        .QN(m2_data_o[16]) );
  OA221X1 U24044 ( .IN1(n18536), .IN2(n2397), .IN3(n18533), .IN4(n2432), .IN5(
        n16327), .Q(n16320) );
  OA221X1 U24045 ( .IN1(n18548), .IN2(n2467), .IN3(n18546), .IN4(n2502), .IN5(
        n16326), .Q(n16321) );
  OA221X1 U24046 ( .IN1(n18560), .IN2(n2607), .IN3(n18558), .IN4(n2642), .IN5(
        n16325), .Q(n16322) );
  NAND4X0 U24047 ( .IN1(n16312), .IN2(n16313), .IN3(n16314), .IN4(n16315), 
        .QN(m2_data_o[17]) );
  OA221X1 U24048 ( .IN1(n18537), .IN2(n2396), .IN3(n18533), .IN4(n2431), .IN5(
        n16319), .Q(n16312) );
  OA221X1 U24049 ( .IN1(n18549), .IN2(n2466), .IN3(n18546), .IN4(n2501), .IN5(
        n16318), .Q(n16313) );
  OA221X1 U24050 ( .IN1(n18560), .IN2(n2606), .IN3(n18559), .IN4(n2641), .IN5(
        n16317), .Q(n16314) );
  NAND4X0 U24051 ( .IN1(n16304), .IN2(n16305), .IN3(n16306), .IN4(n16307), 
        .QN(m2_data_o[18]) );
  OA221X1 U24052 ( .IN1(n18537), .IN2(n2395), .IN3(n18534), .IN4(n2430), .IN5(
        n16311), .Q(n16304) );
  OA221X1 U24053 ( .IN1(n18549), .IN2(n2465), .IN3(n18547), .IN4(n2500), .IN5(
        n16310), .Q(n16305) );
  OA221X1 U24054 ( .IN1(n18561), .IN2(n2605), .IN3(n18557), .IN4(n2640), .IN5(
        n16309), .Q(n16306) );
  NAND4X0 U24055 ( .IN1(n16296), .IN2(n16297), .IN3(n16298), .IN4(n16299), 
        .QN(m2_data_o[19]) );
  OA221X1 U24056 ( .IN1(n18536), .IN2(n2394), .IN3(n18534), .IN4(n2429), .IN5(
        n16303), .Q(n16296) );
  OA221X1 U24057 ( .IN1(n18548), .IN2(n2464), .IN3(n18545), .IN4(n2499), .IN5(
        n16302), .Q(n16297) );
  OA221X1 U24058 ( .IN1(n18562), .IN2(n2604), .IN3(n18557), .IN4(n2639), .IN5(
        n16301), .Q(n16298) );
  NAND4X0 U24059 ( .IN1(n16280), .IN2(n16281), .IN3(n16282), .IN4(n16283), 
        .QN(m2_data_o[20]) );
  OA221X1 U24060 ( .IN1(n18537), .IN2(n2393), .IN3(n16132), .IN4(n2428), .IN5(
        n16287), .Q(n16280) );
  OA221X1 U24061 ( .IN1(n18549), .IN2(n2463), .IN3(n18545), .IN4(n2498), .IN5(
        n16286), .Q(n16281) );
  OA221X1 U24062 ( .IN1(n18560), .IN2(n2603), .IN3(n18558), .IN4(n2638), .IN5(
        n16285), .Q(n16282) );
  NAND4X0 U24063 ( .IN1(n16272), .IN2(n16273), .IN3(n16274), .IN4(n16275), 
        .QN(m2_data_o[21]) );
  OA221X1 U24064 ( .IN1(n18537), .IN2(n2392), .IN3(n16132), .IN4(n2427), .IN5(
        n16279), .Q(n16272) );
  OA221X1 U24065 ( .IN1(n18549), .IN2(n2462), .IN3(n18546), .IN4(n2497), .IN5(
        n16278), .Q(n16273) );
  OA221X1 U24066 ( .IN1(n18560), .IN2(n2602), .IN3(n18558), .IN4(n2637), .IN5(
        n16277), .Q(n16274) );
  NAND4X0 U24067 ( .IN1(n16264), .IN2(n16265), .IN3(n16266), .IN4(n16267), 
        .QN(m2_data_o[22]) );
  OA221X1 U24068 ( .IN1(n18537), .IN2(n2391), .IN3(n16132), .IN4(n2426), .IN5(
        n16271), .Q(n16264) );
  OA221X1 U24069 ( .IN1(n18549), .IN2(n2461), .IN3(n18547), .IN4(n2496), .IN5(
        n16270), .Q(n16265) );
  OA221X1 U24070 ( .IN1(n18561), .IN2(n2601), .IN3(n18558), .IN4(n2636), .IN5(
        n16269), .Q(n16266) );
  NAND4X0 U24071 ( .IN1(n16256), .IN2(n16257), .IN3(n16258), .IN4(n16259), 
        .QN(m2_data_o[23]) );
  OA221X1 U24072 ( .IN1(n18537), .IN2(n2390), .IN3(n16132), .IN4(n2425), .IN5(
        n16263), .Q(n16256) );
  OA221X1 U24073 ( .IN1(n18549), .IN2(n2460), .IN3(n18545), .IN4(n2495), .IN5(
        n16262), .Q(n16257) );
  OA221X1 U24074 ( .IN1(n18562), .IN2(n2600), .IN3(n18558), .IN4(n2635), .IN5(
        n16261), .Q(n16258) );
  NAND4X0 U24075 ( .IN1(n16248), .IN2(n16249), .IN3(n16250), .IN4(n16251), 
        .QN(m2_data_o[24]) );
  OA221X1 U24076 ( .IN1(n18537), .IN2(n2389), .IN3(n18533), .IN4(n2424), .IN5(
        n16255), .Q(n16248) );
  OA221X1 U24077 ( .IN1(n18549), .IN2(n2459), .IN3(n18545), .IN4(n2494), .IN5(
        n16254), .Q(n16249) );
  OA221X1 U24078 ( .IN1(n18561), .IN2(n2599), .IN3(n18559), .IN4(n2634), .IN5(
        n16253), .Q(n16250) );
  NAND4X0 U24079 ( .IN1(n16240), .IN2(n16241), .IN3(n16242), .IN4(n16243), 
        .QN(m2_data_o[25]) );
  OA221X1 U24080 ( .IN1(n18538), .IN2(n2388), .IN3(n18533), .IN4(n2423), .IN5(
        n16247), .Q(n16240) );
  OA221X1 U24081 ( .IN1(n18550), .IN2(n2458), .IN3(n18546), .IN4(n2493), .IN5(
        n16246), .Q(n16241) );
  OA221X1 U24082 ( .IN1(n18561), .IN2(n2598), .IN3(n18557), .IN4(n2633), .IN5(
        n16245), .Q(n16242) );
  NAND4X0 U24083 ( .IN1(n16232), .IN2(n16233), .IN3(n16234), .IN4(n16235), 
        .QN(m2_data_o[26]) );
  OA221X1 U24084 ( .IN1(n18537), .IN2(n2387), .IN3(n16132), .IN4(n2422), .IN5(
        n16239), .Q(n16232) );
  OA221X1 U24085 ( .IN1(n18549), .IN2(n2457), .IN3(n18547), .IN4(n2492), .IN5(
        n16238), .Q(n16233) );
  OA221X1 U24086 ( .IN1(n18561), .IN2(n2597), .IN3(n18558), .IN4(n2632), .IN5(
        n16237), .Q(n16234) );
  NAND4X0 U24087 ( .IN1(n16224), .IN2(n16225), .IN3(n16226), .IN4(n16227), 
        .QN(m2_data_o[27]) );
  OA221X1 U24088 ( .IN1(n18536), .IN2(n2386), .IN3(n16132), .IN4(n2421), .IN5(
        n16231), .Q(n16224) );
  OA221X1 U24089 ( .IN1(n18548), .IN2(n2456), .IN3(n18545), .IN4(n2491), .IN5(
        n16230), .Q(n16225) );
  OA221X1 U24090 ( .IN1(n18561), .IN2(n2596), .IN3(n18559), .IN4(n2631), .IN5(
        n16229), .Q(n16226) );
  NAND4X0 U24091 ( .IN1(n16216), .IN2(n16217), .IN3(n16218), .IN4(n16219), 
        .QN(m2_data_o[28]) );
  OA221X1 U24092 ( .IN1(n18538), .IN2(n2385), .IN3(n16132), .IN4(n2420), .IN5(
        n16223), .Q(n16216) );
  OA221X1 U24093 ( .IN1(n18548), .IN2(n2455), .IN3(n18545), .IN4(n2490), .IN5(
        n16222), .Q(n16217) );
  OA221X1 U24094 ( .IN1(n18562), .IN2(n2595), .IN3(n18559), .IN4(n2630), .IN5(
        n16221), .Q(n16218) );
  NAND4X0 U24095 ( .IN1(n16208), .IN2(n16209), .IN3(n16210), .IN4(n16211), 
        .QN(m2_data_o[29]) );
  OA221X1 U24096 ( .IN1(n18536), .IN2(n2384), .IN3(n18533), .IN4(n2419), .IN5(
        n16215), .Q(n16208) );
  OA221X1 U24097 ( .IN1(n18549), .IN2(n2454), .IN3(n18546), .IN4(n2489), .IN5(
        n16214), .Q(n16209) );
  OA221X1 U24098 ( .IN1(n18560), .IN2(n2594), .IN3(n18557), .IN4(n2629), .IN5(
        n16213), .Q(n16210) );
  NAND4X0 U24099 ( .IN1(n16192), .IN2(n16193), .IN3(n16194), .IN4(n16195), 
        .QN(m2_data_o[30]) );
  OA221X1 U24100 ( .IN1(n18538), .IN2(n2383), .IN3(n18534), .IN4(n2418), .IN5(
        n16199), .Q(n16192) );
  OA221X1 U24101 ( .IN1(n18550), .IN2(n2453), .IN3(n18547), .IN4(n2488), .IN5(
        n16198), .Q(n16193) );
  OA221X1 U24102 ( .IN1(n18561), .IN2(n2593), .IN3(n18558), .IN4(n2628), .IN5(
        n16197), .Q(n16194) );
  NAND4X0 U24103 ( .IN1(n16184), .IN2(n16185), .IN3(n16186), .IN4(n16187), 
        .QN(m2_data_o[31]) );
  OA221X1 U24104 ( .IN1(n18538), .IN2(n2382), .IN3(n18533), .IN4(n2417), .IN5(
        n16191), .Q(n16184) );
  OA221X1 U24105 ( .IN1(n18550), .IN2(n2452), .IN3(n18546), .IN4(n2487), .IN5(
        n16190), .Q(n16185) );
  OA221X1 U24106 ( .IN1(n18561), .IN2(n2592), .IN3(n18559), .IN4(n2627), .IN5(
        n16189), .Q(n16186) );
  NAND4X0 U24107 ( .IN1(n16400), .IN2(n16401), .IN3(n16402), .IN4(n16403), 
        .QN(m1_rty_o) );
  OA221X1 U24108 ( .IN1(n8853), .IN2(n2346), .IN3(n8557), .IN4(n2696), .IN5(
        n16408), .Q(n16400) );
  OA221X1 U24109 ( .IN1(n6597), .IN2(n2416), .IN3(n6301), .IN4(n2451), .IN5(
        n16405), .Q(n16402) );
  OA221X1 U24110 ( .IN1(n4821), .IN2(n2626), .IN3(n4525), .IN4(n2661), .IN5(
        n16404), .Q(n16403) );
  NAND4X0 U24111 ( .IN1(n16409), .IN2(n16410), .IN3(n16411), .IN4(n16412), 
        .QN(m1_err_o) );
  OA221X1 U24112 ( .IN1(n8853), .IN2(n2345), .IN3(n8557), .IN4(n2695), .IN5(
        n16416), .Q(n16409) );
  OA221X1 U24113 ( .IN1(n6597), .IN2(n2415), .IN3(n6301), .IN4(n2450), .IN5(
        n16414), .Q(n16411) );
  OA221X1 U24114 ( .IN1(n4821), .IN2(n2625), .IN3(n4525), .IN4(n2660), .IN5(
        n16413), .Q(n16412) );
  NAND4X0 U24115 ( .IN1(n16689), .IN2(n16690), .IN3(n16691), .IN4(n16692), 
        .QN(m1_ack_o) );
  OA221X1 U24116 ( .IN1(n8853), .IN2(n2344), .IN3(n8557), .IN4(n2694), .IN5(
        n16704), .Q(n16689) );
  OA221X1 U24117 ( .IN1(n6597), .IN2(n2414), .IN3(n6301), .IN4(n2449), .IN5(
        n16700), .Q(n16691) );
  OA221X1 U24118 ( .IN1(n4821), .IN2(n2624), .IN3(n4525), .IN4(n2659), .IN5(
        n16693), .Q(n16692) );
  NAND4X0 U24119 ( .IN1(n16681), .IN2(n16682), .IN3(n16683), .IN4(n16684), 
        .QN(m1_data_o[0]) );
  OA221X1 U24120 ( .IN1(n18488), .IN2(n2413), .IN3(n18485), .IN4(n2448), .IN5(
        n16688), .Q(n16681) );
  OA221X1 U24121 ( .IN1(n18501), .IN2(n2483), .IN3(n18497), .IN4(n2518), .IN5(
        n16687), .Q(n16682) );
  OA221X1 U24122 ( .IN1(n18512), .IN2(n2623), .IN3(n18509), .IN4(n2658), .IN5(
        n16686), .Q(n16683) );
  NAND4X0 U24123 ( .IN1(n16593), .IN2(n16594), .IN3(n16595), .IN4(n16596), 
        .QN(m1_data_o[1]) );
  OA221X1 U24124 ( .IN1(n18490), .IN2(n2412), .IN3(n18486), .IN4(n2447), .IN5(
        n16600), .Q(n16593) );
  OA221X1 U24125 ( .IN1(n18500), .IN2(n2482), .IN3(n18497), .IN4(n2517), .IN5(
        n16599), .Q(n16594) );
  OA221X1 U24126 ( .IN1(n18514), .IN2(n2622), .IN3(n18509), .IN4(n2657), .IN5(
        n16598), .Q(n16595) );
  NAND4X0 U24127 ( .IN1(n16505), .IN2(n16506), .IN3(n16507), .IN4(n16508), 
        .QN(m1_data_o[2]) );
  OA221X1 U24128 ( .IN1(n18488), .IN2(n2411), .IN3(n18485), .IN4(n2446), .IN5(
        n16512), .Q(n16505) );
  OA221X1 U24129 ( .IN1(n18500), .IN2(n2481), .IN3(n18499), .IN4(n2516), .IN5(
        n16511), .Q(n16506) );
  OA221X1 U24130 ( .IN1(n18513), .IN2(n2621), .IN3(n18511), .IN4(n2656), .IN5(
        n16510), .Q(n16507) );
  NAND4X0 U24131 ( .IN1(n16481), .IN2(n16482), .IN3(n16483), .IN4(n16484), 
        .QN(m1_data_o[3]) );
  OA221X1 U24132 ( .IN1(n18489), .IN2(n2410), .IN3(n18487), .IN4(n2445), .IN5(
        n16488), .Q(n16481) );
  OA221X1 U24133 ( .IN1(n18502), .IN2(n2480), .IN3(n18498), .IN4(n2515), .IN5(
        n16487), .Q(n16482) );
  OA221X1 U24134 ( .IN1(n18513), .IN2(n2620), .IN3(n18510), .IN4(n2655), .IN5(
        n16486), .Q(n16483) );
  NAND4X0 U24135 ( .IN1(n16473), .IN2(n16474), .IN3(n16475), .IN4(n16476), 
        .QN(m1_data_o[4]) );
  OA221X1 U24136 ( .IN1(n18489), .IN2(n2409), .IN3(n18485), .IN4(n2444), .IN5(
        n16480), .Q(n16473) );
  OA221X1 U24137 ( .IN1(n18501), .IN2(n2479), .IN3(n18498), .IN4(n2514), .IN5(
        n16479), .Q(n16474) );
  OA221X1 U24138 ( .IN1(n18513), .IN2(n2619), .IN3(n18511), .IN4(n2654), .IN5(
        n16478), .Q(n16475) );
  NAND4X0 U24139 ( .IN1(n16465), .IN2(n16466), .IN3(n16467), .IN4(n16468), 
        .QN(m1_data_o[5]) );
  OA221X1 U24140 ( .IN1(n18488), .IN2(n2408), .IN3(n18486), .IN4(n2443), .IN5(
        n16472), .Q(n16465) );
  OA221X1 U24141 ( .IN1(n18502), .IN2(n2478), .IN3(n18498), .IN4(n2513), .IN5(
        n16471), .Q(n16466) );
  OA221X1 U24142 ( .IN1(n18512), .IN2(n2618), .IN3(n18511), .IN4(n2653), .IN5(
        n16470), .Q(n16467) );
  NAND4X0 U24143 ( .IN1(n16457), .IN2(n16458), .IN3(n16459), .IN4(n16460), 
        .QN(m1_data_o[6]) );
  OA221X1 U24144 ( .IN1(n18490), .IN2(n2407), .IN3(n18487), .IN4(n2442), .IN5(
        n16464), .Q(n16457) );
  OA221X1 U24145 ( .IN1(n18502), .IN2(n2477), .IN3(n18499), .IN4(n2512), .IN5(
        n16463), .Q(n16458) );
  OA221X1 U24146 ( .IN1(n18514), .IN2(n2617), .IN3(n18511), .IN4(n2652), .IN5(
        n16462), .Q(n16459) );
  NAND4X0 U24147 ( .IN1(n16449), .IN2(n16450), .IN3(n16451), .IN4(n16452), 
        .QN(m1_data_o[7]) );
  OA221X1 U24148 ( .IN1(n18490), .IN2(n2406), .IN3(n18487), .IN4(n2441), .IN5(
        n16456), .Q(n16449) );
  OA221X1 U24149 ( .IN1(n18502), .IN2(n2476), .IN3(n18499), .IN4(n2511), .IN5(
        n16455), .Q(n16450) );
  OA221X1 U24150 ( .IN1(n18514), .IN2(n2616), .IN3(n18511), .IN4(n2651), .IN5(
        n16454), .Q(n16451) );
  NAND4X0 U24151 ( .IN1(n16441), .IN2(n16442), .IN3(n16443), .IN4(n16444), 
        .QN(m1_data_o[8]) );
  OA221X1 U24152 ( .IN1(n18490), .IN2(n2405), .IN3(n18487), .IN4(n2440), .IN5(
        n16448), .Q(n16441) );
  OA221X1 U24153 ( .IN1(n18502), .IN2(n2475), .IN3(n18499), .IN4(n2510), .IN5(
        n16447), .Q(n16442) );
  OA221X1 U24154 ( .IN1(n18514), .IN2(n2615), .IN3(n18511), .IN4(n2650), .IN5(
        n16446), .Q(n16443) );
  NAND4X0 U24155 ( .IN1(n16417), .IN2(n16418), .IN3(n16419), .IN4(n16420), 
        .QN(m1_data_o[9]) );
  OA221X1 U24156 ( .IN1(n18490), .IN2(n2404), .IN3(n18487), .IN4(n2439), .IN5(
        n16438), .Q(n16417) );
  OA221X1 U24157 ( .IN1(n18502), .IN2(n2474), .IN3(n18499), .IN4(n2509), .IN5(
        n16433), .Q(n16418) );
  OA221X1 U24158 ( .IN1(n18514), .IN2(n2614), .IN3(n18511), .IN4(n2649), .IN5(
        n16428), .Q(n16419) );
  NAND4X0 U24159 ( .IN1(n16673), .IN2(n16674), .IN3(n16675), .IN4(n16676), 
        .QN(m1_data_o[10]) );
  OA221X1 U24160 ( .IN1(n18490), .IN2(n2403), .IN3(n18485), .IN4(n2438), .IN5(
        n16680), .Q(n16673) );
  OA221X1 U24161 ( .IN1(n18502), .IN2(n2473), .IN3(n18497), .IN4(n2508), .IN5(
        n16679), .Q(n16674) );
  OA221X1 U24162 ( .IN1(n18514), .IN2(n2613), .IN3(n18509), .IN4(n2648), .IN5(
        n16678), .Q(n16675) );
  NAND4X0 U24163 ( .IN1(n16665), .IN2(n16666), .IN3(n16667), .IN4(n16668), 
        .QN(m1_data_o[11]) );
  OA221X1 U24164 ( .IN1(n18489), .IN2(n2402), .IN3(n18485), .IN4(n2437), .IN5(
        n16672), .Q(n16665) );
  OA221X1 U24165 ( .IN1(n18500), .IN2(n2472), .IN3(n18497), .IN4(n2507), .IN5(
        n16671), .Q(n16666) );
  OA221X1 U24166 ( .IN1(n18513), .IN2(n2612), .IN3(n18509), .IN4(n2647), .IN5(
        n16670), .Q(n16667) );
  NAND4X0 U24167 ( .IN1(n16657), .IN2(n16658), .IN3(n16659), .IN4(n16660), 
        .QN(m1_data_o[12]) );
  OA221X1 U24168 ( .IN1(n18488), .IN2(n2401), .IN3(n18485), .IN4(n2436), .IN5(
        n16664), .Q(n16657) );
  OA221X1 U24169 ( .IN1(n18501), .IN2(n2471), .IN3(n18497), .IN4(n2506), .IN5(
        n16663), .Q(n16658) );
  OA221X1 U24170 ( .IN1(n18512), .IN2(n2611), .IN3(n18509), .IN4(n2646), .IN5(
        n16662), .Q(n16659) );
  NAND4X0 U24171 ( .IN1(n16649), .IN2(n16650), .IN3(n16651), .IN4(n16652), 
        .QN(m1_data_o[13]) );
  OA221X1 U24172 ( .IN1(n18488), .IN2(n2400), .IN3(n18486), .IN4(n2435), .IN5(
        n16656), .Q(n16649) );
  OA221X1 U24173 ( .IN1(n18502), .IN2(n2470), .IN3(n18499), .IN4(n2505), .IN5(
        n16655), .Q(n16650) );
  OA221X1 U24174 ( .IN1(n18514), .IN2(n2610), .IN3(n18510), .IN4(n2645), .IN5(
        n16654), .Q(n16651) );
  NAND4X0 U24175 ( .IN1(n16641), .IN2(n16642), .IN3(n16643), .IN4(n16644), 
        .QN(m1_data_o[14]) );
  OA221X1 U24176 ( .IN1(n18490), .IN2(n2399), .IN3(n18486), .IN4(n2434), .IN5(
        n16648), .Q(n16641) );
  OA221X1 U24177 ( .IN1(n18500), .IN2(n2469), .IN3(n18497), .IN4(n2504), .IN5(
        n16647), .Q(n16642) );
  OA221X1 U24178 ( .IN1(n18512), .IN2(n2609), .IN3(n18510), .IN4(n2644), .IN5(
        n16646), .Q(n16643) );
  NAND4X0 U24179 ( .IN1(n16633), .IN2(n16634), .IN3(n16635), .IN4(n16636), 
        .QN(m1_data_o[15]) );
  OA221X1 U24180 ( .IN1(n18489), .IN2(n2398), .IN3(n18486), .IN4(n2433), .IN5(
        n16640), .Q(n16633) );
  OA221X1 U24181 ( .IN1(n18500), .IN2(n2468), .IN3(n18498), .IN4(n2503), .IN5(
        n16639), .Q(n16634) );
  OA221X1 U24182 ( .IN1(n18512), .IN2(n2608), .IN3(n18510), .IN4(n2643), .IN5(
        n16638), .Q(n16635) );
  NAND4X0 U24183 ( .IN1(n16625), .IN2(n16626), .IN3(n16627), .IN4(n16628), 
        .QN(m1_data_o[16]) );
  OA221X1 U24184 ( .IN1(n18488), .IN2(n2397), .IN3(n18486), .IN4(n2432), .IN5(
        n16632), .Q(n16625) );
  OA221X1 U24185 ( .IN1(n18501), .IN2(n2467), .IN3(n18498), .IN4(n2502), .IN5(
        n16631), .Q(n16626) );
  OA221X1 U24186 ( .IN1(n18513), .IN2(n2607), .IN3(n18510), .IN4(n2642), .IN5(
        n16630), .Q(n16627) );
  NAND4X0 U24187 ( .IN1(n16617), .IN2(n16618), .IN3(n16619), .IN4(n16620), 
        .QN(m1_data_o[17]) );
  OA221X1 U24188 ( .IN1(n18489), .IN2(n2396), .IN3(n18487), .IN4(n2431), .IN5(
        n16624), .Q(n16617) );
  OA221X1 U24189 ( .IN1(n18502), .IN2(n2466), .IN3(n18499), .IN4(n2501), .IN5(
        n16623), .Q(n16618) );
  OA221X1 U24190 ( .IN1(n18513), .IN2(n2606), .IN3(n18510), .IN4(n2641), .IN5(
        n16622), .Q(n16619) );
  NAND4X0 U24191 ( .IN1(n16609), .IN2(n16610), .IN3(n16611), .IN4(n16612), 
        .QN(m1_data_o[18]) );
  OA221X1 U24192 ( .IN1(n18489), .IN2(n2395), .IN3(n18485), .IN4(n2430), .IN5(
        n16616), .Q(n16609) );
  OA221X1 U24193 ( .IN1(n18501), .IN2(n2465), .IN3(n18497), .IN4(n2500), .IN5(
        n16615), .Q(n16610) );
  OA221X1 U24194 ( .IN1(n18513), .IN2(n2605), .IN3(n18511), .IN4(n2640), .IN5(
        n16614), .Q(n16611) );
  NAND4X0 U24195 ( .IN1(n16601), .IN2(n16602), .IN3(n16603), .IN4(n16604), 
        .QN(m1_data_o[19]) );
  OA221X1 U24196 ( .IN1(n18490), .IN2(n2394), .IN3(n18486), .IN4(n2429), .IN5(
        n16608), .Q(n16601) );
  OA221X1 U24197 ( .IN1(n18500), .IN2(n2464), .IN3(n18497), .IN4(n2499), .IN5(
        n16607), .Q(n16602) );
  OA221X1 U24198 ( .IN1(n18514), .IN2(n2604), .IN3(n18509), .IN4(n2639), .IN5(
        n16606), .Q(n16603) );
  NAND4X0 U24199 ( .IN1(n16585), .IN2(n16586), .IN3(n16587), .IN4(n16588), 
        .QN(m1_data_o[20]) );
  OA221X1 U24200 ( .IN1(n18488), .IN2(n2393), .IN3(n18485), .IN4(n2428), .IN5(
        n16592), .Q(n16585) );
  OA221X1 U24201 ( .IN1(n18500), .IN2(n2463), .IN3(n18498), .IN4(n2498), .IN5(
        n16591), .Q(n16586) );
  OA221X1 U24202 ( .IN1(n18512), .IN2(n2603), .IN3(n18509), .IN4(n2638), .IN5(
        n16590), .Q(n16587) );
  NAND4X0 U24203 ( .IN1(n16577), .IN2(n16578), .IN3(n16579), .IN4(n16580), 
        .QN(m1_data_o[21]) );
  OA221X1 U24204 ( .IN1(n18488), .IN2(n2392), .IN3(n18486), .IN4(n2427), .IN5(
        n16584), .Q(n16577) );
  OA221X1 U24205 ( .IN1(n18500), .IN2(n2462), .IN3(n18498), .IN4(n2497), .IN5(
        n16583), .Q(n16578) );
  OA221X1 U24206 ( .IN1(n18512), .IN2(n2602), .IN3(n18510), .IN4(n2637), .IN5(
        n16582), .Q(n16579) );
  NAND4X0 U24207 ( .IN1(n16569), .IN2(n16570), .IN3(n16571), .IN4(n16572), 
        .QN(m1_data_o[22]) );
  OA221X1 U24208 ( .IN1(n18488), .IN2(n2391), .IN3(n18487), .IN4(n2426), .IN5(
        n16576), .Q(n16569) );
  OA221X1 U24209 ( .IN1(n18500), .IN2(n2461), .IN3(n18498), .IN4(n2496), .IN5(
        n16575), .Q(n16570) );
  OA221X1 U24210 ( .IN1(n18512), .IN2(n2601), .IN3(n18511), .IN4(n2636), .IN5(
        n16574), .Q(n16571) );
  NAND4X0 U24211 ( .IN1(n16561), .IN2(n16562), .IN3(n16563), .IN4(n16564), 
        .QN(m1_data_o[23]) );
  OA221X1 U24212 ( .IN1(n18488), .IN2(n2390), .IN3(n18485), .IN4(n2425), .IN5(
        n16568), .Q(n16561) );
  OA221X1 U24213 ( .IN1(n18500), .IN2(n2460), .IN3(n18498), .IN4(n2495), .IN5(
        n16567), .Q(n16562) );
  OA221X1 U24214 ( .IN1(n18512), .IN2(n2600), .IN3(n18509), .IN4(n2635), .IN5(
        n16566), .Q(n16563) );
  NAND4X0 U24215 ( .IN1(n16553), .IN2(n16554), .IN3(n16555), .IN4(n16556), 
        .QN(m1_data_o[24]) );
  OA221X1 U24216 ( .IN1(n18489), .IN2(n2389), .IN3(n18487), .IN4(n2424), .IN5(
        n16560), .Q(n16553) );
  OA221X1 U24217 ( .IN1(n18501), .IN2(n2459), .IN3(n18499), .IN4(n2494), .IN5(
        n16559), .Q(n16554) );
  OA221X1 U24218 ( .IN1(n18512), .IN2(n2599), .IN3(n18509), .IN4(n2634), .IN5(
        n16558), .Q(n16555) );
  NAND4X0 U24219 ( .IN1(n16545), .IN2(n16546), .IN3(n16547), .IN4(n16548), 
        .QN(m1_data_o[25]) );
  OA221X1 U24220 ( .IN1(n18489), .IN2(n2388), .IN3(n18487), .IN4(n2423), .IN5(
        n16552), .Q(n16545) );
  OA221X1 U24221 ( .IN1(n18501), .IN2(n2458), .IN3(n18497), .IN4(n2493), .IN5(
        n16551), .Q(n16546) );
  OA221X1 U24222 ( .IN1(n18514), .IN2(n2598), .IN3(n18510), .IN4(n2633), .IN5(
        n16550), .Q(n16547) );
  NAND4X0 U24223 ( .IN1(n16537), .IN2(n16538), .IN3(n16539), .IN4(n16540), 
        .QN(m1_data_o[26]) );
  OA221X1 U24224 ( .IN1(n18489), .IN2(n2387), .IN3(n18485), .IN4(n2422), .IN5(
        n16544), .Q(n16537) );
  OA221X1 U24225 ( .IN1(n18501), .IN2(n2457), .IN3(n18498), .IN4(n2492), .IN5(
        n16543), .Q(n16538) );
  OA221X1 U24226 ( .IN1(n18513), .IN2(n2597), .IN3(n18511), .IN4(n2632), .IN5(
        n16542), .Q(n16539) );
  NAND4X0 U24227 ( .IN1(n16529), .IN2(n16530), .IN3(n16531), .IN4(n16532), 
        .QN(m1_data_o[27]) );
  OA221X1 U24228 ( .IN1(n18489), .IN2(n2386), .IN3(n18486), .IN4(n2421), .IN5(
        n16536), .Q(n16529) );
  OA221X1 U24229 ( .IN1(n18501), .IN2(n2456), .IN3(n18499), .IN4(n2491), .IN5(
        n16535), .Q(n16530) );
  OA221X1 U24230 ( .IN1(n18512), .IN2(n2596), .IN3(n18509), .IN4(n2631), .IN5(
        n16534), .Q(n16531) );
  NAND4X0 U24231 ( .IN1(n16521), .IN2(n16522), .IN3(n16523), .IN4(n16524), 
        .QN(m1_data_o[28]) );
  OA221X1 U24232 ( .IN1(n18490), .IN2(n2385), .IN3(n18486), .IN4(n2420), .IN5(
        n16528), .Q(n16521) );
  OA221X1 U24233 ( .IN1(n18501), .IN2(n2455), .IN3(n18499), .IN4(n2490), .IN5(
        n16527), .Q(n16522) );
  OA221X1 U24234 ( .IN1(n18513), .IN2(n2595), .IN3(n18509), .IN4(n2630), .IN5(
        n16526), .Q(n16523) );
  NAND4X0 U24235 ( .IN1(n16513), .IN2(n16514), .IN3(n16515), .IN4(n16516), 
        .QN(m1_data_o[29]) );
  OA221X1 U24236 ( .IN1(n18489), .IN2(n2384), .IN3(n18487), .IN4(n2419), .IN5(
        n16520), .Q(n16513) );
  OA221X1 U24237 ( .IN1(n18501), .IN2(n2454), .IN3(n18498), .IN4(n2489), .IN5(
        n16519), .Q(n16514) );
  OA221X1 U24238 ( .IN1(n18513), .IN2(n2594), .IN3(n18510), .IN4(n2629), .IN5(
        n16518), .Q(n16515) );
  NAND4X0 U24239 ( .IN1(n16497), .IN2(n16498), .IN3(n16499), .IN4(n16500), 
        .QN(m1_data_o[30]) );
  OA221X1 U24240 ( .IN1(n18488), .IN2(n2383), .IN3(n18485), .IN4(n2418), .IN5(
        n16504), .Q(n16497) );
  OA221X1 U24241 ( .IN1(n18502), .IN2(n2453), .IN3(n18497), .IN4(n2488), .IN5(
        n16503), .Q(n16498) );
  OA221X1 U24242 ( .IN1(n18513), .IN2(n2593), .IN3(n18511), .IN4(n2628), .IN5(
        n16502), .Q(n16499) );
  NAND4X0 U24243 ( .IN1(n16489), .IN2(n16490), .IN3(n16491), .IN4(n16492), 
        .QN(m1_data_o[31]) );
  OA221X1 U24244 ( .IN1(n18490), .IN2(n2382), .IN3(n18487), .IN4(n2417), .IN5(
        n16496), .Q(n16489) );
  OA221X1 U24245 ( .IN1(n18500), .IN2(n2452), .IN3(n18499), .IN4(n2487), .IN5(
        n16495), .Q(n16490) );
  OA221X1 U24246 ( .IN1(n18514), .IN2(n2592), .IN3(n18510), .IN4(n2627), .IN5(
        n16494), .Q(n16491) );
  NAND4X0 U24247 ( .IN1(n16705), .IN2(n16706), .IN3(n16707), .IN4(n16708), 
        .QN(m0_rty_o) );
  OA221X1 U24248 ( .IN1(n8854), .IN2(n2346), .IN3(n8558), .IN4(n2696), .IN5(
        n16713), .Q(n16705) );
  OA221X1 U24249 ( .IN1(n6598), .IN2(n2416), .IN3(n6302), .IN4(n2451), .IN5(
        n16710), .Q(n16707) );
  OA221X1 U24250 ( .IN1(n4822), .IN2(n2626), .IN3(n4526), .IN4(n2661), .IN5(
        n16709), .Q(n16708) );
  NAND4X0 U24251 ( .IN1(n16714), .IN2(n16715), .IN3(n16716), .IN4(n16717), 
        .QN(m0_err_o) );
  OA221X1 U24252 ( .IN1(n8854), .IN2(n2345), .IN3(n8558), .IN4(n2695), .IN5(
        n16721), .Q(n16714) );
  OA221X1 U24253 ( .IN1(n6598), .IN2(n2415), .IN3(n6302), .IN4(n2450), .IN5(
        n16719), .Q(n16716) );
  OA221X1 U24254 ( .IN1(n4822), .IN2(n2625), .IN3(n4526), .IN4(n2660), .IN5(
        n16718), .Q(n16717) );
  NAND4X0 U24255 ( .IN1(n16994), .IN2(n16995), .IN3(n16996), .IN4(n16997), 
        .QN(m0_ack_o) );
  OA221X1 U24256 ( .IN1(n8854), .IN2(n2344), .IN3(n8558), .IN4(n2694), .IN5(
        n17127), .Q(n16994) );
  OA221X1 U24257 ( .IN1(n6598), .IN2(n2414), .IN3(n6302), .IN4(n2449), .IN5(
        n17033), .Q(n16996) );
  OA221X1 U24258 ( .IN1(n4822), .IN2(n2624), .IN3(n4526), .IN4(n2659), .IN5(
        n16998), .Q(n16997) );
  NAND4X0 U24259 ( .IN1(n16986), .IN2(n16987), .IN3(n16988), .IN4(n16989), 
        .QN(m0_data_o[0]) );
  OA221X1 U24260 ( .IN1(n18440), .IN2(n2413), .IN3(n16742), .IN4(n2448), .IN5(
        n16993), .Q(n16986) );
  OA221X1 U24261 ( .IN1(n18452), .IN2(n2483), .IN3(n18449), .IN4(n2518), .IN5(
        n16992), .Q(n16987) );
  OA221X1 U24262 ( .IN1(n18465), .IN2(n2623), .IN3(n18461), .IN4(n2658), .IN5(
        n16991), .Q(n16988) );
  NAND4X0 U24263 ( .IN1(n16898), .IN2(n16899), .IN3(n16900), .IN4(n16901), 
        .QN(m0_data_o[1]) );
  OA221X1 U24264 ( .IN1(n18442), .IN2(n2412), .IN3(n18438), .IN4(n2447), .IN5(
        n16905), .Q(n16898) );
  OA221X1 U24265 ( .IN1(n18454), .IN2(n2482), .IN3(n18449), .IN4(n2517), .IN5(
        n16904), .Q(n16899) );
  OA221X1 U24266 ( .IN1(n18466), .IN2(n2622), .IN3(n18461), .IN4(n2657), .IN5(
        n16903), .Q(n16900) );
  NAND4X0 U24267 ( .IN1(n16810), .IN2(n16811), .IN3(n16812), .IN4(n16813), 
        .QN(m0_data_o[2]) );
  OA221X1 U24268 ( .IN1(n18440), .IN2(n2411), .IN3(n18438), .IN4(n2446), .IN5(
        n16817), .Q(n16810) );
  OA221X1 U24269 ( .IN1(n18454), .IN2(n2481), .IN3(n18451), .IN4(n2516), .IN5(
        n16816), .Q(n16811) );
  OA221X1 U24270 ( .IN1(n18466), .IN2(n2621), .IN3(n18462), .IN4(n2656), .IN5(
        n16815), .Q(n16812) );
  NAND4X0 U24271 ( .IN1(n16786), .IN2(n16787), .IN3(n16788), .IN4(n16789), 
        .QN(m0_data_o[3]) );
  OA221X1 U24272 ( .IN1(n18442), .IN2(n2410), .IN3(n18438), .IN4(n2445), .IN5(
        n16793), .Q(n16786) );
  OA221X1 U24273 ( .IN1(n18454), .IN2(n2480), .IN3(n18450), .IN4(n2515), .IN5(
        n16792), .Q(n16787) );
  OA221X1 U24274 ( .IN1(n18466), .IN2(n2620), .IN3(n18462), .IN4(n2655), .IN5(
        n16791), .Q(n16788) );
  NAND4X0 U24275 ( .IN1(n16778), .IN2(n16779), .IN3(n16780), .IN4(n16781), 
        .QN(m0_data_o[4]) );
  OA221X1 U24276 ( .IN1(n18440), .IN2(n2409), .IN3(n18437), .IN4(n2444), .IN5(
        n16785), .Q(n16778) );
  OA221X1 U24277 ( .IN1(n18452), .IN2(n2479), .IN3(n18451), .IN4(n2514), .IN5(
        n16784), .Q(n16779) );
  OA221X1 U24278 ( .IN1(n18465), .IN2(n2619), .IN3(n18463), .IN4(n2654), .IN5(
        n16783), .Q(n16780) );
  NAND4X0 U24279 ( .IN1(n16770), .IN2(n16771), .IN3(n16772), .IN4(n16773), 
        .QN(m0_data_o[5]) );
  OA221X1 U24280 ( .IN1(n18441), .IN2(n2408), .IN3(n16742), .IN4(n2443), .IN5(
        n16777), .Q(n16770) );
  OA221X1 U24281 ( .IN1(n18453), .IN2(n2478), .IN3(n18451), .IN4(n2513), .IN5(
        n16776), .Q(n16771) );
  OA221X1 U24282 ( .IN1(n18464), .IN2(n2618), .IN3(n18462), .IN4(n2653), .IN5(
        n16775), .Q(n16772) );
  NAND4X0 U24283 ( .IN1(n16762), .IN2(n16763), .IN3(n16764), .IN4(n16765), 
        .QN(m0_data_o[6]) );
  OA221X1 U24284 ( .IN1(n18442), .IN2(n2407), .IN3(n18438), .IN4(n2442), .IN5(
        n16769), .Q(n16762) );
  OA221X1 U24285 ( .IN1(n18454), .IN2(n2477), .IN3(n18451), .IN4(n2512), .IN5(
        n16768), .Q(n16763) );
  OA221X1 U24286 ( .IN1(n18466), .IN2(n2617), .IN3(n18463), .IN4(n2652), .IN5(
        n16767), .Q(n16764) );
  NAND4X0 U24287 ( .IN1(n16754), .IN2(n16755), .IN3(n16756), .IN4(n16757), 
        .QN(m0_data_o[7]) );
  OA221X1 U24288 ( .IN1(n18442), .IN2(n2406), .IN3(n18438), .IN4(n2441), .IN5(
        n16761), .Q(n16754) );
  OA221X1 U24289 ( .IN1(n18454), .IN2(n2476), .IN3(n18451), .IN4(n2511), .IN5(
        n16760), .Q(n16755) );
  OA221X1 U24290 ( .IN1(n18466), .IN2(n2616), .IN3(n18463), .IN4(n2651), .IN5(
        n16759), .Q(n16756) );
  NAND4X0 U24291 ( .IN1(n16746), .IN2(n16747), .IN3(n16748), .IN4(n16749), 
        .QN(m0_data_o[8]) );
  OA221X1 U24292 ( .IN1(n18442), .IN2(n2405), .IN3(n18438), .IN4(n2440), .IN5(
        n16753), .Q(n16746) );
  OA221X1 U24293 ( .IN1(n18454), .IN2(n2475), .IN3(n18451), .IN4(n2510), .IN5(
        n16752), .Q(n16747) );
  OA221X1 U24294 ( .IN1(n18466), .IN2(n2615), .IN3(n18463), .IN4(n2650), .IN5(
        n16751), .Q(n16748) );
  NAND4X0 U24295 ( .IN1(n16722), .IN2(n16723), .IN3(n16724), .IN4(n16725), 
        .QN(m0_data_o[9]) );
  OA221X1 U24296 ( .IN1(n18442), .IN2(n2404), .IN3(n18438), .IN4(n2439), .IN5(
        n16743), .Q(n16722) );
  OA221X1 U24297 ( .IN1(n18454), .IN2(n2474), .IN3(n18451), .IN4(n2509), .IN5(
        n16738), .Q(n16723) );
  OA221X1 U24298 ( .IN1(n18466), .IN2(n2614), .IN3(n18463), .IN4(n2649), .IN5(
        n16733), .Q(n16724) );
  NAND4X0 U24299 ( .IN1(n16978), .IN2(n16979), .IN3(n16980), .IN4(n16981), 
        .QN(m0_data_o[10]) );
  OA221X1 U24300 ( .IN1(n18441), .IN2(n2403), .IN3(n16742), .IN4(n2438), .IN5(
        n16985), .Q(n16978) );
  OA221X1 U24301 ( .IN1(n18454), .IN2(n2473), .IN3(n18449), .IN4(n2508), .IN5(
        n16984), .Q(n16979) );
  OA221X1 U24302 ( .IN1(n18464), .IN2(n2613), .IN3(n18461), .IN4(n2648), .IN5(
        n16983), .Q(n16980) );
  NAND4X0 U24303 ( .IN1(n16970), .IN2(n16971), .IN3(n16972), .IN4(n16973), 
        .QN(m0_data_o[11]) );
  OA221X1 U24304 ( .IN1(n18440), .IN2(n2402), .IN3(n16742), .IN4(n2437), .IN5(
        n16977), .Q(n16970) );
  OA221X1 U24305 ( .IN1(n18452), .IN2(n2472), .IN3(n18449), .IN4(n2507), .IN5(
        n16976), .Q(n16971) );
  OA221X1 U24306 ( .IN1(n18466), .IN2(n2612), .IN3(n18461), .IN4(n2647), .IN5(
        n16975), .Q(n16972) );
  NAND4X0 U24307 ( .IN1(n16962), .IN2(n16963), .IN3(n16964), .IN4(n16965), 
        .QN(m0_data_o[12]) );
  OA221X1 U24308 ( .IN1(n18441), .IN2(n2401), .IN3(n16742), .IN4(n2436), .IN5(
        n16969), .Q(n16962) );
  OA221X1 U24309 ( .IN1(n18453), .IN2(n2471), .IN3(n18449), .IN4(n2506), .IN5(
        n16968), .Q(n16963) );
  OA221X1 U24310 ( .IN1(n18465), .IN2(n2611), .IN3(n18461), .IN4(n2646), .IN5(
        n16967), .Q(n16964) );
  NAND4X0 U24311 ( .IN1(n16954), .IN2(n16955), .IN3(n16956), .IN4(n16957), 
        .QN(m0_data_o[13]) );
  OA221X1 U24312 ( .IN1(n18440), .IN2(n2400), .IN3(n18437), .IN4(n2435), .IN5(
        n16961), .Q(n16954) );
  OA221X1 U24313 ( .IN1(n18452), .IN2(n2470), .IN3(n18450), .IN4(n2505), .IN5(
        n16960), .Q(n16955) );
  OA221X1 U24314 ( .IN1(n18464), .IN2(n2610), .IN3(n18463), .IN4(n2645), .IN5(
        n16959), .Q(n16956) );
  NAND4X0 U24315 ( .IN1(n16946), .IN2(n16947), .IN3(n16948), .IN4(n16949), 
        .QN(m0_data_o[14]) );
  OA221X1 U24316 ( .IN1(n18440), .IN2(n2399), .IN3(n18437), .IN4(n2434), .IN5(
        n16953), .Q(n16946) );
  OA221X1 U24317 ( .IN1(n18452), .IN2(n2469), .IN3(n18450), .IN4(n2504), .IN5(
        n16952), .Q(n16947) );
  OA221X1 U24318 ( .IN1(n18464), .IN2(n2609), .IN3(n18461), .IN4(n2644), .IN5(
        n16951), .Q(n16948) );
  NAND4X0 U24319 ( .IN1(n16938), .IN2(n16939), .IN3(n16940), .IN4(n16941), 
        .QN(m0_data_o[15]) );
  OA221X1 U24320 ( .IN1(n18440), .IN2(n2398), .IN3(n18437), .IN4(n2433), .IN5(
        n16945), .Q(n16938) );
  OA221X1 U24321 ( .IN1(n18452), .IN2(n2468), .IN3(n18450), .IN4(n2503), .IN5(
        n16944), .Q(n16939) );
  OA221X1 U24322 ( .IN1(n18464), .IN2(n2608), .IN3(n18462), .IN4(n2643), .IN5(
        n16943), .Q(n16940) );
  NAND4X0 U24323 ( .IN1(n16930), .IN2(n16931), .IN3(n16932), .IN4(n16933), 
        .QN(m0_data_o[16]) );
  OA221X1 U24324 ( .IN1(n18440), .IN2(n2397), .IN3(n18437), .IN4(n2432), .IN5(
        n16937), .Q(n16930) );
  OA221X1 U24325 ( .IN1(n18452), .IN2(n2467), .IN3(n18450), .IN4(n2502), .IN5(
        n16936), .Q(n16931) );
  OA221X1 U24326 ( .IN1(n18464), .IN2(n2607), .IN3(n18462), .IN4(n2642), .IN5(
        n16935), .Q(n16932) );
  NAND4X0 U24327 ( .IN1(n16922), .IN2(n16923), .IN3(n16924), .IN4(n16925), 
        .QN(m0_data_o[17]) );
  OA221X1 U24328 ( .IN1(n18441), .IN2(n2396), .IN3(n18437), .IN4(n2431), .IN5(
        n16929), .Q(n16922) );
  OA221X1 U24329 ( .IN1(n18453), .IN2(n2466), .IN3(n18450), .IN4(n2501), .IN5(
        n16928), .Q(n16923) );
  OA221X1 U24330 ( .IN1(n18464), .IN2(n2606), .IN3(n18463), .IN4(n2641), .IN5(
        n16927), .Q(n16924) );
  NAND4X0 U24331 ( .IN1(n16914), .IN2(n16915), .IN3(n16916), .IN4(n16917), 
        .QN(m0_data_o[18]) );
  OA221X1 U24332 ( .IN1(n18441), .IN2(n2395), .IN3(n18438), .IN4(n2430), .IN5(
        n16921), .Q(n16914) );
  OA221X1 U24333 ( .IN1(n18453), .IN2(n2465), .IN3(n18451), .IN4(n2500), .IN5(
        n16920), .Q(n16915) );
  OA221X1 U24334 ( .IN1(n18465), .IN2(n2605), .IN3(n18461), .IN4(n2640), .IN5(
        n16919), .Q(n16916) );
  NAND4X0 U24335 ( .IN1(n16906), .IN2(n16907), .IN3(n16908), .IN4(n16909), 
        .QN(m0_data_o[19]) );
  OA221X1 U24336 ( .IN1(n18440), .IN2(n2394), .IN3(n18438), .IN4(n2429), .IN5(
        n16913), .Q(n16906) );
  OA221X1 U24337 ( .IN1(n18452), .IN2(n2464), .IN3(n18449), .IN4(n2499), .IN5(
        n16912), .Q(n16907) );
  OA221X1 U24338 ( .IN1(n18466), .IN2(n2604), .IN3(n18461), .IN4(n2639), .IN5(
        n16911), .Q(n16908) );
  NAND4X0 U24339 ( .IN1(n16890), .IN2(n16891), .IN3(n16892), .IN4(n16893), 
        .QN(m0_data_o[20]) );
  OA221X1 U24340 ( .IN1(n18441), .IN2(n2393), .IN3(n16742), .IN4(n2428), .IN5(
        n16897), .Q(n16890) );
  OA221X1 U24341 ( .IN1(n18453), .IN2(n2463), .IN3(n18449), .IN4(n2498), .IN5(
        n16896), .Q(n16891) );
  OA221X1 U24342 ( .IN1(n18464), .IN2(n2603), .IN3(n18462), .IN4(n2638), .IN5(
        n16895), .Q(n16892) );
  NAND4X0 U24343 ( .IN1(n16882), .IN2(n16883), .IN3(n16884), .IN4(n16885), 
        .QN(m0_data_o[21]) );
  OA221X1 U24344 ( .IN1(n18441), .IN2(n2392), .IN3(n16742), .IN4(n2427), .IN5(
        n16889), .Q(n16882) );
  OA221X1 U24345 ( .IN1(n18453), .IN2(n2462), .IN3(n18450), .IN4(n2497), .IN5(
        n16888), .Q(n16883) );
  OA221X1 U24346 ( .IN1(n18464), .IN2(n2602), .IN3(n18462), .IN4(n2637), .IN5(
        n16887), .Q(n16884) );
  NAND4X0 U24347 ( .IN1(n16874), .IN2(n16875), .IN3(n16876), .IN4(n16877), 
        .QN(m0_data_o[22]) );
  OA221X1 U24348 ( .IN1(n18441), .IN2(n2391), .IN3(n16742), .IN4(n2426), .IN5(
        n16881), .Q(n16874) );
  OA221X1 U24349 ( .IN1(n18453), .IN2(n2461), .IN3(n18451), .IN4(n2496), .IN5(
        n16880), .Q(n16875) );
  OA221X1 U24350 ( .IN1(n18465), .IN2(n2601), .IN3(n18462), .IN4(n2636), .IN5(
        n16879), .Q(n16876) );
  NAND4X0 U24351 ( .IN1(n16866), .IN2(n16867), .IN3(n16868), .IN4(n16869), 
        .QN(m0_data_o[23]) );
  OA221X1 U24352 ( .IN1(n18441), .IN2(n2390), .IN3(n16742), .IN4(n2425), .IN5(
        n16873), .Q(n16866) );
  OA221X1 U24353 ( .IN1(n18453), .IN2(n2460), .IN3(n18449), .IN4(n2495), .IN5(
        n16872), .Q(n16867) );
  OA221X1 U24354 ( .IN1(n18466), .IN2(n2600), .IN3(n18462), .IN4(n2635), .IN5(
        n16871), .Q(n16868) );
  NAND4X0 U24355 ( .IN1(n16858), .IN2(n16859), .IN3(n16860), .IN4(n16861), 
        .QN(m0_data_o[24]) );
  OA221X1 U24356 ( .IN1(n18441), .IN2(n2389), .IN3(n18437), .IN4(n2424), .IN5(
        n16865), .Q(n16858) );
  OA221X1 U24357 ( .IN1(n18453), .IN2(n2459), .IN3(n18449), .IN4(n2494), .IN5(
        n16864), .Q(n16859) );
  OA221X1 U24358 ( .IN1(n18465), .IN2(n2599), .IN3(n18463), .IN4(n2634), .IN5(
        n16863), .Q(n16860) );
  NAND4X0 U24359 ( .IN1(n16850), .IN2(n16851), .IN3(n16852), .IN4(n16853), 
        .QN(m0_data_o[25]) );
  OA221X1 U24360 ( .IN1(n18442), .IN2(n2388), .IN3(n18437), .IN4(n2423), .IN5(
        n16857), .Q(n16850) );
  OA221X1 U24361 ( .IN1(n18454), .IN2(n2458), .IN3(n18450), .IN4(n2493), .IN5(
        n16856), .Q(n16851) );
  OA221X1 U24362 ( .IN1(n18465), .IN2(n2598), .IN3(n18461), .IN4(n2633), .IN5(
        n16855), .Q(n16852) );
  NAND4X0 U24363 ( .IN1(n16842), .IN2(n16843), .IN3(n16844), .IN4(n16845), 
        .QN(m0_data_o[26]) );
  OA221X1 U24364 ( .IN1(n18441), .IN2(n2387), .IN3(n16742), .IN4(n2422), .IN5(
        n16849), .Q(n16842) );
  OA221X1 U24365 ( .IN1(n18453), .IN2(n2457), .IN3(n18451), .IN4(n2492), .IN5(
        n16848), .Q(n16843) );
  OA221X1 U24366 ( .IN1(n18465), .IN2(n2597), .IN3(n18462), .IN4(n2632), .IN5(
        n16847), .Q(n16844) );
  NAND4X0 U24367 ( .IN1(n16834), .IN2(n16835), .IN3(n16836), .IN4(n16837), 
        .QN(m0_data_o[27]) );
  OA221X1 U24368 ( .IN1(n18440), .IN2(n2386), .IN3(n16742), .IN4(n2421), .IN5(
        n16841), .Q(n16834) );
  OA221X1 U24369 ( .IN1(n18452), .IN2(n2456), .IN3(n18449), .IN4(n2491), .IN5(
        n16840), .Q(n16835) );
  OA221X1 U24370 ( .IN1(n18465), .IN2(n2596), .IN3(n18463), .IN4(n2631), .IN5(
        n16839), .Q(n16836) );
  NAND4X0 U24371 ( .IN1(n16826), .IN2(n16827), .IN3(n16828), .IN4(n16829), 
        .QN(m0_data_o[28]) );
  OA221X1 U24372 ( .IN1(n18442), .IN2(n2385), .IN3(n16742), .IN4(n2420), .IN5(
        n16833), .Q(n16826) );
  OA221X1 U24373 ( .IN1(n18452), .IN2(n2455), .IN3(n18449), .IN4(n2490), .IN5(
        n16832), .Q(n16827) );
  OA221X1 U24374 ( .IN1(n18466), .IN2(n2595), .IN3(n18463), .IN4(n2630), .IN5(
        n16831), .Q(n16828) );
  NAND4X0 U24375 ( .IN1(n16818), .IN2(n16819), .IN3(n16820), .IN4(n16821), 
        .QN(m0_data_o[29]) );
  OA221X1 U24376 ( .IN1(n18440), .IN2(n2384), .IN3(n18437), .IN4(n2419), .IN5(
        n16825), .Q(n16818) );
  OA221X1 U24377 ( .IN1(n18453), .IN2(n2454), .IN3(n18450), .IN4(n2489), .IN5(
        n16824), .Q(n16819) );
  OA221X1 U24378 ( .IN1(n18464), .IN2(n2594), .IN3(n18461), .IN4(n2629), .IN5(
        n16823), .Q(n16820) );
  NAND4X0 U24379 ( .IN1(n16802), .IN2(n16803), .IN3(n16804), .IN4(n16805), 
        .QN(m0_data_o[30]) );
  OA221X1 U24380 ( .IN1(n18442), .IN2(n2383), .IN3(n18438), .IN4(n2418), .IN5(
        n16809), .Q(n16802) );
  OA221X1 U24381 ( .IN1(n18454), .IN2(n2453), .IN3(n18451), .IN4(n2488), .IN5(
        n16808), .Q(n16803) );
  OA221X1 U24382 ( .IN1(n18465), .IN2(n2593), .IN3(n18462), .IN4(n2628), .IN5(
        n16807), .Q(n16804) );
  NAND4X0 U24383 ( .IN1(n16794), .IN2(n16795), .IN3(n16796), .IN4(n16797), 
        .QN(m0_data_o[31]) );
  OA221X1 U24384 ( .IN1(n18442), .IN2(n2382), .IN3(n18437), .IN4(n2417), .IN5(
        n16801), .Q(n16794) );
  OA221X1 U24385 ( .IN1(n18454), .IN2(n2452), .IN3(n18450), .IN4(n2487), .IN5(
        n16800), .Q(n16795) );
  OA221X1 U24386 ( .IN1(n18465), .IN2(n2592), .IN3(n18463), .IN4(n2627), .IN5(
        n16799), .Q(n16796) );
  NAND4X0 U24387 ( .IN1(n18164), .IN2(n13670), .IN3(n13671), .IN4(n13672), 
        .QN(n13629) );
  NOR2X0 U24388 ( .IN1(n13677), .IN2(n13678), .QN(n13671) );
  NOR4X0 U24389 ( .IN1(n13673), .IN2(n13674), .IN3(n13675), .IN4(n13676), .QN(
        n13672) );
  NAND4X0 U24390 ( .IN1(n18165), .IN2(n13361), .IN3(n13362), .IN4(n13363), 
        .QN(n13320) );
  NOR2X0 U24391 ( .IN1(n13368), .IN2(n13369), .QN(n13362) );
  NOR4X0 U24392 ( .IN1(n13364), .IN2(n13365), .IN3(n13366), .IN4(n13367), .QN(
        n13363) );
  NAND4X0 U24393 ( .IN1(n18166), .IN2(n11195), .IN3(n11196), .IN4(n11197), 
        .QN(n11154) );
  NOR2X0 U24394 ( .IN1(n11202), .IN2(n11203), .QN(n11196) );
  NOR4X0 U24395 ( .IN1(n11198), .IN2(n11199), .IN3(n11200), .IN4(n11201), .QN(
        n11197) );
  NAND4X0 U24396 ( .IN1(n18168), .IN2(n13052), .IN3(n13053), .IN4(n13054), 
        .QN(n13011) );
  NOR2X0 U24397 ( .IN1(n13059), .IN2(n13060), .QN(n13053) );
  NOR4X0 U24398 ( .IN1(n13055), .IN2(n13056), .IN3(n13057), .IN4(n13058), .QN(
        n13054) );
  NAND4X0 U24399 ( .IN1(n18170), .IN2(n12743), .IN3(n12744), .IN4(n12745), 
        .QN(n12702) );
  NOR2X0 U24400 ( .IN1(n12750), .IN2(n12751), .QN(n12744) );
  NOR4X0 U24401 ( .IN1(n12746), .IN2(n12747), .IN3(n12748), .IN4(n12749), .QN(
        n12745) );
  NAND4X0 U24402 ( .IN1(n18172), .IN2(n10886), .IN3(n10887), .IN4(n10888), 
        .QN(n10845) );
  NOR2X0 U24403 ( .IN1(n10893), .IN2(n10894), .QN(n10887) );
  NOR4X0 U24404 ( .IN1(n10889), .IN2(n10890), .IN3(n10891), .IN4(n10892), .QN(
        n10888) );
  NAND4X0 U24405 ( .IN1(n18174), .IN2(n10576), .IN3(n10577), .IN4(n10578), 
        .QN(n10535) );
  NOR2X0 U24406 ( .IN1(n10583), .IN2(n10584), .QN(n10577) );
  NOR4X0 U24407 ( .IN1(n10579), .IN2(n10580), .IN3(n10581), .IN4(n10582), .QN(
        n10578) );
  NAND4X0 U24408 ( .IN1(n18176), .IN2(n12434), .IN3(n12435), .IN4(n12436), 
        .QN(n12393) );
  NOR2X0 U24409 ( .IN1(n12441), .IN2(n12442), .QN(n12435) );
  NOR4X0 U24410 ( .IN1(n12437), .IN2(n12438), .IN3(n12439), .IN4(n12440), .QN(
        n12436) );
  NAND4X0 U24411 ( .IN1(n18177), .IN2(n12125), .IN3(n12126), .IN4(n12127), 
        .QN(n12084) );
  NOR2X0 U24412 ( .IN1(n12132), .IN2(n12133), .QN(n12126) );
  NOR4X0 U24413 ( .IN1(n12128), .IN2(n12129), .IN3(n12130), .IN4(n12131), .QN(
        n12127) );
  NAND4X0 U24414 ( .IN1(n18179), .IN2(n10267), .IN3(n10268), .IN4(n10269), 
        .QN(n10226) );
  NOR2X0 U24415 ( .IN1(n10274), .IN2(n10275), .QN(n10268) );
  NOR4X0 U24416 ( .IN1(n10270), .IN2(n10271), .IN3(n10272), .IN4(n10273), .QN(
        n10269) );
  NAND4X0 U24417 ( .IN1(n18181), .IN2(n9957), .IN3(n9958), .IN4(n9959), .QN(
        n9916) );
  NOR2X0 U24418 ( .IN1(n9964), .IN2(n9965), .QN(n9958) );
  NOR4X0 U24419 ( .IN1(n9960), .IN2(n9961), .IN3(n9962), .IN4(n9963), .QN(
        n9959) );
  NAND4X0 U24420 ( .IN1(n18183), .IN2(n11815), .IN3(n11816), .IN4(n11817), 
        .QN(n11774) );
  NOR2X0 U24421 ( .IN1(n11822), .IN2(n11823), .QN(n11816) );
  NOR4X0 U24422 ( .IN1(n11818), .IN2(n11819), .IN3(n11820), .IN4(n11821), .QN(
        n11817) );
  NAND4X0 U24423 ( .IN1(n18185), .IN2(n11505), .IN3(n11506), .IN4(n11507), 
        .QN(n11464) );
  NOR2X0 U24424 ( .IN1(n11512), .IN2(n11513), .QN(n11506) );
  NOR4X0 U24425 ( .IN1(n11508), .IN2(n11509), .IN3(n11510), .IN4(n11511), .QN(
        n11507) );
  NAND4X0 U24426 ( .IN1(n18186), .IN2(n9647), .IN3(n9648), .IN4(n9649), .QN(
        n9606) );
  NOR2X0 U24427 ( .IN1(n9654), .IN2(n9655), .QN(n9648) );
  NOR4X0 U24428 ( .IN1(n9650), .IN2(n9651), .IN3(n9652), .IN4(n9653), .QN(
        n9649) );
  NAND4X0 U24429 ( .IN1(n18188), .IN2(n9336), .IN3(n9337), .IN4(n9338), .QN(
        n9295) );
  NOR2X0 U24430 ( .IN1(n9343), .IN2(n9344), .QN(n9337) );
  NOR4X0 U24431 ( .IN1(n9339), .IN2(n9340), .IN3(n9341), .IN4(n9342), .QN(
        n9338) );
  AO221X1 U24432 ( .IN1(n13989), .IN2(n13990), .IN3(n13987), .IN4(n4226), 
        .IN5(n13991), .Q(n13954) );
  NOR2X0 U24433 ( .IN1(n13968), .IN2(n13965), .QN(n13989) );
  AO22X1 U24434 ( .IN1(n4224), .IN2(n13990), .IN3(n4223), .IN4(n13992), .Q(
        n13991) );
  INVX0 U24435 ( .IN(n13967), .QN(n4224) );
  AO221X1 U24436 ( .IN1(n14129), .IN2(n14130), .IN3(n14127), .IN4(n4234), 
        .IN5(n14131), .Q(n14094) );
  NOR2X0 U24437 ( .IN1(n14108), .IN2(n14105), .QN(n14129) );
  AO22X1 U24438 ( .IN1(n4232), .IN2(n14130), .IN3(n4231), .IN4(n14132), .Q(
        n14131) );
  INVX0 U24439 ( .IN(n14107), .QN(n4232) );
  ISOLANDX1 U24440 ( .D(n13909), .ISO(n3390), .Q(n13880) );
  ISOLANDX1 U24441 ( .D(n13600), .ISO(n3391), .Q(n13571) );
  ISOLANDX1 U24442 ( .D(n11434), .ISO(n3383), .Q(n11405) );
  ISOLANDX1 U24443 ( .D(n13291), .ISO(n3392), .Q(n13262) );
  ISOLANDX1 U24444 ( .D(n12982), .ISO(n3393), .Q(n12953) );
  ISOLANDX1 U24445 ( .D(n11125), .ISO(n3384), .Q(n11096) );
  ISOLANDX1 U24446 ( .D(n10815), .ISO(n3385), .Q(n10786) );
  ISOLANDX1 U24447 ( .D(n12673), .ISO(n3394), .Q(n12644) );
  ISOLANDX1 U24448 ( .D(n12364), .ISO(n3395), .Q(n12335) );
  ISOLANDX1 U24449 ( .D(n10506), .ISO(n3386), .Q(n10477) );
  ISOLANDX1 U24450 ( .D(n10196), .ISO(n3387), .Q(n10167) );
  ISOLANDX1 U24451 ( .D(n12054), .ISO(n3396), .Q(n12025) );
  ISOLANDX1 U24452 ( .D(n11744), .ISO(n3397), .Q(n11715) );
  ISOLANDX1 U24453 ( .D(n9886), .ISO(n3388), .Q(n9857) );
  ISOLANDX1 U24454 ( .D(n9575), .ISO(n3389), .Q(n9546) );
  ISOLANDX1 U24455 ( .D(n14183), .ISO(n3381), .Q(n14154) );
  AO21X1 U24456 ( .IN1(n3881), .IN2(n13909), .IN3(n3878), .Q(n13918) );
  AO21X1 U24457 ( .IN1(n3836), .IN2(n13600), .IN3(n3833), .Q(n13609) );
  AO21X1 U24458 ( .IN1(n4196), .IN2(n11434), .IN3(n4193), .Q(n11443) );
  AO21X1 U24459 ( .IN1(n3791), .IN2(n13291), .IN3(n3788), .Q(n13300) );
  AO21X1 U24460 ( .IN1(n3746), .IN2(n12982), .IN3(n3743), .Q(n12991) );
  AO21X1 U24461 ( .IN1(n4151), .IN2(n11125), .IN3(n4148), .Q(n11134) );
  AO21X1 U24462 ( .IN1(n4106), .IN2(n10815), .IN3(n4103), .Q(n10824) );
  AO21X1 U24463 ( .IN1(n3701), .IN2(n12673), .IN3(n3698), .Q(n12682) );
  AO21X1 U24464 ( .IN1(n3656), .IN2(n12364), .IN3(n3653), .Q(n12373) );
  AO21X1 U24465 ( .IN1(n4061), .IN2(n10506), .IN3(n4058), .Q(n10515) );
  AO21X1 U24466 ( .IN1(n4016), .IN2(n10196), .IN3(n4013), .Q(n10205) );
  AO21X1 U24467 ( .IN1(n3611), .IN2(n12054), .IN3(n3608), .Q(n12063) );
  AO21X1 U24468 ( .IN1(n3566), .IN2(n11744), .IN3(n3563), .Q(n11753) );
  AO21X1 U24469 ( .IN1(n3971), .IN2(n9886), .IN3(n3968), .Q(n9895) );
  AO21X1 U24470 ( .IN1(n3926), .IN2(n9575), .IN3(n3923), .Q(n9584) );
  AO21X1 U24471 ( .IN1(n4241), .IN2(n14183), .IN3(n4238), .Q(n14192) );
  NAND2X0 U24472 ( .IN1(n13880), .IN2(n13888), .QN(n13898) );
  NAND2X0 U24473 ( .IN1(n13571), .IN2(n13579), .QN(n13589) );
  NAND2X0 U24474 ( .IN1(n11405), .IN2(n11413), .QN(n11423) );
  NAND2X0 U24475 ( .IN1(n13262), .IN2(n13270), .QN(n13280) );
  NAND2X0 U24476 ( .IN1(n12953), .IN2(n12961), .QN(n12971) );
  NAND2X0 U24477 ( .IN1(n11096), .IN2(n11104), .QN(n11114) );
  NAND2X0 U24478 ( .IN1(n10786), .IN2(n10794), .QN(n10804) );
  NAND2X0 U24479 ( .IN1(n12644), .IN2(n12652), .QN(n12662) );
  NAND2X0 U24480 ( .IN1(n12335), .IN2(n12343), .QN(n12353) );
  NAND2X0 U24481 ( .IN1(n10477), .IN2(n10485), .QN(n10495) );
  NAND2X0 U24482 ( .IN1(n10167), .IN2(n10175), .QN(n10185) );
  NAND2X0 U24483 ( .IN1(n12025), .IN2(n12033), .QN(n12043) );
  NAND2X0 U24484 ( .IN1(n11715), .IN2(n11723), .QN(n11733) );
  NAND2X0 U24485 ( .IN1(n9857), .IN2(n9865), .QN(n9875) );
  NAND2X0 U24486 ( .IN1(n9546), .IN2(n9554), .QN(n9564) );
  NAND2X0 U24487 ( .IN1(n14154), .IN2(n14162), .QN(n14172) );
  AND4X1 U24488 ( .IN1(n13987), .IN2(n3400), .IN3(n18157), .IN4(n13944), .Q(
        n13992) );
  NAND3X0 U24489 ( .IN1(n13944), .IN2(n3258), .IN3(n18157), .QN(n13963) );
  NAND3X0 U24490 ( .IN1(n3382), .IN2(n3260), .IN3(n18158), .QN(n14103) );
  AND4X1 U24491 ( .IN1(n14127), .IN2(n3401), .IN3(n18158), .IN4(n3382), .Q(
        n14132) );
  AND3X1 U24492 ( .IN1(n13880), .IN2(n13883), .IN3(n3497), .Q(n13921) );
  AND3X1 U24493 ( .IN1(n13571), .IN2(n13574), .IN3(n3501), .Q(n13612) );
  AND3X1 U24494 ( .IN1(n11405), .IN2(n11408), .IN3(n3469), .Q(n11446) );
  AND3X1 U24495 ( .IN1(n13262), .IN2(n13265), .IN3(n3505), .Q(n13303) );
  AND3X1 U24496 ( .IN1(n12953), .IN2(n12956), .IN3(n3509), .Q(n12994) );
  AND3X1 U24497 ( .IN1(n11096), .IN2(n11099), .IN3(n3473), .Q(n11137) );
  AND3X1 U24498 ( .IN1(n10786), .IN2(n10789), .IN3(n3477), .Q(n10827) );
  AND3X1 U24499 ( .IN1(n12644), .IN2(n12647), .IN3(n3513), .Q(n12685) );
  AND3X1 U24500 ( .IN1(n12335), .IN2(n12338), .IN3(n3517), .Q(n12376) );
  AND3X1 U24501 ( .IN1(n10477), .IN2(n10480), .IN3(n3481), .Q(n10518) );
  AND3X1 U24502 ( .IN1(n10167), .IN2(n10170), .IN3(n3485), .Q(n10208) );
  AND3X1 U24503 ( .IN1(n12025), .IN2(n12028), .IN3(n3521), .Q(n12066) );
  AND3X1 U24504 ( .IN1(n11715), .IN2(n11718), .IN3(n3525), .Q(n11756) );
  AND3X1 U24505 ( .IN1(n9857), .IN2(n9860), .IN3(n3489), .Q(n9898) );
  AND3X1 U24506 ( .IN1(n9546), .IN2(n9549), .IN3(n3493), .Q(n9587) );
  AND3X1 U24507 ( .IN1(n14154), .IN2(n14157), .IN3(n3463), .Q(n14195) );
  AO221X1 U24508 ( .IN1(n3879), .IN2(n13921), .IN3(n3880), .IN4(n13922), .IN5(
        n13923), .Q(n13879) );
  INVX0 U24509 ( .IN(n13901), .QN(n3880) );
  AO22X1 U24510 ( .IN1(n3497), .IN2(n3882), .IN3(n13924), .IN4(n13922), .Q(
        n13923) );
  NOR2X0 U24511 ( .IN1(n3146), .IN2(n3224), .QN(n13924) );
  AO221X1 U24512 ( .IN1(n3834), .IN2(n13612), .IN3(n3835), .IN4(n13613), .IN5(
        n13614), .Q(n13570) );
  INVX0 U24513 ( .IN(n13592), .QN(n3835) );
  AO22X1 U24514 ( .IN1(n3501), .IN2(n3837), .IN3(n13615), .IN4(n13613), .Q(
        n13614) );
  NOR2X0 U24515 ( .IN1(n3152), .IN2(n3228), .QN(n13615) );
  AO221X1 U24516 ( .IN1(n4194), .IN2(n11446), .IN3(n4195), .IN4(n11447), .IN5(
        n11448), .Q(n11404) );
  INVX0 U24517 ( .IN(n11426), .QN(n4195) );
  AO22X1 U24518 ( .IN1(n3469), .IN2(n4197), .IN3(n11449), .IN4(n11447), .Q(
        n11448) );
  NOR2X0 U24519 ( .IN1(n3104), .IN2(n3196), .QN(n11449) );
  AO221X1 U24520 ( .IN1(n3789), .IN2(n13303), .IN3(n3790), .IN4(n13304), .IN5(
        n13305), .Q(n13261) );
  INVX0 U24521 ( .IN(n13283), .QN(n3790) );
  AO22X1 U24522 ( .IN1(n3505), .IN2(n3792), .IN3(n13306), .IN4(n13304), .Q(
        n13305) );
  NOR2X0 U24523 ( .IN1(n3158), .IN2(n3232), .QN(n13306) );
  AO221X1 U24524 ( .IN1(n3744), .IN2(n12994), .IN3(n3745), .IN4(n12995), .IN5(
        n12996), .Q(n12952) );
  INVX0 U24525 ( .IN(n12974), .QN(n3745) );
  AO22X1 U24526 ( .IN1(n3509), .IN2(n3747), .IN3(n12997), .IN4(n12995), .Q(
        n12996) );
  NOR2X0 U24527 ( .IN1(n3164), .IN2(n3236), .QN(n12997) );
  AO221X1 U24528 ( .IN1(n4149), .IN2(n11137), .IN3(n4150), .IN4(n11138), .IN5(
        n11139), .Q(n11095) );
  INVX0 U24529 ( .IN(n11117), .QN(n4150) );
  AO22X1 U24530 ( .IN1(n3473), .IN2(n4152), .IN3(n11140), .IN4(n11138), .Q(
        n11139) );
  NOR2X0 U24531 ( .IN1(n3110), .IN2(n3200), .QN(n11140) );
  AO221X1 U24532 ( .IN1(n4104), .IN2(n10827), .IN3(n4105), .IN4(n10828), .IN5(
        n10829), .Q(n10785) );
  INVX0 U24533 ( .IN(n10807), .QN(n4105) );
  AO22X1 U24534 ( .IN1(n3477), .IN2(n4107), .IN3(n10830), .IN4(n10828), .Q(
        n10829) );
  NOR2X0 U24535 ( .IN1(n3116), .IN2(n3204), .QN(n10830) );
  AO221X1 U24536 ( .IN1(n3699), .IN2(n12685), .IN3(n3700), .IN4(n12686), .IN5(
        n12687), .Q(n12643) );
  INVX0 U24537 ( .IN(n12665), .QN(n3700) );
  AO22X1 U24538 ( .IN1(n3513), .IN2(n3702), .IN3(n12688), .IN4(n12686), .Q(
        n12687) );
  NOR2X0 U24539 ( .IN1(n3170), .IN2(n3240), .QN(n12688) );
  AO221X1 U24540 ( .IN1(n3654), .IN2(n12376), .IN3(n3655), .IN4(n12377), .IN5(
        n12378), .Q(n12334) );
  INVX0 U24541 ( .IN(n12356), .QN(n3655) );
  AO22X1 U24542 ( .IN1(n3517), .IN2(n3657), .IN3(n12379), .IN4(n12377), .Q(
        n12378) );
  NOR2X0 U24543 ( .IN1(n3176), .IN2(n3244), .QN(n12379) );
  AO221X1 U24544 ( .IN1(n4059), .IN2(n10518), .IN3(n4060), .IN4(n10519), .IN5(
        n10520), .Q(n10476) );
  INVX0 U24545 ( .IN(n10498), .QN(n4060) );
  AO22X1 U24546 ( .IN1(n3481), .IN2(n4062), .IN3(n10521), .IN4(n10519), .Q(
        n10520) );
  NOR2X0 U24547 ( .IN1(n3122), .IN2(n3208), .QN(n10521) );
  AO221X1 U24548 ( .IN1(n4014), .IN2(n10208), .IN3(n4015), .IN4(n10209), .IN5(
        n10210), .Q(n10166) );
  INVX0 U24549 ( .IN(n10188), .QN(n4015) );
  AO22X1 U24550 ( .IN1(n3485), .IN2(n4017), .IN3(n10211), .IN4(n10209), .Q(
        n10210) );
  NOR2X0 U24551 ( .IN1(n3128), .IN2(n3212), .QN(n10211) );
  AO221X1 U24552 ( .IN1(n3609), .IN2(n12066), .IN3(n3610), .IN4(n12067), .IN5(
        n12068), .Q(n12024) );
  INVX0 U24553 ( .IN(n12046), .QN(n3610) );
  AO22X1 U24554 ( .IN1(n3521), .IN2(n3612), .IN3(n12069), .IN4(n12067), .Q(
        n12068) );
  NOR2X0 U24555 ( .IN1(n3182), .IN2(n3248), .QN(n12069) );
  AO221X1 U24556 ( .IN1(n3564), .IN2(n11756), .IN3(n3565), .IN4(n11757), .IN5(
        n11758), .Q(n11714) );
  INVX0 U24557 ( .IN(n11736), .QN(n3565) );
  AO22X1 U24558 ( .IN1(n3525), .IN2(n3567), .IN3(n11759), .IN4(n11757), .Q(
        n11758) );
  NOR2X0 U24559 ( .IN1(n3188), .IN2(n3252), .QN(n11759) );
  AO221X1 U24560 ( .IN1(n3969), .IN2(n9898), .IN3(n3970), .IN4(n9899), .IN5(
        n9900), .Q(n9856) );
  INVX0 U24561 ( .IN(n9878), .QN(n3970) );
  AO22X1 U24562 ( .IN1(n3489), .IN2(n3972), .IN3(n9901), .IN4(n9899), .Q(n9900) );
  NOR2X0 U24563 ( .IN1(n3134), .IN2(n3216), .QN(n9901) );
  AO221X1 U24564 ( .IN1(n3924), .IN2(n9587), .IN3(n3925), .IN4(n9588), .IN5(
        n9589), .Q(n9545) );
  INVX0 U24565 ( .IN(n9567), .QN(n3925) );
  AO22X1 U24566 ( .IN1(n3493), .IN2(n3927), .IN3(n9590), .IN4(n9588), .Q(n9589) );
  NOR2X0 U24567 ( .IN1(n3140), .IN2(n3220), .QN(n9590) );
  AO221X1 U24568 ( .IN1(n4239), .IN2(n14195), .IN3(n4240), .IN4(n14196), .IN5(
        n14197), .Q(n14153) );
  INVX0 U24569 ( .IN(n14175), .QN(n4240) );
  AO22X1 U24570 ( .IN1(n3463), .IN2(n4242), .IN3(n14198), .IN4(n14196), .Q(
        n14197) );
  NOR2X0 U24571 ( .IN1(n3094), .IN2(n3190), .QN(n14198) );
  OA221X1 U24572 ( .IN1(n18812), .IN2(n2833), .IN3(n14808), .IN4(n18810), 
        .IN5(n14809), .Q(n14807) );
  OA22X1 U24573 ( .IN1(n18806), .IN2(n2798), .IN3(n18803), .IN4(n2763), .Q(
        n14809) );
  OA221X1 U24574 ( .IN1(n18813), .IN2(n2832), .IN3(n14709), .IN4(n18811), 
        .IN5(n14710), .Q(n14708) );
  OA22X1 U24575 ( .IN1(n18807), .IN2(n2797), .IN3(n18804), .IN4(n2762), .Q(
        n14710) );
  OA221X1 U24576 ( .IN1(n18813), .IN2(n2831), .IN3(n14610), .IN4(n18811), 
        .IN5(n14611), .Q(n14609) );
  OA22X1 U24577 ( .IN1(n18806), .IN2(n2796), .IN3(n18804), .IN4(n2761), .Q(
        n14611) );
  OA221X1 U24578 ( .IN1(n18814), .IN2(n2830), .IN3(n14583), .IN4(n18811), 
        .IN5(n14584), .Q(n14582) );
  OA22X1 U24579 ( .IN1(n18808), .IN2(n2795), .IN3(n18805), .IN4(n2760), .Q(
        n14584) );
  OA221X1 U24580 ( .IN1(n18812), .IN2(n2829), .IN3(n14574), .IN4(n18810), 
        .IN5(n14575), .Q(n14573) );
  OA22X1 U24581 ( .IN1(n18807), .IN2(n2794), .IN3(n18803), .IN4(n2759), .Q(
        n14575) );
  OA221X1 U24582 ( .IN1(n18814), .IN2(n2828), .IN3(n14565), .IN4(n18810), 
        .IN5(n14566), .Q(n14564) );
  OA22X1 U24583 ( .IN1(n18807), .IN2(n2793), .IN3(n18804), .IN4(n2758), .Q(
        n14566) );
  OA221X1 U24584 ( .IN1(n18814), .IN2(n2827), .IN3(n14556), .IN4(n18810), 
        .IN5(n14557), .Q(n14555) );
  OA22X1 U24585 ( .IN1(n18808), .IN2(n2792), .IN3(n18805), .IN4(n2757), .Q(
        n14557) );
  OA221X1 U24586 ( .IN1(n18814), .IN2(n2826), .IN3(n14547), .IN4(n18810), 
        .IN5(n14548), .Q(n14546) );
  OA22X1 U24587 ( .IN1(n18808), .IN2(n2791), .IN3(n18805), .IN4(n2756), .Q(
        n14548) );
  OA221X1 U24588 ( .IN1(n18814), .IN2(n2825), .IN3(n14538), .IN4(n18810), 
        .IN5(n14539), .Q(n14537) );
  OA22X1 U24589 ( .IN1(n18808), .IN2(n2790), .IN3(n18805), .IN4(n2755), .Q(
        n14539) );
  OA221X1 U24590 ( .IN1(n18814), .IN2(n2824), .IN3(n14514), .IN4(n18811), 
        .IN5(n14516), .Q(n14512) );
  OA22X1 U24591 ( .IN1(n18808), .IN2(n2789), .IN3(n18805), .IN4(n2754), .Q(
        n14516) );
  OA221X1 U24592 ( .IN1(n18812), .IN2(n2823), .IN3(n14799), .IN4(n18810), 
        .IN5(n14800), .Q(n14798) );
  OA22X1 U24593 ( .IN1(n18806), .IN2(n2788), .IN3(n18803), .IN4(n2753), .Q(
        n14800) );
  OA221X1 U24594 ( .IN1(n18812), .IN2(n2822), .IN3(n14790), .IN4(n18810), 
        .IN5(n14791), .Q(n14789) );
  OA22X1 U24595 ( .IN1(n18806), .IN2(n2787), .IN3(n18803), .IN4(n2752), .Q(
        n14791) );
  OA221X1 U24596 ( .IN1(n18812), .IN2(n2821), .IN3(n14781), .IN4(n18811), 
        .IN5(n14782), .Q(n14780) );
  OA22X1 U24597 ( .IN1(n18806), .IN2(n2786), .IN3(n18803), .IN4(n2751), .Q(
        n14782) );
  OA221X1 U24598 ( .IN1(n18812), .IN2(n2820), .IN3(n14772), .IN4(n18809), 
        .IN5(n14773), .Q(n14771) );
  OA22X1 U24599 ( .IN1(n18806), .IN2(n2785), .IN3(n18804), .IN4(n2750), .Q(
        n14773) );
  OA221X1 U24600 ( .IN1(n18813), .IN2(n2819), .IN3(n14763), .IN4(n18811), 
        .IN5(n14764), .Q(n14762) );
  OA22X1 U24601 ( .IN1(n18807), .IN2(n2784), .IN3(n18804), .IN4(n2749), .Q(
        n14764) );
  OA221X1 U24602 ( .IN1(n18814), .IN2(n2818), .IN3(n14754), .IN4(n18811), 
        .IN5(n14755), .Q(n14753) );
  OA22X1 U24603 ( .IN1(n18808), .IN2(n2783), .IN3(n18804), .IN4(n2748), .Q(
        n14755) );
  OA221X1 U24604 ( .IN1(n18813), .IN2(n2817), .IN3(n18809), .IN4(n14745), 
        .IN5(n14746), .Q(n14744) );
  OA22X1 U24605 ( .IN1(n18808), .IN2(n2782), .IN3(n18804), .IN4(n2747), .Q(
        n14746) );
  OA221X1 U24606 ( .IN1(n18813), .IN2(n2816), .IN3(n18809), .IN4(n14736), 
        .IN5(n14737), .Q(n14735) );
  OA22X1 U24607 ( .IN1(n18807), .IN2(n2781), .IN3(n18805), .IN4(n2746), .Q(
        n14737) );
  OA221X1 U24608 ( .IN1(n18813), .IN2(n2815), .IN3(n18811), .IN4(n14727), 
        .IN5(n14728), .Q(n14726) );
  OA22X1 U24609 ( .IN1(n18807), .IN2(n2780), .IN3(n18805), .IN4(n2745), .Q(
        n14728) );
  OA221X1 U24610 ( .IN1(n18813), .IN2(n2814), .IN3(n18809), .IN4(n14718), 
        .IN5(n14719), .Q(n14717) );
  OA22X1 U24611 ( .IN1(n18807), .IN2(n2779), .IN3(n18803), .IN4(n2744), .Q(
        n14719) );
  OA221X1 U24612 ( .IN1(n18813), .IN2(n2813), .IN3(n18809), .IN4(n14700), 
        .IN5(n14701), .Q(n14699) );
  OA22X1 U24613 ( .IN1(n18808), .IN2(n2778), .IN3(n18805), .IN4(n2743), .Q(
        n14701) );
  OA221X1 U24614 ( .IN1(n18814), .IN2(n2812), .IN3(n18809), .IN4(n14691), 
        .IN5(n14692), .Q(n14690) );
  OA22X1 U24615 ( .IN1(n18808), .IN2(n2777), .IN3(n18803), .IN4(n2742), .Q(
        n14692) );
  OA221X1 U24616 ( .IN1(n18813), .IN2(n2811), .IN3(n18810), .IN4(n14682), 
        .IN5(n14683), .Q(n14681) );
  OA22X1 U24617 ( .IN1(n18808), .IN2(n2776), .IN3(n18804), .IN4(n2741), .Q(
        n14683) );
  OA221X1 U24618 ( .IN1(n18812), .IN2(n2810), .IN3(n18809), .IN4(n14673), 
        .IN5(n14674), .Q(n14672) );
  OA22X1 U24619 ( .IN1(n18806), .IN2(n2775), .IN3(n18804), .IN4(n2740), .Q(
        n14674) );
  OA221X1 U24620 ( .IN1(n18814), .IN2(n2809), .IN3(n18809), .IN4(n14664), 
        .IN5(n14665), .Q(n14663) );
  OA22X1 U24621 ( .IN1(n18807), .IN2(n2774), .IN3(n18804), .IN4(n2739), .Q(
        n14665) );
  OA221X1 U24622 ( .IN1(n18814), .IN2(n2808), .IN3(n18810), .IN4(n14655), 
        .IN5(n14656), .Q(n14654) );
  OA22X1 U24623 ( .IN1(n18807), .IN2(n2773), .IN3(n18803), .IN4(n2738), .Q(
        n14656) );
  OA221X1 U24624 ( .IN1(n18812), .IN2(n2807), .IN3(n18811), .IN4(n14646), 
        .IN5(n14647), .Q(n14645) );
  OA22X1 U24625 ( .IN1(n18808), .IN2(n2772), .IN3(n18803), .IN4(n2737), .Q(
        n14647) );
  OA221X1 U24626 ( .IN1(n18812), .IN2(n2806), .IN3(n18810), .IN4(n14637), 
        .IN5(n14638), .Q(n14636) );
  OA22X1 U24627 ( .IN1(n18806), .IN2(n2771), .IN3(n18804), .IN4(n2736), .Q(
        n14638) );
  OA221X1 U24628 ( .IN1(n18812), .IN2(n2805), .IN3(n18811), .IN4(n14628), 
        .IN5(n14629), .Q(n14627) );
  OA22X1 U24629 ( .IN1(n18806), .IN2(n2770), .IN3(n18805), .IN4(n2735), .Q(
        n14629) );
  OA221X1 U24630 ( .IN1(n18813), .IN2(n2804), .IN3(n18809), .IN4(n14619), 
        .IN5(n14620), .Q(n14618) );
  OA22X1 U24631 ( .IN1(n18806), .IN2(n2769), .IN3(n18805), .IN4(n2734), .Q(
        n14620) );
  OA221X1 U24632 ( .IN1(n18813), .IN2(n2803), .IN3(n18809), .IN4(n14601), 
        .IN5(n14602), .Q(n14600) );
  OA22X1 U24633 ( .IN1(n18806), .IN2(n2768), .IN3(n18803), .IN4(n2733), .Q(
        n14602) );
  OA221X1 U24634 ( .IN1(n18812), .IN2(n2802), .IN3(n18809), .IN4(n14592), 
        .IN5(n14593), .Q(n14591) );
  OA22X1 U24635 ( .IN1(n18807), .IN2(n2767), .IN3(n18803), .IN4(n2732), .Q(
        n14593) );
  OA221X1 U24636 ( .IN1(n18764), .IN2(n2833), .IN3(n14808), .IN4(n18762), 
        .IN5(n15160), .Q(n15159) );
  OA22X1 U24637 ( .IN1(n18758), .IN2(n2798), .IN3(n18755), .IN4(n2763), .Q(
        n15160) );
  OA221X1 U24638 ( .IN1(n18766), .IN2(n2832), .IN3(n14709), .IN4(n18763), 
        .IN5(n15072), .Q(n15071) );
  OA22X1 U24639 ( .IN1(n18758), .IN2(n2797), .IN3(n18756), .IN4(n2762), .Q(
        n15072) );
  OA221X1 U24640 ( .IN1(n18764), .IN2(n2831), .IN3(n14610), .IN4(n18763), 
        .IN5(n14984), .Q(n14983) );
  OA22X1 U24641 ( .IN1(n18760), .IN2(n2796), .IN3(n18755), .IN4(n2761), .Q(
        n14984) );
  OA221X1 U24642 ( .IN1(n18764), .IN2(n2830), .IN3(n14583), .IN4(n18763), 
        .IN5(n14960), .Q(n14959) );
  OA22X1 U24643 ( .IN1(n18758), .IN2(n2795), .IN3(n14900), .IN4(n2760), .Q(
        n14960) );
  OA221X1 U24644 ( .IN1(n18766), .IN2(n2829), .IN3(n14574), .IN4(n18762), 
        .IN5(n14952), .Q(n14951) );
  OA22X1 U24645 ( .IN1(n18758), .IN2(n2794), .IN3(n14900), .IN4(n2759), .Q(
        n14952) );
  OA221X1 U24646 ( .IN1(n18765), .IN2(n2828), .IN3(n14565), .IN4(n18762), 
        .IN5(n14944), .Q(n14943) );
  OA22X1 U24647 ( .IN1(n18760), .IN2(n2793), .IN3(n14900), .IN4(n2758), .Q(
        n14944) );
  OA221X1 U24648 ( .IN1(n18766), .IN2(n2827), .IN3(n14556), .IN4(n18762), 
        .IN5(n14936), .Q(n14935) );
  OA22X1 U24649 ( .IN1(n18760), .IN2(n2792), .IN3(n18756), .IN4(n2757), .Q(
        n14936) );
  OA221X1 U24650 ( .IN1(n18766), .IN2(n2826), .IN3(n14547), .IN4(n18762), 
        .IN5(n14928), .Q(n14927) );
  OA22X1 U24651 ( .IN1(n18759), .IN2(n2791), .IN3(n18756), .IN4(n2756), .Q(
        n14928) );
  OA221X1 U24652 ( .IN1(n18766), .IN2(n2825), .IN3(n14538), .IN4(n18762), 
        .IN5(n14920), .Q(n14919) );
  OA22X1 U24653 ( .IN1(n18758), .IN2(n2790), .IN3(n18756), .IN4(n2755), .Q(
        n14920) );
  OA221X1 U24654 ( .IN1(n18766), .IN2(n2824), .IN3(n14514), .IN4(n18763), 
        .IN5(n14898), .Q(n14895) );
  OA22X1 U24655 ( .IN1(n18760), .IN2(n2789), .IN3(n18756), .IN4(n2754), .Q(
        n14898) );
  OA221X1 U24656 ( .IN1(n18764), .IN2(n2823), .IN3(n14799), .IN4(n18762), 
        .IN5(n15152), .Q(n15151) );
  OA22X1 U24657 ( .IN1(n18758), .IN2(n2788), .IN3(n18755), .IN4(n2753), .Q(
        n15152) );
  OA221X1 U24658 ( .IN1(n18764), .IN2(n2822), .IN3(n14790), .IN4(n18762), 
        .IN5(n15144), .Q(n15143) );
  OA22X1 U24659 ( .IN1(n18758), .IN2(n2787), .IN3(n18755), .IN4(n2752), .Q(
        n15144) );
  OA221X1 U24660 ( .IN1(n18764), .IN2(n2821), .IN3(n14781), .IN4(n18763), 
        .IN5(n15136), .Q(n15135) );
  OA22X1 U24661 ( .IN1(n18758), .IN2(n2786), .IN3(n18755), .IN4(n2751), .Q(
        n15136) );
  OA221X1 U24662 ( .IN1(n18765), .IN2(n2820), .IN3(n14772), .IN4(n18761), 
        .IN5(n15128), .Q(n15127) );
  OA22X1 U24663 ( .IN1(n18759), .IN2(n2785), .IN3(n14900), .IN4(n2750), .Q(
        n15128) );
  OA221X1 U24664 ( .IN1(n18765), .IN2(n2819), .IN3(n14763), .IN4(n18763), 
        .IN5(n15120), .Q(n15119) );
  OA22X1 U24665 ( .IN1(n18759), .IN2(n2784), .IN3(n14900), .IN4(n2749), .Q(
        n15120) );
  OA221X1 U24666 ( .IN1(n18765), .IN2(n2818), .IN3(n14754), .IN4(n18763), 
        .IN5(n15112), .Q(n15111) );
  OA22X1 U24667 ( .IN1(n18759), .IN2(n2783), .IN3(n14900), .IN4(n2748), .Q(
        n15112) );
  OA221X1 U24668 ( .IN1(n18765), .IN2(n2817), .IN3(n18761), .IN4(n14745), 
        .IN5(n15104), .Q(n15103) );
  OA22X1 U24669 ( .IN1(n18759), .IN2(n2782), .IN3(n18756), .IN4(n2747), .Q(
        n15104) );
  OA221X1 U24670 ( .IN1(n18765), .IN2(n2816), .IN3(n18761), .IN4(n14736), 
        .IN5(n15096), .Q(n15095) );
  OA22X1 U24671 ( .IN1(n18759), .IN2(n2781), .IN3(n18756), .IN4(n2746), .Q(
        n15096) );
  OA221X1 U24672 ( .IN1(n18765), .IN2(n2815), .IN3(n18763), .IN4(n14727), 
        .IN5(n15088), .Q(n15087) );
  OA22X1 U24673 ( .IN1(n18760), .IN2(n2780), .IN3(n14900), .IN4(n2745), .Q(
        n15088) );
  OA221X1 U24674 ( .IN1(n18766), .IN2(n2814), .IN3(n18761), .IN4(n14718), 
        .IN5(n15080), .Q(n15079) );
  OA22X1 U24675 ( .IN1(n18758), .IN2(n2779), .IN3(n18756), .IN4(n2744), .Q(
        n15080) );
  OA221X1 U24676 ( .IN1(n18764), .IN2(n2813), .IN3(n18761), .IN4(n14700), 
        .IN5(n15064), .Q(n15063) );
  OA22X1 U24677 ( .IN1(n18760), .IN2(n2778), .IN3(n14900), .IN4(n2743), .Q(
        n15064) );
  OA221X1 U24678 ( .IN1(n18765), .IN2(n2812), .IN3(n18761), .IN4(n14691), 
        .IN5(n15056), .Q(n15055) );
  OA22X1 U24679 ( .IN1(n18760), .IN2(n2777), .IN3(n14900), .IN4(n2742), .Q(
        n15056) );
  OA221X1 U24680 ( .IN1(n18764), .IN2(n2811), .IN3(n18762), .IN4(n14682), 
        .IN5(n15048), .Q(n15047) );
  OA22X1 U24681 ( .IN1(n18760), .IN2(n2776), .IN3(n18755), .IN4(n2741), .Q(
        n15048) );
  OA221X1 U24682 ( .IN1(n18766), .IN2(n2810), .IN3(n18761), .IN4(n14673), 
        .IN5(n15040), .Q(n15039) );
  OA22X1 U24683 ( .IN1(n18760), .IN2(n2775), .IN3(n14900), .IN4(n2740), .Q(
        n15040) );
  OA221X1 U24684 ( .IN1(n18766), .IN2(n2809), .IN3(n18761), .IN4(n14664), 
        .IN5(n15032), .Q(n15031) );
  OA22X1 U24685 ( .IN1(n18760), .IN2(n2774), .IN3(n18755), .IN4(n2739), .Q(
        n15032) );
  OA221X1 U24686 ( .IN1(n18766), .IN2(n2808), .IN3(n18762), .IN4(n14655), 
        .IN5(n15024), .Q(n15023) );
  OA22X1 U24687 ( .IN1(n18759), .IN2(n2773), .IN3(n18755), .IN4(n2738), .Q(
        n15024) );
  OA221X1 U24688 ( .IN1(n18764), .IN2(n2807), .IN3(n18763), .IN4(n14646), 
        .IN5(n15016), .Q(n15015) );
  OA22X1 U24689 ( .IN1(n18760), .IN2(n2772), .IN3(n14900), .IN4(n2737), .Q(
        n15016) );
  OA221X1 U24690 ( .IN1(n18764), .IN2(n2806), .IN3(n18762), .IN4(n14637), 
        .IN5(n15008), .Q(n15007) );
  OA22X1 U24691 ( .IN1(n18759), .IN2(n2771), .IN3(n18755), .IN4(n2736), .Q(
        n15008) );
  OA221X1 U24692 ( .IN1(n18765), .IN2(n2805), .IN3(n18763), .IN4(n14628), 
        .IN5(n15000), .Q(n14999) );
  OA22X1 U24693 ( .IN1(n18759), .IN2(n2770), .IN3(n14900), .IN4(n2735), .Q(
        n15000) );
  OA221X1 U24694 ( .IN1(n18764), .IN2(n2804), .IN3(n18761), .IN4(n14619), 
        .IN5(n14992), .Q(n14991) );
  OA22X1 U24695 ( .IN1(n18758), .IN2(n2769), .IN3(n18755), .IN4(n2734), .Q(
        n14992) );
  OA221X1 U24696 ( .IN1(n18766), .IN2(n2803), .IN3(n18761), .IN4(n14601), 
        .IN5(n14976), .Q(n14975) );
  OA22X1 U24697 ( .IN1(n18758), .IN2(n2768), .IN3(n18756), .IN4(n2733), .Q(
        n14976) );
  OA221X1 U24698 ( .IN1(n18765), .IN2(n2802), .IN3(n18761), .IN4(n14592), 
        .IN5(n14968), .Q(n14967) );
  OA22X1 U24699 ( .IN1(n18759), .IN2(n2767), .IN3(n18756), .IN4(n2732), .Q(
        n14968) );
  OA221X1 U24700 ( .IN1(n18716), .IN2(n2833), .IN3(n14808), .IN4(n18714), 
        .IN5(n15465), .Q(n15464) );
  OA22X1 U24701 ( .IN1(n18710), .IN2(n2798), .IN3(n18707), .IN4(n2763), .Q(
        n15465) );
  OA221X1 U24702 ( .IN1(n18717), .IN2(n2832), .IN3(n14709), .IN4(n18715), 
        .IN5(n15377), .Q(n15376) );
  OA22X1 U24703 ( .IN1(n18711), .IN2(n2797), .IN3(n18708), .IN4(n2762), .Q(
        n15377) );
  OA221X1 U24704 ( .IN1(n18717), .IN2(n2831), .IN3(n14610), .IN4(n18715), 
        .IN5(n15289), .Q(n15288) );
  OA22X1 U24705 ( .IN1(n18710), .IN2(n2796), .IN3(n18708), .IN4(n2761), .Q(
        n15289) );
  OA221X1 U24706 ( .IN1(n18718), .IN2(n2830), .IN3(n14583), .IN4(n18715), 
        .IN5(n15265), .Q(n15264) );
  OA22X1 U24707 ( .IN1(n18712), .IN2(n2795), .IN3(n18709), .IN4(n2760), .Q(
        n15265) );
  OA221X1 U24708 ( .IN1(n18716), .IN2(n2829), .IN3(n14574), .IN4(n18714), 
        .IN5(n15257), .Q(n15256) );
  OA22X1 U24709 ( .IN1(n18711), .IN2(n2794), .IN3(n18707), .IN4(n2759), .Q(
        n15257) );
  OA221X1 U24710 ( .IN1(n18718), .IN2(n2828), .IN3(n14565), .IN4(n18714), 
        .IN5(n15249), .Q(n15248) );
  OA22X1 U24711 ( .IN1(n18711), .IN2(n2793), .IN3(n18708), .IN4(n2758), .Q(
        n15249) );
  OA221X1 U24712 ( .IN1(n18718), .IN2(n2827), .IN3(n14556), .IN4(n18714), 
        .IN5(n15241), .Q(n15240) );
  OA22X1 U24713 ( .IN1(n18712), .IN2(n2792), .IN3(n18709), .IN4(n2757), .Q(
        n15241) );
  OA221X1 U24714 ( .IN1(n18718), .IN2(n2826), .IN3(n14547), .IN4(n18714), 
        .IN5(n15233), .Q(n15232) );
  OA22X1 U24715 ( .IN1(n18712), .IN2(n2791), .IN3(n18709), .IN4(n2756), .Q(
        n15233) );
  OA221X1 U24716 ( .IN1(n18718), .IN2(n2825), .IN3(n14538), .IN4(n18714), 
        .IN5(n15225), .Q(n15224) );
  OA22X1 U24717 ( .IN1(n18712), .IN2(n2790), .IN3(n18709), .IN4(n2755), .Q(
        n15225) );
  OA221X1 U24718 ( .IN1(n18718), .IN2(n2824), .IN3(n14514), .IN4(n18715), 
        .IN5(n15203), .Q(n15200) );
  OA22X1 U24719 ( .IN1(n18712), .IN2(n2789), .IN3(n18709), .IN4(n2754), .Q(
        n15203) );
  OA221X1 U24720 ( .IN1(n18716), .IN2(n2823), .IN3(n14799), .IN4(n18714), 
        .IN5(n15457), .Q(n15456) );
  OA22X1 U24721 ( .IN1(n18710), .IN2(n2788), .IN3(n18707), .IN4(n2753), .Q(
        n15457) );
  OA221X1 U24722 ( .IN1(n18716), .IN2(n2822), .IN3(n14790), .IN4(n18714), 
        .IN5(n15449), .Q(n15448) );
  OA22X1 U24723 ( .IN1(n18710), .IN2(n2787), .IN3(n18707), .IN4(n2752), .Q(
        n15449) );
  OA221X1 U24724 ( .IN1(n18716), .IN2(n2821), .IN3(n14781), .IN4(n18715), 
        .IN5(n15441), .Q(n15440) );
  OA22X1 U24725 ( .IN1(n18710), .IN2(n2786), .IN3(n18707), .IN4(n2751), .Q(
        n15441) );
  OA221X1 U24726 ( .IN1(n18716), .IN2(n2820), .IN3(n14772), .IN4(n18713), 
        .IN5(n15433), .Q(n15432) );
  OA22X1 U24727 ( .IN1(n18710), .IN2(n2785), .IN3(n18708), .IN4(n2750), .Q(
        n15433) );
  OA221X1 U24728 ( .IN1(n18717), .IN2(n2819), .IN3(n14763), .IN4(n18715), 
        .IN5(n15425), .Q(n15424) );
  OA22X1 U24729 ( .IN1(n18711), .IN2(n2784), .IN3(n18708), .IN4(n2749), .Q(
        n15425) );
  OA221X1 U24730 ( .IN1(n18718), .IN2(n2818), .IN3(n14754), .IN4(n18715), 
        .IN5(n15417), .Q(n15416) );
  OA22X1 U24731 ( .IN1(n18712), .IN2(n2783), .IN3(n18708), .IN4(n2748), .Q(
        n15417) );
  OA221X1 U24732 ( .IN1(n18717), .IN2(n2817), .IN3(n18713), .IN4(n14745), 
        .IN5(n15409), .Q(n15408) );
  OA22X1 U24733 ( .IN1(n18712), .IN2(n2782), .IN3(n18708), .IN4(n2747), .Q(
        n15409) );
  OA221X1 U24734 ( .IN1(n18717), .IN2(n2816), .IN3(n18713), .IN4(n14736), 
        .IN5(n15401), .Q(n15400) );
  OA22X1 U24735 ( .IN1(n18711), .IN2(n2781), .IN3(n18709), .IN4(n2746), .Q(
        n15401) );
  OA221X1 U24736 ( .IN1(n18717), .IN2(n2815), .IN3(n18715), .IN4(n14727), 
        .IN5(n15393), .Q(n15392) );
  OA22X1 U24737 ( .IN1(n18711), .IN2(n2780), .IN3(n18709), .IN4(n2745), .Q(
        n15393) );
  OA221X1 U24738 ( .IN1(n18717), .IN2(n2814), .IN3(n18713), .IN4(n14718), 
        .IN5(n15385), .Q(n15384) );
  OA22X1 U24739 ( .IN1(n18711), .IN2(n2779), .IN3(n18707), .IN4(n2744), .Q(
        n15385) );
  OA221X1 U24740 ( .IN1(n18717), .IN2(n2813), .IN3(n18713), .IN4(n14700), 
        .IN5(n15369), .Q(n15368) );
  OA22X1 U24741 ( .IN1(n18712), .IN2(n2778), .IN3(n18709), .IN4(n2743), .Q(
        n15369) );
  OA221X1 U24742 ( .IN1(n18718), .IN2(n2812), .IN3(n18713), .IN4(n14691), 
        .IN5(n15361), .Q(n15360) );
  OA22X1 U24743 ( .IN1(n18712), .IN2(n2777), .IN3(n18707), .IN4(n2742), .Q(
        n15361) );
  OA221X1 U24744 ( .IN1(n18717), .IN2(n2811), .IN3(n18714), .IN4(n14682), 
        .IN5(n15353), .Q(n15352) );
  OA22X1 U24745 ( .IN1(n18712), .IN2(n2776), .IN3(n18708), .IN4(n2741), .Q(
        n15353) );
  OA221X1 U24746 ( .IN1(n18716), .IN2(n2810), .IN3(n18713), .IN4(n14673), 
        .IN5(n15345), .Q(n15344) );
  OA22X1 U24747 ( .IN1(n18710), .IN2(n2775), .IN3(n18708), .IN4(n2740), .Q(
        n15345) );
  OA221X1 U24748 ( .IN1(n18718), .IN2(n2809), .IN3(n18713), .IN4(n14664), 
        .IN5(n15337), .Q(n15336) );
  OA22X1 U24749 ( .IN1(n18711), .IN2(n2774), .IN3(n18708), .IN4(n2739), .Q(
        n15337) );
  OA221X1 U24750 ( .IN1(n18718), .IN2(n2808), .IN3(n18714), .IN4(n14655), 
        .IN5(n15329), .Q(n15328) );
  OA22X1 U24751 ( .IN1(n18711), .IN2(n2773), .IN3(n18707), .IN4(n2738), .Q(
        n15329) );
  OA221X1 U24752 ( .IN1(n18716), .IN2(n2807), .IN3(n18715), .IN4(n14646), 
        .IN5(n15321), .Q(n15320) );
  OA22X1 U24753 ( .IN1(n18712), .IN2(n2772), .IN3(n18707), .IN4(n2737), .Q(
        n15321) );
  OA221X1 U24754 ( .IN1(n18716), .IN2(n2806), .IN3(n18714), .IN4(n14637), 
        .IN5(n15313), .Q(n15312) );
  OA22X1 U24755 ( .IN1(n18710), .IN2(n2771), .IN3(n18708), .IN4(n2736), .Q(
        n15313) );
  OA221X1 U24756 ( .IN1(n18716), .IN2(n2805), .IN3(n18715), .IN4(n14628), 
        .IN5(n15305), .Q(n15304) );
  OA22X1 U24757 ( .IN1(n18710), .IN2(n2770), .IN3(n18709), .IN4(n2735), .Q(
        n15305) );
  OA221X1 U24758 ( .IN1(n18717), .IN2(n2804), .IN3(n18713), .IN4(n14619), 
        .IN5(n15297), .Q(n15296) );
  OA22X1 U24759 ( .IN1(n18710), .IN2(n2769), .IN3(n18709), .IN4(n2734), .Q(
        n15297) );
  OA221X1 U24760 ( .IN1(n18717), .IN2(n2803), .IN3(n18713), .IN4(n14601), 
        .IN5(n15281), .Q(n15280) );
  OA22X1 U24761 ( .IN1(n18710), .IN2(n2768), .IN3(n18707), .IN4(n2733), .Q(
        n15281) );
  OA221X1 U24762 ( .IN1(n18716), .IN2(n2802), .IN3(n18713), .IN4(n14592), 
        .IN5(n15273), .Q(n15272) );
  OA22X1 U24763 ( .IN1(n18711), .IN2(n2767), .IN3(n18707), .IN4(n2732), .Q(
        n15273) );
  OA221X1 U24764 ( .IN1(n18668), .IN2(n2833), .IN3(n14808), .IN4(n18666), 
        .IN5(n15770), .Q(n15769) );
  OA22X1 U24765 ( .IN1(n18662), .IN2(n2798), .IN3(n18659), .IN4(n2763), .Q(
        n15770) );
  OA221X1 U24766 ( .IN1(n18670), .IN2(n2832), .IN3(n14709), .IN4(n18667), 
        .IN5(n15682), .Q(n15681) );
  OA22X1 U24767 ( .IN1(n18662), .IN2(n2797), .IN3(n18660), .IN4(n2762), .Q(
        n15682) );
  OA221X1 U24768 ( .IN1(n18668), .IN2(n2831), .IN3(n14610), .IN4(n18667), 
        .IN5(n15594), .Q(n15593) );
  OA22X1 U24769 ( .IN1(n18664), .IN2(n2796), .IN3(n18659), .IN4(n2761), .Q(
        n15594) );
  OA221X1 U24770 ( .IN1(n18668), .IN2(n2830), .IN3(n14583), .IN4(n18667), 
        .IN5(n15570), .Q(n15569) );
  OA22X1 U24771 ( .IN1(n18662), .IN2(n2795), .IN3(n15510), .IN4(n2760), .Q(
        n15570) );
  OA221X1 U24772 ( .IN1(n18670), .IN2(n2829), .IN3(n14574), .IN4(n18666), 
        .IN5(n15562), .Q(n15561) );
  OA22X1 U24773 ( .IN1(n18662), .IN2(n2794), .IN3(n15510), .IN4(n2759), .Q(
        n15562) );
  OA221X1 U24774 ( .IN1(n18669), .IN2(n2828), .IN3(n14565), .IN4(n18666), 
        .IN5(n15554), .Q(n15553) );
  OA22X1 U24775 ( .IN1(n18664), .IN2(n2793), .IN3(n15510), .IN4(n2758), .Q(
        n15554) );
  OA221X1 U24776 ( .IN1(n18670), .IN2(n2827), .IN3(n14556), .IN4(n18666), 
        .IN5(n15546), .Q(n15545) );
  OA22X1 U24777 ( .IN1(n18664), .IN2(n2792), .IN3(n18660), .IN4(n2757), .Q(
        n15546) );
  OA221X1 U24778 ( .IN1(n18670), .IN2(n2826), .IN3(n14547), .IN4(n18666), 
        .IN5(n15538), .Q(n15537) );
  OA22X1 U24779 ( .IN1(n18663), .IN2(n2791), .IN3(n18660), .IN4(n2756), .Q(
        n15538) );
  OA221X1 U24780 ( .IN1(n18670), .IN2(n2825), .IN3(n14538), .IN4(n18666), 
        .IN5(n15530), .Q(n15529) );
  OA22X1 U24781 ( .IN1(n18662), .IN2(n2790), .IN3(n18660), .IN4(n2755), .Q(
        n15530) );
  OA221X1 U24782 ( .IN1(n18670), .IN2(n2824), .IN3(n14514), .IN4(n18667), 
        .IN5(n15508), .Q(n15505) );
  OA22X1 U24783 ( .IN1(n18664), .IN2(n2789), .IN3(n18660), .IN4(n2754), .Q(
        n15508) );
  OA221X1 U24784 ( .IN1(n18668), .IN2(n2823), .IN3(n14799), .IN4(n18666), 
        .IN5(n15762), .Q(n15761) );
  OA22X1 U24785 ( .IN1(n18662), .IN2(n2788), .IN3(n18659), .IN4(n2753), .Q(
        n15762) );
  OA221X1 U24786 ( .IN1(n18668), .IN2(n2822), .IN3(n14790), .IN4(n18666), 
        .IN5(n15754), .Q(n15753) );
  OA22X1 U24787 ( .IN1(n18662), .IN2(n2787), .IN3(n18659), .IN4(n2752), .Q(
        n15754) );
  OA221X1 U24788 ( .IN1(n18668), .IN2(n2821), .IN3(n14781), .IN4(n18667), 
        .IN5(n15746), .Q(n15745) );
  OA22X1 U24789 ( .IN1(n18662), .IN2(n2786), .IN3(n18659), .IN4(n2751), .Q(
        n15746) );
  OA221X1 U24790 ( .IN1(n18669), .IN2(n2820), .IN3(n14772), .IN4(n18665), 
        .IN5(n15738), .Q(n15737) );
  OA22X1 U24791 ( .IN1(n18663), .IN2(n2785), .IN3(n15510), .IN4(n2750), .Q(
        n15738) );
  OA221X1 U24792 ( .IN1(n18669), .IN2(n2819), .IN3(n14763), .IN4(n18667), 
        .IN5(n15730), .Q(n15729) );
  OA22X1 U24793 ( .IN1(n18663), .IN2(n2784), .IN3(n15510), .IN4(n2749), .Q(
        n15730) );
  OA221X1 U24794 ( .IN1(n18669), .IN2(n2818), .IN3(n14754), .IN4(n18667), 
        .IN5(n15722), .Q(n15721) );
  OA22X1 U24795 ( .IN1(n18663), .IN2(n2783), .IN3(n15510), .IN4(n2748), .Q(
        n15722) );
  OA221X1 U24796 ( .IN1(n18669), .IN2(n2817), .IN3(n18665), .IN4(n14745), 
        .IN5(n15714), .Q(n15713) );
  OA22X1 U24797 ( .IN1(n18663), .IN2(n2782), .IN3(n18660), .IN4(n2747), .Q(
        n15714) );
  OA221X1 U24798 ( .IN1(n18669), .IN2(n2816), .IN3(n18665), .IN4(n14736), 
        .IN5(n15706), .Q(n15705) );
  OA22X1 U24799 ( .IN1(n18663), .IN2(n2781), .IN3(n18660), .IN4(n2746), .Q(
        n15706) );
  OA221X1 U24800 ( .IN1(n18669), .IN2(n2815), .IN3(n18667), .IN4(n14727), 
        .IN5(n15698), .Q(n15697) );
  OA22X1 U24801 ( .IN1(n18664), .IN2(n2780), .IN3(n15510), .IN4(n2745), .Q(
        n15698) );
  OA221X1 U24802 ( .IN1(n18670), .IN2(n2814), .IN3(n18665), .IN4(n14718), 
        .IN5(n15690), .Q(n15689) );
  OA22X1 U24803 ( .IN1(n18662), .IN2(n2779), .IN3(n18660), .IN4(n2744), .Q(
        n15690) );
  OA221X1 U24804 ( .IN1(n18668), .IN2(n2813), .IN3(n18665), .IN4(n14700), 
        .IN5(n15674), .Q(n15673) );
  OA22X1 U24805 ( .IN1(n18664), .IN2(n2778), .IN3(n15510), .IN4(n2743), .Q(
        n15674) );
  OA221X1 U24806 ( .IN1(n18669), .IN2(n2812), .IN3(n18665), .IN4(n14691), 
        .IN5(n15666), .Q(n15665) );
  OA22X1 U24807 ( .IN1(n18664), .IN2(n2777), .IN3(n15510), .IN4(n2742), .Q(
        n15666) );
  OA221X1 U24808 ( .IN1(n18668), .IN2(n2811), .IN3(n18666), .IN4(n14682), 
        .IN5(n15658), .Q(n15657) );
  OA22X1 U24809 ( .IN1(n18664), .IN2(n2776), .IN3(n18659), .IN4(n2741), .Q(
        n15658) );
  OA221X1 U24810 ( .IN1(n18670), .IN2(n2810), .IN3(n18665), .IN4(n14673), 
        .IN5(n15650), .Q(n15649) );
  OA22X1 U24811 ( .IN1(n18664), .IN2(n2775), .IN3(n15510), .IN4(n2740), .Q(
        n15650) );
  OA221X1 U24812 ( .IN1(n18670), .IN2(n2809), .IN3(n18665), .IN4(n14664), 
        .IN5(n15642), .Q(n15641) );
  OA22X1 U24813 ( .IN1(n18664), .IN2(n2774), .IN3(n18659), .IN4(n2739), .Q(
        n15642) );
  OA221X1 U24814 ( .IN1(n18670), .IN2(n2808), .IN3(n18666), .IN4(n14655), 
        .IN5(n15634), .Q(n15633) );
  OA22X1 U24815 ( .IN1(n18663), .IN2(n2773), .IN3(n18659), .IN4(n2738), .Q(
        n15634) );
  OA221X1 U24816 ( .IN1(n18668), .IN2(n2807), .IN3(n18667), .IN4(n14646), 
        .IN5(n15626), .Q(n15625) );
  OA22X1 U24817 ( .IN1(n18664), .IN2(n2772), .IN3(n15510), .IN4(n2737), .Q(
        n15626) );
  OA221X1 U24818 ( .IN1(n18668), .IN2(n2806), .IN3(n18666), .IN4(n14637), 
        .IN5(n15618), .Q(n15617) );
  OA22X1 U24819 ( .IN1(n18663), .IN2(n2771), .IN3(n18659), .IN4(n2736), .Q(
        n15618) );
  OA221X1 U24820 ( .IN1(n18669), .IN2(n2805), .IN3(n18667), .IN4(n14628), 
        .IN5(n15610), .Q(n15609) );
  OA22X1 U24821 ( .IN1(n18663), .IN2(n2770), .IN3(n15510), .IN4(n2735), .Q(
        n15610) );
  OA221X1 U24822 ( .IN1(n18668), .IN2(n2804), .IN3(n18665), .IN4(n14619), 
        .IN5(n15602), .Q(n15601) );
  OA22X1 U24823 ( .IN1(n18662), .IN2(n2769), .IN3(n18659), .IN4(n2734), .Q(
        n15602) );
  OA221X1 U24824 ( .IN1(n18670), .IN2(n2803), .IN3(n18665), .IN4(n14601), 
        .IN5(n15586), .Q(n15585) );
  OA22X1 U24825 ( .IN1(n18662), .IN2(n2768), .IN3(n18660), .IN4(n2733), .Q(
        n15586) );
  OA221X1 U24826 ( .IN1(n18669), .IN2(n2802), .IN3(n18665), .IN4(n14592), 
        .IN5(n15578), .Q(n15577) );
  OA22X1 U24827 ( .IN1(n18663), .IN2(n2767), .IN3(n18660), .IN4(n2732), .Q(
        n15578) );
  OA221X1 U24828 ( .IN1(n18620), .IN2(n2833), .IN3(n14808), .IN4(n18618), 
        .IN5(n16075), .Q(n16074) );
  OA22X1 U24829 ( .IN1(n18614), .IN2(n2798), .IN3(n18611), .IN4(n2763), .Q(
        n16075) );
  OA221X1 U24830 ( .IN1(n18621), .IN2(n2832), .IN3(n14709), .IN4(n18619), 
        .IN5(n15987), .Q(n15986) );
  OA22X1 U24831 ( .IN1(n18615), .IN2(n2797), .IN3(n18612), .IN4(n2762), .Q(
        n15987) );
  OA221X1 U24832 ( .IN1(n18621), .IN2(n2831), .IN3(n14610), .IN4(n18619), 
        .IN5(n15899), .Q(n15898) );
  OA22X1 U24833 ( .IN1(n18614), .IN2(n2796), .IN3(n18612), .IN4(n2761), .Q(
        n15899) );
  OA221X1 U24834 ( .IN1(n18622), .IN2(n2830), .IN3(n14583), .IN4(n18619), 
        .IN5(n15875), .Q(n15874) );
  OA22X1 U24835 ( .IN1(n18616), .IN2(n2795), .IN3(n18613), .IN4(n2760), .Q(
        n15875) );
  OA221X1 U24836 ( .IN1(n18620), .IN2(n2829), .IN3(n14574), .IN4(n18618), 
        .IN5(n15867), .Q(n15866) );
  OA22X1 U24837 ( .IN1(n18615), .IN2(n2794), .IN3(n18611), .IN4(n2759), .Q(
        n15867) );
  OA221X1 U24838 ( .IN1(n18622), .IN2(n2828), .IN3(n14565), .IN4(n18618), 
        .IN5(n15859), .Q(n15858) );
  OA22X1 U24839 ( .IN1(n18615), .IN2(n2793), .IN3(n18612), .IN4(n2758), .Q(
        n15859) );
  OA221X1 U24840 ( .IN1(n18622), .IN2(n2827), .IN3(n14556), .IN4(n18618), 
        .IN5(n15851), .Q(n15850) );
  OA22X1 U24841 ( .IN1(n18616), .IN2(n2792), .IN3(n18613), .IN4(n2757), .Q(
        n15851) );
  OA221X1 U24842 ( .IN1(n18622), .IN2(n2826), .IN3(n14547), .IN4(n18618), 
        .IN5(n15843), .Q(n15842) );
  OA22X1 U24843 ( .IN1(n18616), .IN2(n2791), .IN3(n18613), .IN4(n2756), .Q(
        n15843) );
  OA221X1 U24844 ( .IN1(n18622), .IN2(n2825), .IN3(n14538), .IN4(n18618), 
        .IN5(n15835), .Q(n15834) );
  OA22X1 U24845 ( .IN1(n18616), .IN2(n2790), .IN3(n18613), .IN4(n2755), .Q(
        n15835) );
  OA221X1 U24846 ( .IN1(n18622), .IN2(n2824), .IN3(n14514), .IN4(n18619), 
        .IN5(n15813), .Q(n15810) );
  OA22X1 U24847 ( .IN1(n18616), .IN2(n2789), .IN3(n18613), .IN4(n2754), .Q(
        n15813) );
  OA221X1 U24848 ( .IN1(n18620), .IN2(n2823), .IN3(n14799), .IN4(n18618), 
        .IN5(n16067), .Q(n16066) );
  OA22X1 U24849 ( .IN1(n18614), .IN2(n2788), .IN3(n18611), .IN4(n2753), .Q(
        n16067) );
  OA221X1 U24850 ( .IN1(n18620), .IN2(n2822), .IN3(n14790), .IN4(n18618), 
        .IN5(n16059), .Q(n16058) );
  OA22X1 U24851 ( .IN1(n18614), .IN2(n2787), .IN3(n18611), .IN4(n2752), .Q(
        n16059) );
  OA221X1 U24852 ( .IN1(n18620), .IN2(n2821), .IN3(n14781), .IN4(n18619), 
        .IN5(n16051), .Q(n16050) );
  OA22X1 U24853 ( .IN1(n18614), .IN2(n2786), .IN3(n18611), .IN4(n2751), .Q(
        n16051) );
  OA221X1 U24854 ( .IN1(n18620), .IN2(n2820), .IN3(n14772), .IN4(n18617), 
        .IN5(n16043), .Q(n16042) );
  OA22X1 U24855 ( .IN1(n18614), .IN2(n2785), .IN3(n18612), .IN4(n2750), .Q(
        n16043) );
  OA221X1 U24856 ( .IN1(n18621), .IN2(n2819), .IN3(n14763), .IN4(n18619), 
        .IN5(n16035), .Q(n16034) );
  OA22X1 U24857 ( .IN1(n18615), .IN2(n2784), .IN3(n18612), .IN4(n2749), .Q(
        n16035) );
  OA221X1 U24858 ( .IN1(n18622), .IN2(n2818), .IN3(n14754), .IN4(n18619), 
        .IN5(n16027), .Q(n16026) );
  OA22X1 U24859 ( .IN1(n18616), .IN2(n2783), .IN3(n18612), .IN4(n2748), .Q(
        n16027) );
  OA221X1 U24860 ( .IN1(n18621), .IN2(n2817), .IN3(n18617), .IN4(n14745), 
        .IN5(n16019), .Q(n16018) );
  OA22X1 U24861 ( .IN1(n18616), .IN2(n2782), .IN3(n18612), .IN4(n2747), .Q(
        n16019) );
  OA221X1 U24862 ( .IN1(n18621), .IN2(n2816), .IN3(n18617), .IN4(n14736), 
        .IN5(n16011), .Q(n16010) );
  OA22X1 U24863 ( .IN1(n18615), .IN2(n2781), .IN3(n18613), .IN4(n2746), .Q(
        n16011) );
  OA221X1 U24864 ( .IN1(n18621), .IN2(n2815), .IN3(n18619), .IN4(n14727), 
        .IN5(n16003), .Q(n16002) );
  OA22X1 U24865 ( .IN1(n18615), .IN2(n2780), .IN3(n18613), .IN4(n2745), .Q(
        n16003) );
  OA221X1 U24866 ( .IN1(n18621), .IN2(n2814), .IN3(n18617), .IN4(n14718), 
        .IN5(n15995), .Q(n15994) );
  OA22X1 U24867 ( .IN1(n18615), .IN2(n2779), .IN3(n18611), .IN4(n2744), .Q(
        n15995) );
  OA221X1 U24868 ( .IN1(n18621), .IN2(n2813), .IN3(n18617), .IN4(n14700), 
        .IN5(n15979), .Q(n15978) );
  OA22X1 U24869 ( .IN1(n18616), .IN2(n2778), .IN3(n18613), .IN4(n2743), .Q(
        n15979) );
  OA221X1 U24870 ( .IN1(n18622), .IN2(n2812), .IN3(n18617), .IN4(n14691), 
        .IN5(n15971), .Q(n15970) );
  OA22X1 U24871 ( .IN1(n18616), .IN2(n2777), .IN3(n18611), .IN4(n2742), .Q(
        n15971) );
  OA221X1 U24872 ( .IN1(n18621), .IN2(n2811), .IN3(n18618), .IN4(n14682), 
        .IN5(n15963), .Q(n15962) );
  OA22X1 U24873 ( .IN1(n18616), .IN2(n2776), .IN3(n18612), .IN4(n2741), .Q(
        n15963) );
  OA221X1 U24874 ( .IN1(n18620), .IN2(n2810), .IN3(n18617), .IN4(n14673), 
        .IN5(n15955), .Q(n15954) );
  OA22X1 U24875 ( .IN1(n18614), .IN2(n2775), .IN3(n18612), .IN4(n2740), .Q(
        n15955) );
  OA221X1 U24876 ( .IN1(n18622), .IN2(n2809), .IN3(n18617), .IN4(n14664), 
        .IN5(n15947), .Q(n15946) );
  OA22X1 U24877 ( .IN1(n18615), .IN2(n2774), .IN3(n18612), .IN4(n2739), .Q(
        n15947) );
  OA221X1 U24878 ( .IN1(n18622), .IN2(n2808), .IN3(n18618), .IN4(n14655), 
        .IN5(n15939), .Q(n15938) );
  OA22X1 U24879 ( .IN1(n18615), .IN2(n2773), .IN3(n18611), .IN4(n2738), .Q(
        n15939) );
  OA221X1 U24880 ( .IN1(n18620), .IN2(n2807), .IN3(n18619), .IN4(n14646), 
        .IN5(n15931), .Q(n15930) );
  OA22X1 U24881 ( .IN1(n18616), .IN2(n2772), .IN3(n18611), .IN4(n2737), .Q(
        n15931) );
  OA221X1 U24882 ( .IN1(n18620), .IN2(n2806), .IN3(n18618), .IN4(n14637), 
        .IN5(n15923), .Q(n15922) );
  OA22X1 U24883 ( .IN1(n18614), .IN2(n2771), .IN3(n18612), .IN4(n2736), .Q(
        n15923) );
  OA221X1 U24884 ( .IN1(n18620), .IN2(n2805), .IN3(n18619), .IN4(n14628), 
        .IN5(n15915), .Q(n15914) );
  OA22X1 U24885 ( .IN1(n18614), .IN2(n2770), .IN3(n18613), .IN4(n2735), .Q(
        n15915) );
  OA221X1 U24886 ( .IN1(n18621), .IN2(n2804), .IN3(n18617), .IN4(n14619), 
        .IN5(n15907), .Q(n15906) );
  OA22X1 U24887 ( .IN1(n18614), .IN2(n2769), .IN3(n18613), .IN4(n2734), .Q(
        n15907) );
  OA221X1 U24888 ( .IN1(n18621), .IN2(n2803), .IN3(n18617), .IN4(n14601), 
        .IN5(n15891), .Q(n15890) );
  OA22X1 U24889 ( .IN1(n18614), .IN2(n2768), .IN3(n18611), .IN4(n2733), .Q(
        n15891) );
  OA221X1 U24890 ( .IN1(n18620), .IN2(n2802), .IN3(n18617), .IN4(n14592), 
        .IN5(n15883), .Q(n15882) );
  OA22X1 U24891 ( .IN1(n18615), .IN2(n2767), .IN3(n18611), .IN4(n2732), .Q(
        n15883) );
  OA221X1 U24892 ( .IN1(n18572), .IN2(n2833), .IN3(n14808), .IN4(n18570), 
        .IN5(n16380), .Q(n16379) );
  OA22X1 U24893 ( .IN1(n18566), .IN2(n2798), .IN3(n18563), .IN4(n2763), .Q(
        n16380) );
  OA221X1 U24894 ( .IN1(n18574), .IN2(n2832), .IN3(n14709), .IN4(n18571), 
        .IN5(n16292), .Q(n16291) );
  OA22X1 U24895 ( .IN1(n18566), .IN2(n2797), .IN3(n18564), .IN4(n2762), .Q(
        n16292) );
  OA221X1 U24896 ( .IN1(n18572), .IN2(n2831), .IN3(n14610), .IN4(n18571), 
        .IN5(n16204), .Q(n16203) );
  OA22X1 U24897 ( .IN1(n18568), .IN2(n2796), .IN3(n18563), .IN4(n2761), .Q(
        n16204) );
  OA221X1 U24898 ( .IN1(n18572), .IN2(n2830), .IN3(n14583), .IN4(n18571), 
        .IN5(n16180), .Q(n16179) );
  OA22X1 U24899 ( .IN1(n18566), .IN2(n2795), .IN3(n16120), .IN4(n2760), .Q(
        n16180) );
  OA221X1 U24900 ( .IN1(n18574), .IN2(n2829), .IN3(n14574), .IN4(n18570), 
        .IN5(n16172), .Q(n16171) );
  OA22X1 U24901 ( .IN1(n18566), .IN2(n2794), .IN3(n16120), .IN4(n2759), .Q(
        n16172) );
  OA221X1 U24902 ( .IN1(n18573), .IN2(n2828), .IN3(n14565), .IN4(n18570), 
        .IN5(n16164), .Q(n16163) );
  OA22X1 U24903 ( .IN1(n18568), .IN2(n2793), .IN3(n16120), .IN4(n2758), .Q(
        n16164) );
  OA221X1 U24904 ( .IN1(n18574), .IN2(n2827), .IN3(n14556), .IN4(n18570), 
        .IN5(n16156), .Q(n16155) );
  OA22X1 U24905 ( .IN1(n18568), .IN2(n2792), .IN3(n18564), .IN4(n2757), .Q(
        n16156) );
  OA221X1 U24906 ( .IN1(n18574), .IN2(n2826), .IN3(n14547), .IN4(n18570), 
        .IN5(n16148), .Q(n16147) );
  OA22X1 U24907 ( .IN1(n18567), .IN2(n2791), .IN3(n18564), .IN4(n2756), .Q(
        n16148) );
  OA221X1 U24908 ( .IN1(n18574), .IN2(n2825), .IN3(n14538), .IN4(n18570), 
        .IN5(n16140), .Q(n16139) );
  OA22X1 U24909 ( .IN1(n18566), .IN2(n2790), .IN3(n18564), .IN4(n2755), .Q(
        n16140) );
  OA221X1 U24910 ( .IN1(n18574), .IN2(n2824), .IN3(n14514), .IN4(n18571), 
        .IN5(n16118), .Q(n16115) );
  OA22X1 U24911 ( .IN1(n18568), .IN2(n2789), .IN3(n18564), .IN4(n2754), .Q(
        n16118) );
  OA221X1 U24912 ( .IN1(n18572), .IN2(n2823), .IN3(n14799), .IN4(n18570), 
        .IN5(n16372), .Q(n16371) );
  OA22X1 U24913 ( .IN1(n18566), .IN2(n2788), .IN3(n18563), .IN4(n2753), .Q(
        n16372) );
  OA221X1 U24914 ( .IN1(n18572), .IN2(n2822), .IN3(n14790), .IN4(n18570), 
        .IN5(n16364), .Q(n16363) );
  OA22X1 U24915 ( .IN1(n18566), .IN2(n2787), .IN3(n18563), .IN4(n2752), .Q(
        n16364) );
  OA221X1 U24916 ( .IN1(n18572), .IN2(n2821), .IN3(n14781), .IN4(n18571), 
        .IN5(n16356), .Q(n16355) );
  OA22X1 U24917 ( .IN1(n18566), .IN2(n2786), .IN3(n18563), .IN4(n2751), .Q(
        n16356) );
  OA221X1 U24918 ( .IN1(n18573), .IN2(n2820), .IN3(n14772), .IN4(n18569), 
        .IN5(n16348), .Q(n16347) );
  OA22X1 U24919 ( .IN1(n18567), .IN2(n2785), .IN3(n16120), .IN4(n2750), .Q(
        n16348) );
  OA221X1 U24920 ( .IN1(n18573), .IN2(n2819), .IN3(n14763), .IN4(n18571), 
        .IN5(n16340), .Q(n16339) );
  OA22X1 U24921 ( .IN1(n18567), .IN2(n2784), .IN3(n16120), .IN4(n2749), .Q(
        n16340) );
  OA221X1 U24922 ( .IN1(n18573), .IN2(n2818), .IN3(n14754), .IN4(n18571), 
        .IN5(n16332), .Q(n16331) );
  OA22X1 U24923 ( .IN1(n18567), .IN2(n2783), .IN3(n16120), .IN4(n2748), .Q(
        n16332) );
  OA221X1 U24924 ( .IN1(n18573), .IN2(n2817), .IN3(n18569), .IN4(n14745), 
        .IN5(n16324), .Q(n16323) );
  OA22X1 U24925 ( .IN1(n18567), .IN2(n2782), .IN3(n18564), .IN4(n2747), .Q(
        n16324) );
  OA221X1 U24926 ( .IN1(n18573), .IN2(n2816), .IN3(n18569), .IN4(n14736), 
        .IN5(n16316), .Q(n16315) );
  OA22X1 U24927 ( .IN1(n18567), .IN2(n2781), .IN3(n18564), .IN4(n2746), .Q(
        n16316) );
  OA221X1 U24928 ( .IN1(n18573), .IN2(n2815), .IN3(n18571), .IN4(n14727), 
        .IN5(n16308), .Q(n16307) );
  OA22X1 U24929 ( .IN1(n18568), .IN2(n2780), .IN3(n16120), .IN4(n2745), .Q(
        n16308) );
  OA221X1 U24930 ( .IN1(n18574), .IN2(n2814), .IN3(n18569), .IN4(n14718), 
        .IN5(n16300), .Q(n16299) );
  OA22X1 U24931 ( .IN1(n18566), .IN2(n2779), .IN3(n18564), .IN4(n2744), .Q(
        n16300) );
  OA221X1 U24932 ( .IN1(n18572), .IN2(n2813), .IN3(n18569), .IN4(n14700), 
        .IN5(n16284), .Q(n16283) );
  OA22X1 U24933 ( .IN1(n18568), .IN2(n2778), .IN3(n16120), .IN4(n2743), .Q(
        n16284) );
  OA221X1 U24934 ( .IN1(n18573), .IN2(n2812), .IN3(n18569), .IN4(n14691), 
        .IN5(n16276), .Q(n16275) );
  OA22X1 U24935 ( .IN1(n18568), .IN2(n2777), .IN3(n16120), .IN4(n2742), .Q(
        n16276) );
  OA221X1 U24936 ( .IN1(n18572), .IN2(n2811), .IN3(n18570), .IN4(n14682), 
        .IN5(n16268), .Q(n16267) );
  OA22X1 U24937 ( .IN1(n18568), .IN2(n2776), .IN3(n18563), .IN4(n2741), .Q(
        n16268) );
  OA221X1 U24938 ( .IN1(n18574), .IN2(n2810), .IN3(n18569), .IN4(n14673), 
        .IN5(n16260), .Q(n16259) );
  OA22X1 U24939 ( .IN1(n18568), .IN2(n2775), .IN3(n16120), .IN4(n2740), .Q(
        n16260) );
  OA221X1 U24940 ( .IN1(n18574), .IN2(n2809), .IN3(n18569), .IN4(n14664), 
        .IN5(n16252), .Q(n16251) );
  OA22X1 U24941 ( .IN1(n18568), .IN2(n2774), .IN3(n18563), .IN4(n2739), .Q(
        n16252) );
  OA221X1 U24942 ( .IN1(n18574), .IN2(n2808), .IN3(n18570), .IN4(n14655), 
        .IN5(n16244), .Q(n16243) );
  OA22X1 U24943 ( .IN1(n18567), .IN2(n2773), .IN3(n18563), .IN4(n2738), .Q(
        n16244) );
  OA221X1 U24944 ( .IN1(n18572), .IN2(n2807), .IN3(n18571), .IN4(n14646), 
        .IN5(n16236), .Q(n16235) );
  OA22X1 U24945 ( .IN1(n18568), .IN2(n2772), .IN3(n16120), .IN4(n2737), .Q(
        n16236) );
  OA221X1 U24946 ( .IN1(n18572), .IN2(n2806), .IN3(n18570), .IN4(n14637), 
        .IN5(n16228), .Q(n16227) );
  OA22X1 U24947 ( .IN1(n18567), .IN2(n2771), .IN3(n18563), .IN4(n2736), .Q(
        n16228) );
  OA221X1 U24948 ( .IN1(n18573), .IN2(n2805), .IN3(n18571), .IN4(n14628), 
        .IN5(n16220), .Q(n16219) );
  OA22X1 U24949 ( .IN1(n18567), .IN2(n2770), .IN3(n16120), .IN4(n2735), .Q(
        n16220) );
  OA221X1 U24950 ( .IN1(n18572), .IN2(n2804), .IN3(n18569), .IN4(n14619), 
        .IN5(n16212), .Q(n16211) );
  OA22X1 U24951 ( .IN1(n18566), .IN2(n2769), .IN3(n18563), .IN4(n2734), .Q(
        n16212) );
  OA221X1 U24952 ( .IN1(n18574), .IN2(n2803), .IN3(n18569), .IN4(n14601), 
        .IN5(n16196), .Q(n16195) );
  OA22X1 U24953 ( .IN1(n18566), .IN2(n2768), .IN3(n18564), .IN4(n2733), .Q(
        n16196) );
  OA221X1 U24954 ( .IN1(n18573), .IN2(n2802), .IN3(n18569), .IN4(n14592), 
        .IN5(n16188), .Q(n16187) );
  OA22X1 U24955 ( .IN1(n18567), .IN2(n2767), .IN3(n18564), .IN4(n2732), .Q(
        n16188) );
  OA221X1 U24956 ( .IN1(n18524), .IN2(n2833), .IN3(n14808), .IN4(n18522), 
        .IN5(n16685), .Q(n16684) );
  OA22X1 U24957 ( .IN1(n18518), .IN2(n2798), .IN3(n18515), .IN4(n2763), .Q(
        n16685) );
  OA221X1 U24958 ( .IN1(n18525), .IN2(n2832), .IN3(n14709), .IN4(n18523), 
        .IN5(n16597), .Q(n16596) );
  OA22X1 U24959 ( .IN1(n18519), .IN2(n2797), .IN3(n18516), .IN4(n2762), .Q(
        n16597) );
  OA221X1 U24960 ( .IN1(n18525), .IN2(n2831), .IN3(n14610), .IN4(n18523), 
        .IN5(n16509), .Q(n16508) );
  OA22X1 U24961 ( .IN1(n18518), .IN2(n2796), .IN3(n18516), .IN4(n2761), .Q(
        n16509) );
  OA221X1 U24962 ( .IN1(n18526), .IN2(n2830), .IN3(n14583), .IN4(n18523), 
        .IN5(n16485), .Q(n16484) );
  OA22X1 U24963 ( .IN1(n18520), .IN2(n2795), .IN3(n18517), .IN4(n2760), .Q(
        n16485) );
  OA221X1 U24964 ( .IN1(n18524), .IN2(n2829), .IN3(n14574), .IN4(n18522), 
        .IN5(n16477), .Q(n16476) );
  OA22X1 U24965 ( .IN1(n18519), .IN2(n2794), .IN3(n18515), .IN4(n2759), .Q(
        n16477) );
  OA221X1 U24966 ( .IN1(n18526), .IN2(n2828), .IN3(n14565), .IN4(n18522), 
        .IN5(n16469), .Q(n16468) );
  OA22X1 U24967 ( .IN1(n18519), .IN2(n2793), .IN3(n18516), .IN4(n2758), .Q(
        n16469) );
  OA221X1 U24968 ( .IN1(n18526), .IN2(n2827), .IN3(n14556), .IN4(n18522), 
        .IN5(n16461), .Q(n16460) );
  OA22X1 U24969 ( .IN1(n18520), .IN2(n2792), .IN3(n18517), .IN4(n2757), .Q(
        n16461) );
  OA221X1 U24970 ( .IN1(n18526), .IN2(n2826), .IN3(n14547), .IN4(n18522), 
        .IN5(n16453), .Q(n16452) );
  OA22X1 U24971 ( .IN1(n18520), .IN2(n2791), .IN3(n18517), .IN4(n2756), .Q(
        n16453) );
  OA221X1 U24972 ( .IN1(n18526), .IN2(n2825), .IN3(n14538), .IN4(n18522), 
        .IN5(n16445), .Q(n16444) );
  OA22X1 U24973 ( .IN1(n18520), .IN2(n2790), .IN3(n18517), .IN4(n2755), .Q(
        n16445) );
  OA221X1 U24974 ( .IN1(n18526), .IN2(n2824), .IN3(n14514), .IN4(n18523), 
        .IN5(n16423), .Q(n16420) );
  OA22X1 U24975 ( .IN1(n18520), .IN2(n2789), .IN3(n18517), .IN4(n2754), .Q(
        n16423) );
  OA221X1 U24976 ( .IN1(n18524), .IN2(n2823), .IN3(n14799), .IN4(n18522), 
        .IN5(n16677), .Q(n16676) );
  OA22X1 U24977 ( .IN1(n18518), .IN2(n2788), .IN3(n18515), .IN4(n2753), .Q(
        n16677) );
  OA221X1 U24978 ( .IN1(n18524), .IN2(n2822), .IN3(n14790), .IN4(n18522), 
        .IN5(n16669), .Q(n16668) );
  OA22X1 U24979 ( .IN1(n18518), .IN2(n2787), .IN3(n18515), .IN4(n2752), .Q(
        n16669) );
  OA221X1 U24980 ( .IN1(n18524), .IN2(n2821), .IN3(n14781), .IN4(n18523), 
        .IN5(n16661), .Q(n16660) );
  OA22X1 U24981 ( .IN1(n18518), .IN2(n2786), .IN3(n18515), .IN4(n2751), .Q(
        n16661) );
  OA221X1 U24982 ( .IN1(n18524), .IN2(n2820), .IN3(n14772), .IN4(n18521), 
        .IN5(n16653), .Q(n16652) );
  OA22X1 U24983 ( .IN1(n18518), .IN2(n2785), .IN3(n18516), .IN4(n2750), .Q(
        n16653) );
  OA221X1 U24984 ( .IN1(n18525), .IN2(n2819), .IN3(n14763), .IN4(n18523), 
        .IN5(n16645), .Q(n16644) );
  OA22X1 U24985 ( .IN1(n18519), .IN2(n2784), .IN3(n18516), .IN4(n2749), .Q(
        n16645) );
  OA221X1 U24986 ( .IN1(n18526), .IN2(n2818), .IN3(n14754), .IN4(n18523), 
        .IN5(n16637), .Q(n16636) );
  OA22X1 U24987 ( .IN1(n18520), .IN2(n2783), .IN3(n18516), .IN4(n2748), .Q(
        n16637) );
  OA221X1 U24988 ( .IN1(n18525), .IN2(n2817), .IN3(n18521), .IN4(n14745), 
        .IN5(n16629), .Q(n16628) );
  OA22X1 U24989 ( .IN1(n18520), .IN2(n2782), .IN3(n18516), .IN4(n2747), .Q(
        n16629) );
  OA221X1 U24990 ( .IN1(n18525), .IN2(n2816), .IN3(n18521), .IN4(n14736), 
        .IN5(n16621), .Q(n16620) );
  OA22X1 U24991 ( .IN1(n18519), .IN2(n2781), .IN3(n18517), .IN4(n2746), .Q(
        n16621) );
  OA221X1 U24992 ( .IN1(n18525), .IN2(n2815), .IN3(n18523), .IN4(n14727), 
        .IN5(n16613), .Q(n16612) );
  OA22X1 U24993 ( .IN1(n18519), .IN2(n2780), .IN3(n18517), .IN4(n2745), .Q(
        n16613) );
  OA221X1 U24994 ( .IN1(n18525), .IN2(n2814), .IN3(n18521), .IN4(n14718), 
        .IN5(n16605), .Q(n16604) );
  OA22X1 U24995 ( .IN1(n18519), .IN2(n2779), .IN3(n18515), .IN4(n2744), .Q(
        n16605) );
  OA221X1 U24996 ( .IN1(n18525), .IN2(n2813), .IN3(n18521), .IN4(n14700), 
        .IN5(n16589), .Q(n16588) );
  OA22X1 U24997 ( .IN1(n18520), .IN2(n2778), .IN3(n18517), .IN4(n2743), .Q(
        n16589) );
  OA221X1 U24998 ( .IN1(n18526), .IN2(n2812), .IN3(n18521), .IN4(n14691), 
        .IN5(n16581), .Q(n16580) );
  OA22X1 U24999 ( .IN1(n18520), .IN2(n2777), .IN3(n18515), .IN4(n2742), .Q(
        n16581) );
  OA221X1 U25000 ( .IN1(n18525), .IN2(n2811), .IN3(n18522), .IN4(n14682), 
        .IN5(n16573), .Q(n16572) );
  OA22X1 U25001 ( .IN1(n18520), .IN2(n2776), .IN3(n18516), .IN4(n2741), .Q(
        n16573) );
  OA221X1 U25002 ( .IN1(n18524), .IN2(n2810), .IN3(n18521), .IN4(n14673), 
        .IN5(n16565), .Q(n16564) );
  OA22X1 U25003 ( .IN1(n18518), .IN2(n2775), .IN3(n18516), .IN4(n2740), .Q(
        n16565) );
  OA221X1 U25004 ( .IN1(n18526), .IN2(n2809), .IN3(n18521), .IN4(n14664), 
        .IN5(n16557), .Q(n16556) );
  OA22X1 U25005 ( .IN1(n18519), .IN2(n2774), .IN3(n18516), .IN4(n2739), .Q(
        n16557) );
  OA221X1 U25006 ( .IN1(n18526), .IN2(n2808), .IN3(n18522), .IN4(n14655), 
        .IN5(n16549), .Q(n16548) );
  OA22X1 U25007 ( .IN1(n18519), .IN2(n2773), .IN3(n18515), .IN4(n2738), .Q(
        n16549) );
  OA221X1 U25008 ( .IN1(n18524), .IN2(n2807), .IN3(n18523), .IN4(n14646), 
        .IN5(n16541), .Q(n16540) );
  OA22X1 U25009 ( .IN1(n18520), .IN2(n2772), .IN3(n18515), .IN4(n2737), .Q(
        n16541) );
  OA221X1 U25010 ( .IN1(n18524), .IN2(n2806), .IN3(n18522), .IN4(n14637), 
        .IN5(n16533), .Q(n16532) );
  OA22X1 U25011 ( .IN1(n18518), .IN2(n2771), .IN3(n18516), .IN4(n2736), .Q(
        n16533) );
  OA221X1 U25012 ( .IN1(n18524), .IN2(n2805), .IN3(n18523), .IN4(n14628), 
        .IN5(n16525), .Q(n16524) );
  OA22X1 U25013 ( .IN1(n18518), .IN2(n2770), .IN3(n18517), .IN4(n2735), .Q(
        n16525) );
  OA221X1 U25014 ( .IN1(n18525), .IN2(n2804), .IN3(n18521), .IN4(n14619), 
        .IN5(n16517), .Q(n16516) );
  OA22X1 U25015 ( .IN1(n18518), .IN2(n2769), .IN3(n18517), .IN4(n2734), .Q(
        n16517) );
  OA221X1 U25016 ( .IN1(n18525), .IN2(n2803), .IN3(n18521), .IN4(n14601), 
        .IN5(n16501), .Q(n16500) );
  OA22X1 U25017 ( .IN1(n18518), .IN2(n2768), .IN3(n18515), .IN4(n2733), .Q(
        n16501) );
  OA221X1 U25018 ( .IN1(n18524), .IN2(n2802), .IN3(n18521), .IN4(n14592), 
        .IN5(n16493), .Q(n16492) );
  OA22X1 U25019 ( .IN1(n18519), .IN2(n2767), .IN3(n18515), .IN4(n2732), .Q(
        n16493) );
  OA221X1 U25020 ( .IN1(n18476), .IN2(n2833), .IN3(n14808), .IN4(n18474), 
        .IN5(n16990), .Q(n16989) );
  OA22X1 U25021 ( .IN1(n18470), .IN2(n2798), .IN3(n18467), .IN4(n2763), .Q(
        n16990) );
  OA221X1 U25022 ( .IN1(n18478), .IN2(n2832), .IN3(n14709), .IN4(n18475), 
        .IN5(n16902), .Q(n16901) );
  OA22X1 U25023 ( .IN1(n18470), .IN2(n2797), .IN3(n18468), .IN4(n2762), .Q(
        n16902) );
  OA221X1 U25024 ( .IN1(n18476), .IN2(n2831), .IN3(n14610), .IN4(n18475), 
        .IN5(n16814), .Q(n16813) );
  OA22X1 U25025 ( .IN1(n18472), .IN2(n2796), .IN3(n18467), .IN4(n2761), .Q(
        n16814) );
  OA221X1 U25026 ( .IN1(n18476), .IN2(n2830), .IN3(n14583), .IN4(n18475), 
        .IN5(n16790), .Q(n16789) );
  OA22X1 U25027 ( .IN1(n18470), .IN2(n2795), .IN3(n16730), .IN4(n2760), .Q(
        n16790) );
  OA221X1 U25028 ( .IN1(n18478), .IN2(n2829), .IN3(n14574), .IN4(n18474), 
        .IN5(n16782), .Q(n16781) );
  OA22X1 U25029 ( .IN1(n18470), .IN2(n2794), .IN3(n16730), .IN4(n2759), .Q(
        n16782) );
  OA221X1 U25030 ( .IN1(n18477), .IN2(n2828), .IN3(n14565), .IN4(n18474), 
        .IN5(n16774), .Q(n16773) );
  OA22X1 U25031 ( .IN1(n18472), .IN2(n2793), .IN3(n16730), .IN4(n2758), .Q(
        n16774) );
  OA221X1 U25032 ( .IN1(n18478), .IN2(n2827), .IN3(n14556), .IN4(n18474), 
        .IN5(n16766), .Q(n16765) );
  OA22X1 U25033 ( .IN1(n18472), .IN2(n2792), .IN3(n18468), .IN4(n2757), .Q(
        n16766) );
  OA221X1 U25034 ( .IN1(n18478), .IN2(n2826), .IN3(n14547), .IN4(n18474), 
        .IN5(n16758), .Q(n16757) );
  OA22X1 U25035 ( .IN1(n18471), .IN2(n2791), .IN3(n18468), .IN4(n2756), .Q(
        n16758) );
  OA221X1 U25036 ( .IN1(n18478), .IN2(n2825), .IN3(n14538), .IN4(n18474), 
        .IN5(n16750), .Q(n16749) );
  OA22X1 U25037 ( .IN1(n18470), .IN2(n2790), .IN3(n18468), .IN4(n2755), .Q(
        n16750) );
  OA221X1 U25038 ( .IN1(n18478), .IN2(n2824), .IN3(n14514), .IN4(n18475), 
        .IN5(n16728), .Q(n16725) );
  OA22X1 U25039 ( .IN1(n18472), .IN2(n2789), .IN3(n18468), .IN4(n2754), .Q(
        n16728) );
  OA221X1 U25040 ( .IN1(n18476), .IN2(n2823), .IN3(n14799), .IN4(n18474), 
        .IN5(n16982), .Q(n16981) );
  OA22X1 U25041 ( .IN1(n18470), .IN2(n2788), .IN3(n18467), .IN4(n2753), .Q(
        n16982) );
  OA221X1 U25042 ( .IN1(n18476), .IN2(n2822), .IN3(n14790), .IN4(n18474), 
        .IN5(n16974), .Q(n16973) );
  OA22X1 U25043 ( .IN1(n18470), .IN2(n2787), .IN3(n18467), .IN4(n2752), .Q(
        n16974) );
  OA221X1 U25044 ( .IN1(n18476), .IN2(n2821), .IN3(n14781), .IN4(n18475), 
        .IN5(n16966), .Q(n16965) );
  OA22X1 U25045 ( .IN1(n18470), .IN2(n2786), .IN3(n18467), .IN4(n2751), .Q(
        n16966) );
  OA221X1 U25046 ( .IN1(n18477), .IN2(n2820), .IN3(n14772), .IN4(n18473), 
        .IN5(n16958), .Q(n16957) );
  OA22X1 U25047 ( .IN1(n18471), .IN2(n2785), .IN3(n16730), .IN4(n2750), .Q(
        n16958) );
  OA221X1 U25048 ( .IN1(n18477), .IN2(n2819), .IN3(n14763), .IN4(n18475), 
        .IN5(n16950), .Q(n16949) );
  OA22X1 U25049 ( .IN1(n18471), .IN2(n2784), .IN3(n16730), .IN4(n2749), .Q(
        n16950) );
  OA221X1 U25050 ( .IN1(n18477), .IN2(n2818), .IN3(n14754), .IN4(n18475), 
        .IN5(n16942), .Q(n16941) );
  OA22X1 U25051 ( .IN1(n18471), .IN2(n2783), .IN3(n16730), .IN4(n2748), .Q(
        n16942) );
  OA221X1 U25052 ( .IN1(n18477), .IN2(n2817), .IN3(n18473), .IN4(n14745), 
        .IN5(n16934), .Q(n16933) );
  OA22X1 U25053 ( .IN1(n18471), .IN2(n2782), .IN3(n18468), .IN4(n2747), .Q(
        n16934) );
  OA221X1 U25054 ( .IN1(n18477), .IN2(n2816), .IN3(n18473), .IN4(n14736), 
        .IN5(n16926), .Q(n16925) );
  OA22X1 U25055 ( .IN1(n18471), .IN2(n2781), .IN3(n18468), .IN4(n2746), .Q(
        n16926) );
  OA221X1 U25056 ( .IN1(n18477), .IN2(n2815), .IN3(n18475), .IN4(n14727), 
        .IN5(n16918), .Q(n16917) );
  OA22X1 U25057 ( .IN1(n18472), .IN2(n2780), .IN3(n16730), .IN4(n2745), .Q(
        n16918) );
  OA221X1 U25058 ( .IN1(n18478), .IN2(n2814), .IN3(n18473), .IN4(n14718), 
        .IN5(n16910), .Q(n16909) );
  OA22X1 U25059 ( .IN1(n18470), .IN2(n2779), .IN3(n18468), .IN4(n2744), .Q(
        n16910) );
  OA221X1 U25060 ( .IN1(n18476), .IN2(n2813), .IN3(n18473), .IN4(n14700), 
        .IN5(n16894), .Q(n16893) );
  OA22X1 U25061 ( .IN1(n18472), .IN2(n2778), .IN3(n16730), .IN4(n2743), .Q(
        n16894) );
  OA221X1 U25062 ( .IN1(n18477), .IN2(n2812), .IN3(n18473), .IN4(n14691), 
        .IN5(n16886), .Q(n16885) );
  OA22X1 U25063 ( .IN1(n18472), .IN2(n2777), .IN3(n16730), .IN4(n2742), .Q(
        n16886) );
  OA221X1 U25064 ( .IN1(n18476), .IN2(n2811), .IN3(n18474), .IN4(n14682), 
        .IN5(n16878), .Q(n16877) );
  OA22X1 U25065 ( .IN1(n18472), .IN2(n2776), .IN3(n18467), .IN4(n2741), .Q(
        n16878) );
  OA221X1 U25066 ( .IN1(n18478), .IN2(n2810), .IN3(n18473), .IN4(n14673), 
        .IN5(n16870), .Q(n16869) );
  OA22X1 U25067 ( .IN1(n18472), .IN2(n2775), .IN3(n16730), .IN4(n2740), .Q(
        n16870) );
  OA221X1 U25068 ( .IN1(n18478), .IN2(n2809), .IN3(n18473), .IN4(n14664), 
        .IN5(n16862), .Q(n16861) );
  OA22X1 U25069 ( .IN1(n18472), .IN2(n2774), .IN3(n18467), .IN4(n2739), .Q(
        n16862) );
  OA221X1 U25070 ( .IN1(n18478), .IN2(n2808), .IN3(n18474), .IN4(n14655), 
        .IN5(n16854), .Q(n16853) );
  OA22X1 U25071 ( .IN1(n18471), .IN2(n2773), .IN3(n18467), .IN4(n2738), .Q(
        n16854) );
  OA221X1 U25072 ( .IN1(n18476), .IN2(n2807), .IN3(n18475), .IN4(n14646), 
        .IN5(n16846), .Q(n16845) );
  OA22X1 U25073 ( .IN1(n18472), .IN2(n2772), .IN3(n16730), .IN4(n2737), .Q(
        n16846) );
  OA221X1 U25074 ( .IN1(n18476), .IN2(n2806), .IN3(n18474), .IN4(n14637), 
        .IN5(n16838), .Q(n16837) );
  OA22X1 U25075 ( .IN1(n18471), .IN2(n2771), .IN3(n18467), .IN4(n2736), .Q(
        n16838) );
  OA221X1 U25076 ( .IN1(n18477), .IN2(n2805), .IN3(n18475), .IN4(n14628), 
        .IN5(n16830), .Q(n16829) );
  OA22X1 U25077 ( .IN1(n18471), .IN2(n2770), .IN3(n16730), .IN4(n2735), .Q(
        n16830) );
  OA221X1 U25078 ( .IN1(n18476), .IN2(n2804), .IN3(n18473), .IN4(n14619), 
        .IN5(n16822), .Q(n16821) );
  OA22X1 U25079 ( .IN1(n18470), .IN2(n2769), .IN3(n18467), .IN4(n2734), .Q(
        n16822) );
  OA221X1 U25080 ( .IN1(n18478), .IN2(n2803), .IN3(n18473), .IN4(n14601), 
        .IN5(n16806), .Q(n16805) );
  OA22X1 U25081 ( .IN1(n18470), .IN2(n2768), .IN3(n18468), .IN4(n2733), .Q(
        n16806) );
  OA221X1 U25082 ( .IN1(n18477), .IN2(n2802), .IN3(n18473), .IN4(n14592), 
        .IN5(n16798), .Q(n16797) );
  OA22X1 U25083 ( .IN1(n18471), .IN2(n2767), .IN3(n18468), .IN4(n2732), .Q(
        n16798) );
  OA221X1 U25084 ( .IN1(n14496), .IN2(n14497), .IN3(n6887), .IN4(n2381), .IN5(
        n14498), .Q(n14491) );
  OA22X1 U25085 ( .IN1(n7367), .IN2(n2836), .IN3(n7663), .IN4(n2801), .Q(
        n14498) );
  OA221X1 U25086 ( .IN1(n14496), .IN2(n14506), .IN3(n6887), .IN4(n2380), .IN5(
        n14507), .Q(n14501) );
  OA22X1 U25087 ( .IN1(n7367), .IN2(n2835), .IN3(n7663), .IN4(n2800), .Q(
        n14507) );
  OA221X1 U25088 ( .IN1(n14851), .IN2(n14496), .IN3(n6887), .IN4(n2379), .IN5(
        n14852), .Q(n14814) );
  OA22X1 U25089 ( .IN1(n7367), .IN2(n2834), .IN3(n7663), .IN4(n2799), .Q(
        n14852) );
  OA221X1 U25090 ( .IN1(n14881), .IN2(n14497), .IN3(n6888), .IN4(n2381), .IN5(
        n14882), .Q(n14876) );
  OA22X1 U25091 ( .IN1(n7368), .IN2(n2836), .IN3(n7664), .IN4(n2801), .Q(
        n14882) );
  OA221X1 U25092 ( .IN1(n14881), .IN2(n14506), .IN3(n6888), .IN4(n2380), .IN5(
        n14890), .Q(n14885) );
  OA22X1 U25093 ( .IN1(n7368), .IN2(n2835), .IN3(n7664), .IN4(n2800), .Q(
        n14890) );
  OA221X1 U25094 ( .IN1(n14851), .IN2(n14881), .IN3(n6888), .IN4(n2379), .IN5(
        n15178), .Q(n15165) );
  OA22X1 U25095 ( .IN1(n7368), .IN2(n2834), .IN3(n7664), .IN4(n2799), .Q(
        n15178) );
  OA221X1 U25096 ( .IN1(n15186), .IN2(n14497), .IN3(n6889), .IN4(n2381), .IN5(
        n15187), .Q(n15181) );
  OA22X1 U25097 ( .IN1(n7369), .IN2(n2836), .IN3(n7665), .IN4(n2801), .Q(
        n15187) );
  OA221X1 U25098 ( .IN1(n15186), .IN2(n14506), .IN3(n6889), .IN4(n2380), .IN5(
        n15195), .Q(n15190) );
  OA22X1 U25099 ( .IN1(n7369), .IN2(n2835), .IN3(n7665), .IN4(n2800), .Q(
        n15195) );
  OA221X1 U25100 ( .IN1(n14851), .IN2(n15186), .IN3(n6889), .IN4(n2379), .IN5(
        n15483), .Q(n15470) );
  OA22X1 U25101 ( .IN1(n7369), .IN2(n2834), .IN3(n7665), .IN4(n2799), .Q(
        n15483) );
  OA221X1 U25102 ( .IN1(n15491), .IN2(n14497), .IN3(n6890), .IN4(n2381), .IN5(
        n15492), .Q(n15486) );
  OA22X1 U25103 ( .IN1(n7370), .IN2(n2836), .IN3(n7666), .IN4(n2801), .Q(
        n15492) );
  OA221X1 U25104 ( .IN1(n15491), .IN2(n14506), .IN3(n6890), .IN4(n2380), .IN5(
        n15500), .Q(n15495) );
  OA22X1 U25105 ( .IN1(n7370), .IN2(n2835), .IN3(n7666), .IN4(n2800), .Q(
        n15500) );
  OA221X1 U25106 ( .IN1(n14851), .IN2(n15491), .IN3(n6890), .IN4(n2379), .IN5(
        n15788), .Q(n15775) );
  OA22X1 U25107 ( .IN1(n7370), .IN2(n2834), .IN3(n7666), .IN4(n2799), .Q(
        n15788) );
  OA221X1 U25108 ( .IN1(n15796), .IN2(n14497), .IN3(n6891), .IN4(n2381), .IN5(
        n15797), .Q(n15791) );
  OA22X1 U25109 ( .IN1(n7371), .IN2(n2836), .IN3(n7667), .IN4(n2801), .Q(
        n15797) );
  OA221X1 U25110 ( .IN1(n15796), .IN2(n14506), .IN3(n6891), .IN4(n2380), .IN5(
        n15805), .Q(n15800) );
  OA22X1 U25111 ( .IN1(n7371), .IN2(n2835), .IN3(n7667), .IN4(n2800), .Q(
        n15805) );
  OA221X1 U25112 ( .IN1(n14851), .IN2(n15796), .IN3(n6891), .IN4(n2379), .IN5(
        n16093), .Q(n16080) );
  OA22X1 U25113 ( .IN1(n7371), .IN2(n2834), .IN3(n7667), .IN4(n2799), .Q(
        n16093) );
  OA221X1 U25114 ( .IN1(n16101), .IN2(n14497), .IN3(n6892), .IN4(n2381), .IN5(
        n16102), .Q(n16096) );
  OA22X1 U25115 ( .IN1(n7372), .IN2(n2836), .IN3(n7668), .IN4(n2801), .Q(
        n16102) );
  OA221X1 U25116 ( .IN1(n16101), .IN2(n14506), .IN3(n6892), .IN4(n2380), .IN5(
        n16110), .Q(n16105) );
  OA22X1 U25117 ( .IN1(n7372), .IN2(n2835), .IN3(n7668), .IN4(n2800), .Q(
        n16110) );
  OA221X1 U25118 ( .IN1(n14851), .IN2(n16101), .IN3(n6892), .IN4(n2379), .IN5(
        n16398), .Q(n16385) );
  OA22X1 U25119 ( .IN1(n7372), .IN2(n2834), .IN3(n7668), .IN4(n2799), .Q(
        n16398) );
  OA221X1 U25120 ( .IN1(n16406), .IN2(n14497), .IN3(n6893), .IN4(n2381), .IN5(
        n16407), .Q(n16401) );
  OA22X1 U25121 ( .IN1(n7373), .IN2(n2836), .IN3(n7669), .IN4(n2801), .Q(
        n16407) );
  OA221X1 U25122 ( .IN1(n16406), .IN2(n14506), .IN3(n6893), .IN4(n2380), .IN5(
        n16415), .Q(n16410) );
  OA22X1 U25123 ( .IN1(n7373), .IN2(n2835), .IN3(n7669), .IN4(n2800), .Q(
        n16415) );
  OA221X1 U25124 ( .IN1(n14851), .IN2(n16406), .IN3(n6893), .IN4(n2379), .IN5(
        n16703), .Q(n16690) );
  OA22X1 U25125 ( .IN1(n7373), .IN2(n2834), .IN3(n7669), .IN4(n2799), .Q(
        n16703) );
  OA221X1 U25126 ( .IN1(n16711), .IN2(n14497), .IN3(n6894), .IN4(n2381), .IN5(
        n16712), .Q(n16706) );
  OA22X1 U25127 ( .IN1(n7374), .IN2(n2836), .IN3(n7670), .IN4(n2801), .Q(
        n16712) );
  OA221X1 U25128 ( .IN1(n16711), .IN2(n14506), .IN3(n6894), .IN4(n2380), .IN5(
        n16720), .Q(n16715) );
  OA22X1 U25129 ( .IN1(n7374), .IN2(n2835), .IN3(n7670), .IN4(n2800), .Q(
        n16720) );
  OA221X1 U25130 ( .IN1(n14851), .IN2(n16711), .IN3(n6894), .IN4(n2379), .IN5(
        n17064), .Q(n16995) );
  OA22X1 U25131 ( .IN1(n7374), .IN2(n2834), .IN3(n7670), .IN4(n2799), .Q(
        n17064) );
  AO21X1 U25132 ( .IN1(n14046), .IN2(n14047), .IN3(n14044), .Q(n14004) );
  NAND3X0 U25133 ( .IN1(n14048), .IN2(n3254), .IN3(n14020), .QN(n14047) );
  OA22X1 U25134 ( .IN1(n18163), .IN2(n13863), .IN3(n13634), .IN4(n13844), .Q(
        n13866) );
  OA22X1 U25135 ( .IN1(n18164), .IN2(n13732), .IN3(n13670), .IN4(n13715), .Q(
        n13735) );
  OA22X1 U25136 ( .IN1(n18159), .IN2(n13554), .IN3(n13325), .IN4(n13535), .Q(
        n13557) );
  OA22X1 U25137 ( .IN1(n18165), .IN2(n13423), .IN3(n13361), .IN4(n13406), .Q(
        n13426) );
  OA22X1 U25138 ( .IN1(n18160), .IN2(n11388), .IN3(n11159), .IN4(n11369), .Q(
        n11391) );
  OA22X1 U25139 ( .IN1(n18166), .IN2(n11257), .IN3(n11195), .IN4(n11240), .Q(
        n11260) );
  OA22X1 U25140 ( .IN1(n18167), .IN2(n13245), .IN3(n13016), .IN4(n13226), .Q(
        n13248) );
  OA22X1 U25141 ( .IN1(n18168), .IN2(n13114), .IN3(n13052), .IN4(n13097), .Q(
        n13117) );
  OA22X1 U25142 ( .IN1(n18169), .IN2(n12936), .IN3(n12707), .IN4(n12917), .Q(
        n12939) );
  OA22X1 U25143 ( .IN1(n18170), .IN2(n12805), .IN3(n12743), .IN4(n12788), .Q(
        n12808) );
  OA22X1 U25144 ( .IN1(n18171), .IN2(n11079), .IN3(n10850), .IN4(n11060), .Q(
        n11082) );
  OA22X1 U25145 ( .IN1(n18172), .IN2(n10948), .IN3(n10886), .IN4(n10931), .Q(
        n10951) );
  OA22X1 U25146 ( .IN1(n18173), .IN2(n10769), .IN3(n10540), .IN4(n10750), .Q(
        n10772) );
  OA22X1 U25147 ( .IN1(n18174), .IN2(n10638), .IN3(n10576), .IN4(n10621), .Q(
        n10641) );
  OA22X1 U25148 ( .IN1(n18175), .IN2(n12627), .IN3(n12398), .IN4(n12608), .Q(
        n12630) );
  OA22X1 U25149 ( .IN1(n18176), .IN2(n12496), .IN3(n12434), .IN4(n12479), .Q(
        n12499) );
  OA22X1 U25150 ( .IN1(n18161), .IN2(n12318), .IN3(n12089), .IN4(n12299), .Q(
        n12321) );
  OA22X1 U25151 ( .IN1(n18177), .IN2(n12187), .IN3(n12125), .IN4(n12170), .Q(
        n12190) );
  OA22X1 U25152 ( .IN1(n18178), .IN2(n10460), .IN3(n10231), .IN4(n10441), .Q(
        n10463) );
  OA22X1 U25153 ( .IN1(n18179), .IN2(n10329), .IN3(n10267), .IN4(n10312), .Q(
        n10332) );
  OA22X1 U25154 ( .IN1(n18180), .IN2(n10150), .IN3(n9921), .IN4(n10131), .Q(
        n10153) );
  OA22X1 U25155 ( .IN1(n18181), .IN2(n10019), .IN3(n9957), .IN4(n10002), .Q(
        n10022) );
  OA22X1 U25156 ( .IN1(n18182), .IN2(n12008), .IN3(n11779), .IN4(n11989), .Q(
        n12011) );
  OA22X1 U25157 ( .IN1(n18183), .IN2(n11877), .IN3(n11815), .IN4(n11860), .Q(
        n11880) );
  OA22X1 U25158 ( .IN1(n18184), .IN2(n11698), .IN3(n11469), .IN4(n11679), .Q(
        n11701) );
  OA22X1 U25159 ( .IN1(n18185), .IN2(n11567), .IN3(n11505), .IN4(n11550), .Q(
        n11570) );
  OA22X1 U25160 ( .IN1(n18162), .IN2(n9840), .IN3(n9611), .IN4(n9821), .Q(
        n9843) );
  OA22X1 U25161 ( .IN1(n18186), .IN2(n9709), .IN3(n9647), .IN4(n9692), .Q(
        n9712) );
  OA22X1 U25162 ( .IN1(n18187), .IN2(n9529), .IN3(n9300), .IN4(n9510), .Q(
        n9532) );
  OA22X1 U25163 ( .IN1(n18188), .IN2(n9398), .IN3(n9336), .IN4(n9381), .Q(
        n9401) );
  AO21X1 U25164 ( .IN1(n13844), .IN2(n13845), .IN3(n18163), .Q(n13813) );
  NAND3X0 U25165 ( .IN1(n13634), .IN2(n3322), .IN3(n13814), .QN(n13845) );
  AO21X1 U25166 ( .IN1(n13715), .IN2(n13716), .IN3(n18164), .Q(n13688) );
  NAND3X0 U25167 ( .IN1(n13670), .IN2(n3318), .IN3(n13689), .QN(n13716) );
  AO21X1 U25168 ( .IN1(n13535), .IN2(n13536), .IN3(n18159), .Q(n13504) );
  NAND3X0 U25169 ( .IN1(n13325), .IN2(n3330), .IN3(n13505), .QN(n13536) );
  AO21X1 U25170 ( .IN1(n13406), .IN2(n13407), .IN3(n18165), .Q(n13379) );
  NAND3X0 U25171 ( .IN1(n13361), .IN2(n3326), .IN3(n13380), .QN(n13407) );
  AO21X1 U25172 ( .IN1(n11369), .IN2(n11370), .IN3(n18160), .Q(n11338) );
  NAND3X0 U25173 ( .IN1(n11159), .IN2(n3266), .IN3(n11339), .QN(n11370) );
  AO21X1 U25174 ( .IN1(n11240), .IN2(n11241), .IN3(n18166), .Q(n11213) );
  NAND3X0 U25175 ( .IN1(n11195), .IN2(n3262), .IN3(n11214), .QN(n11241) );
  AO21X1 U25176 ( .IN1(n13226), .IN2(n13227), .IN3(n18167), .Q(n13195) );
  NAND3X0 U25177 ( .IN1(n13016), .IN2(n3338), .IN3(n13196), .QN(n13227) );
  AO21X1 U25178 ( .IN1(n13097), .IN2(n13098), .IN3(n18168), .Q(n13070) );
  NAND3X0 U25179 ( .IN1(n13052), .IN2(n3334), .IN3(n13071), .QN(n13098) );
  AO21X1 U25180 ( .IN1(n12917), .IN2(n12918), .IN3(n18169), .Q(n12886) );
  NAND3X0 U25181 ( .IN1(n12707), .IN2(n3346), .IN3(n12887), .QN(n12918) );
  AO21X1 U25182 ( .IN1(n12788), .IN2(n12789), .IN3(n18170), .Q(n12761) );
  NAND3X0 U25183 ( .IN1(n12743), .IN2(n3342), .IN3(n12762), .QN(n12789) );
  AO21X1 U25184 ( .IN1(n11060), .IN2(n11061), .IN3(n18171), .Q(n11029) );
  NAND3X0 U25185 ( .IN1(n10850), .IN2(n3274), .IN3(n11030), .QN(n11061) );
  AO21X1 U25186 ( .IN1(n10931), .IN2(n10932), .IN3(n18172), .Q(n10904) );
  NAND3X0 U25187 ( .IN1(n10886), .IN2(n3270), .IN3(n10905), .QN(n10932) );
  AO21X1 U25188 ( .IN1(n10750), .IN2(n10751), .IN3(n18173), .Q(n10719) );
  NAND3X0 U25189 ( .IN1(n10540), .IN2(n3282), .IN3(n10720), .QN(n10751) );
  AO21X1 U25190 ( .IN1(n10621), .IN2(n10622), .IN3(n18174), .Q(n10594) );
  NAND3X0 U25191 ( .IN1(n10576), .IN2(n3278), .IN3(n10595), .QN(n10622) );
  AO21X1 U25192 ( .IN1(n12608), .IN2(n12609), .IN3(n18175), .Q(n12577) );
  NAND3X0 U25193 ( .IN1(n12398), .IN2(n3354), .IN3(n12578), .QN(n12609) );
  AO21X1 U25194 ( .IN1(n12479), .IN2(n12480), .IN3(n18176), .Q(n12452) );
  NAND3X0 U25195 ( .IN1(n12434), .IN2(n3350), .IN3(n12453), .QN(n12480) );
  AO21X1 U25196 ( .IN1(n12299), .IN2(n12300), .IN3(n18161), .Q(n12268) );
  NAND3X0 U25197 ( .IN1(n12089), .IN2(n3362), .IN3(n12269), .QN(n12300) );
  AO21X1 U25198 ( .IN1(n12170), .IN2(n12171), .IN3(n18177), .Q(n12143) );
  NAND3X0 U25199 ( .IN1(n12125), .IN2(n3358), .IN3(n12144), .QN(n12171) );
  AO21X1 U25200 ( .IN1(n10441), .IN2(n10442), .IN3(n18178), .Q(n10410) );
  NAND3X0 U25201 ( .IN1(n10231), .IN2(n3290), .IN3(n10411), .QN(n10442) );
  AO21X1 U25202 ( .IN1(n10312), .IN2(n10313), .IN3(n18179), .Q(n10285) );
  NAND3X0 U25203 ( .IN1(n10267), .IN2(n3286), .IN3(n10286), .QN(n10313) );
  AO21X1 U25204 ( .IN1(n10131), .IN2(n10132), .IN3(n18180), .Q(n10100) );
  NAND3X0 U25205 ( .IN1(n9921), .IN2(n3298), .IN3(n10101), .QN(n10132) );
  AO21X1 U25206 ( .IN1(n10002), .IN2(n10003), .IN3(n18181), .Q(n9975) );
  NAND3X0 U25207 ( .IN1(n9957), .IN2(n3294), .IN3(n9976), .QN(n10003) );
  AO21X1 U25208 ( .IN1(n11989), .IN2(n11990), .IN3(n18182), .Q(n11958) );
  NAND3X0 U25209 ( .IN1(n11779), .IN2(n3370), .IN3(n11959), .QN(n11990) );
  AO21X1 U25210 ( .IN1(n11860), .IN2(n11861), .IN3(n18183), .Q(n11833) );
  NAND3X0 U25211 ( .IN1(n11815), .IN2(n3366), .IN3(n11834), .QN(n11861) );
  AO21X1 U25212 ( .IN1(n11679), .IN2(n11680), .IN3(n18184), .Q(n11648) );
  NAND3X0 U25213 ( .IN1(n11469), .IN2(n3378), .IN3(n11649), .QN(n11680) );
  AO21X1 U25214 ( .IN1(n11550), .IN2(n11551), .IN3(n18185), .Q(n11523) );
  NAND3X0 U25215 ( .IN1(n11505), .IN2(n3374), .IN3(n11524), .QN(n11551) );
  AO21X1 U25216 ( .IN1(n9821), .IN2(n9822), .IN3(n18162), .Q(n9790) );
  NAND3X0 U25217 ( .IN1(n9611), .IN2(n3306), .IN3(n9791), .QN(n9822) );
  AO21X1 U25218 ( .IN1(n9692), .IN2(n9693), .IN3(n18186), .Q(n9665) );
  NAND3X0 U25219 ( .IN1(n9647), .IN2(n3302), .IN3(n9666), .QN(n9693) );
  AO21X1 U25220 ( .IN1(n9510), .IN2(n9511), .IN3(n18187), .Q(n9479) );
  NAND3X0 U25221 ( .IN1(n9300), .IN2(n3314), .IN3(n9480), .QN(n9511) );
  AO21X1 U25222 ( .IN1(n9381), .IN2(n9382), .IN3(n18188), .Q(n9354) );
  NAND3X0 U25223 ( .IN1(n9336), .IN2(n3310), .IN3(n9355), .QN(n9382) );
  OA21X1 U25224 ( .IN1(n14032), .IN2(n14039), .IN3(n14022), .Q(n14028) );
  OA21X1 U25225 ( .IN1(n13899), .IN2(n3433), .IN3(n13917), .Q(n13895) );
  OA21X1 U25226 ( .IN1(n13590), .IN2(n3437), .IN3(n13608), .Q(n13586) );
  OA21X1 U25227 ( .IN1(n11424), .IN2(n3405), .IN3(n11442), .Q(n11420) );
  OA21X1 U25228 ( .IN1(n13281), .IN2(n3441), .IN3(n13299), .Q(n13277) );
  OA21X1 U25229 ( .IN1(n12972), .IN2(n3445), .IN3(n12990), .Q(n12968) );
  OA21X1 U25230 ( .IN1(n11115), .IN2(n3409), .IN3(n11133), .Q(n11111) );
  OA21X1 U25231 ( .IN1(n10805), .IN2(n3413), .IN3(n10823), .Q(n10801) );
  OA21X1 U25232 ( .IN1(n12663), .IN2(n3449), .IN3(n12681), .Q(n12659) );
  OA21X1 U25233 ( .IN1(n12354), .IN2(n3453), .IN3(n12372), .Q(n12350) );
  OA21X1 U25234 ( .IN1(n10496), .IN2(n3417), .IN3(n10514), .Q(n10492) );
  OA21X1 U25235 ( .IN1(n10186), .IN2(n3421), .IN3(n10204), .Q(n10182) );
  OA21X1 U25236 ( .IN1(n12044), .IN2(n3457), .IN3(n12062), .Q(n12040) );
  OA21X1 U25237 ( .IN1(n11734), .IN2(n3461), .IN3(n11752), .Q(n11730) );
  OA21X1 U25238 ( .IN1(n9876), .IN2(n3425), .IN3(n9894), .Q(n9872) );
  OA21X1 U25239 ( .IN1(n9565), .IN2(n3429), .IN3(n9583), .Q(n9561) );
  OA21X1 U25240 ( .IN1(n13964), .IN2(n13971), .IN3(n13983), .Q(n13960) );
  OA21X1 U25241 ( .IN1(n14173), .IN2(n3399), .IN3(n14191), .Q(n14169) );
  OA21X1 U25242 ( .IN1(n14104), .IN2(n14111), .IN3(n14123), .Q(n14100) );
  AND2X1 U25243 ( .IN1(n13984), .IN2(n13985), .Q(n13964) );
  NAND3X0 U25244 ( .IN1(n18157), .IN2(n13944), .IN3(n4223), .QN(n13985) );
  AND2X1 U25245 ( .IN1(n14124), .IN2(n14125), .Q(n14104) );
  NAND3X0 U25246 ( .IN1(n18158), .IN2(n3382), .IN3(n4231), .QN(n14125) );
  ISOLANDX1 U25247 ( .D(n14132), .ISO(n14090), .Q(n14130) );
  ISOLANDX1 U25248 ( .D(n13992), .ISO(n13950), .Q(n13990) );
  AOI21X1 U25249 ( .IN1(n3865), .IN2(n18163), .IN3(n3862), .QN(n13851) );
  AOI21X1 U25250 ( .IN1(n3873), .IN2(n18164), .IN3(n3870), .QN(n13721) );
  AOI21X1 U25251 ( .IN1(n3820), .IN2(n18159), .IN3(n3817), .QN(n13542) );
  AOI21X1 U25252 ( .IN1(n3828), .IN2(n18165), .IN3(n3825), .QN(n13412) );
  AOI21X1 U25253 ( .IN1(n4180), .IN2(n18160), .IN3(n4177), .QN(n11376) );
  AOI21X1 U25254 ( .IN1(n4188), .IN2(n18166), .IN3(n4185), .QN(n11246) );
  AOI21X1 U25255 ( .IN1(n3775), .IN2(n18167), .IN3(n3772), .QN(n13233) );
  AOI21X1 U25256 ( .IN1(n3783), .IN2(n18168), .IN3(n3780), .QN(n13103) );
  AOI21X1 U25257 ( .IN1(n3730), .IN2(n18169), .IN3(n3727), .QN(n12924) );
  AOI21X1 U25258 ( .IN1(n3738), .IN2(n18170), .IN3(n3735), .QN(n12794) );
  AOI21X1 U25259 ( .IN1(n4135), .IN2(n18171), .IN3(n4132), .QN(n11067) );
  AOI21X1 U25260 ( .IN1(n4143), .IN2(n18172), .IN3(n4140), .QN(n10937) );
  AOI21X1 U25261 ( .IN1(n4090), .IN2(n18173), .IN3(n4087), .QN(n10757) );
  AOI21X1 U25262 ( .IN1(n4098), .IN2(n18174), .IN3(n4095), .QN(n10627) );
  AOI21X1 U25263 ( .IN1(n3685), .IN2(n18175), .IN3(n3682), .QN(n12615) );
  AOI21X1 U25264 ( .IN1(n3693), .IN2(n18176), .IN3(n3690), .QN(n12485) );
  AOI21X1 U25265 ( .IN1(n3640), .IN2(n18161), .IN3(n3637), .QN(n12306) );
  AOI21X1 U25266 ( .IN1(n3648), .IN2(n18177), .IN3(n3645), .QN(n12176) );
  AOI21X1 U25267 ( .IN1(n4045), .IN2(n18178), .IN3(n4042), .QN(n10448) );
  AOI21X1 U25268 ( .IN1(n4053), .IN2(n18179), .IN3(n4050), .QN(n10318) );
  AOI21X1 U25269 ( .IN1(n4000), .IN2(n18180), .IN3(n3997), .QN(n10138) );
  AOI21X1 U25270 ( .IN1(n4008), .IN2(n18181), .IN3(n4005), .QN(n10008) );
  AOI21X1 U25271 ( .IN1(n3595), .IN2(n18182), .IN3(n3592), .QN(n11996) );
  AOI21X1 U25272 ( .IN1(n3603), .IN2(n18183), .IN3(n3600), .QN(n11866) );
  AOI21X1 U25273 ( .IN1(n3550), .IN2(n18184), .IN3(n3547), .QN(n11686) );
  AOI21X1 U25274 ( .IN1(n3558), .IN2(n18185), .IN3(n3555), .QN(n11556) );
  AOI21X1 U25275 ( .IN1(n3955), .IN2(n18162), .IN3(n3952), .QN(n9828) );
  AOI21X1 U25276 ( .IN1(n3963), .IN2(n18186), .IN3(n3960), .QN(n9698) );
  AOI21X1 U25277 ( .IN1(n3910), .IN2(n18187), .IN3(n3907), .QN(n9517) );
  AOI21X1 U25278 ( .IN1(n3918), .IN2(n18188), .IN3(n3915), .QN(n9387) );
  AOI21X1 U25279 ( .IN1(n4225), .IN2(n18157), .IN3(n4222), .QN(n13984) );
  AOI21X1 U25280 ( .IN1(n4233), .IN2(n18158), .IN3(n4230), .QN(n14124) );
  OA21X1 U25281 ( .IN1(n13980), .IN2(n13981), .IN3(n13982), .Q(n13975) );
  OA21X1 U25282 ( .IN1(n13971), .IN2(n13963), .IN3(n13960), .Q(n13981) );
  OA21X1 U25283 ( .IN1(n14120), .IN2(n14121), .IN3(n14122), .Q(n14115) );
  OA21X1 U25284 ( .IN1(n14111), .IN2(n14103), .IN3(n14100), .Q(n14121) );
  NAND3X0 U25285 ( .IN1(n13814), .IN2(n13838), .IN3(n3321), .QN(n13806) );
  NAND3X0 U25286 ( .IN1(n13689), .IN2(n13677), .IN3(n3317), .QN(n13681) );
  NAND3X0 U25287 ( .IN1(n13505), .IN2(n13529), .IN3(n3329), .QN(n13497) );
  NAND3X0 U25288 ( .IN1(n13380), .IN2(n13368), .IN3(n3325), .QN(n13372) );
  NAND3X0 U25289 ( .IN1(n11339), .IN2(n11363), .IN3(n3265), .QN(n11331) );
  NAND3X0 U25290 ( .IN1(n11214), .IN2(n11202), .IN3(n3261), .QN(n11206) );
  NAND3X0 U25291 ( .IN1(n13196), .IN2(n13220), .IN3(n3337), .QN(n13188) );
  NAND3X0 U25292 ( .IN1(n13071), .IN2(n13059), .IN3(n3333), .QN(n13063) );
  NAND3X0 U25293 ( .IN1(n12887), .IN2(n12911), .IN3(n3345), .QN(n12879) );
  NAND3X0 U25294 ( .IN1(n12762), .IN2(n12750), .IN3(n3341), .QN(n12754) );
  NAND3X0 U25295 ( .IN1(n11030), .IN2(n11054), .IN3(n3273), .QN(n11022) );
  NAND3X0 U25296 ( .IN1(n10905), .IN2(n10893), .IN3(n3269), .QN(n10897) );
  NAND3X0 U25297 ( .IN1(n10720), .IN2(n10744), .IN3(n3281), .QN(n10712) );
  NAND3X0 U25298 ( .IN1(n10595), .IN2(n10583), .IN3(n3277), .QN(n10587) );
  NAND3X0 U25299 ( .IN1(n12578), .IN2(n12602), .IN3(n3353), .QN(n12570) );
  NAND3X0 U25300 ( .IN1(n12453), .IN2(n12441), .IN3(n3349), .QN(n12445) );
  NAND3X0 U25301 ( .IN1(n12269), .IN2(n12293), .IN3(n3361), .QN(n12261) );
  NAND3X0 U25302 ( .IN1(n12144), .IN2(n12132), .IN3(n3357), .QN(n12136) );
  NAND3X0 U25303 ( .IN1(n10411), .IN2(n10435), .IN3(n3289), .QN(n10403) );
  NAND3X0 U25304 ( .IN1(n10286), .IN2(n10274), .IN3(n3285), .QN(n10278) );
  NAND3X0 U25305 ( .IN1(n10101), .IN2(n10125), .IN3(n3297), .QN(n10093) );
  NAND3X0 U25306 ( .IN1(n9976), .IN2(n9964), .IN3(n3293), .QN(n9968) );
  NAND3X0 U25307 ( .IN1(n11959), .IN2(n11983), .IN3(n3369), .QN(n11951) );
  NAND3X0 U25308 ( .IN1(n11834), .IN2(n11822), .IN3(n3365), .QN(n11826) );
  NAND3X0 U25309 ( .IN1(n11649), .IN2(n11673), .IN3(n3377), .QN(n11641) );
  NAND3X0 U25310 ( .IN1(n11524), .IN2(n11512), .IN3(n3373), .QN(n11516) );
  NAND3X0 U25311 ( .IN1(n9791), .IN2(n9815), .IN3(n3305), .QN(n9783) );
  NAND3X0 U25312 ( .IN1(n9666), .IN2(n9654), .IN3(n3301), .QN(n9658) );
  NAND3X0 U25313 ( .IN1(n9480), .IN2(n9504), .IN3(n3313), .QN(n9472) );
  NAND3X0 U25314 ( .IN1(n9355), .IN2(n9343), .IN3(n3309), .QN(n9347) );
  AOI221X1 U25315 ( .IN1(n13919), .IN2(n3497), .IN3(n3323), .IN4(n13920), 
        .IN5(n13879), .QN(n13890) );
  AO221X1 U25316 ( .IN1(n13887), .IN2(n3882), .IN3(n2978), .IN4(n13894), .IN5(
        n13925), .Q(n13920) );
  ISOLANDX1 U25317 ( .D(n13918), .ISO(n3433), .Q(n13919) );
  INVX0 U25318 ( .IN(n13897), .QN(n2978) );
  AOI221X1 U25319 ( .IN1(n13610), .IN2(n3501), .IN3(n3331), .IN4(n13611), 
        .IN5(n13570), .QN(n13581) );
  AO221X1 U25320 ( .IN1(n13578), .IN2(n3837), .IN3(n2994), .IN4(n13585), .IN5(
        n13616), .Q(n13611) );
  ISOLANDX1 U25321 ( .D(n13609), .ISO(n3437), .Q(n13610) );
  INVX0 U25322 ( .IN(n13588), .QN(n2994) );
  AOI221X1 U25323 ( .IN1(n11444), .IN2(n3469), .IN3(n3267), .IN4(n11445), 
        .IN5(n11404), .QN(n11415) );
  AO221X1 U25324 ( .IN1(n11412), .IN2(n4197), .IN3(n2866), .IN4(n11419), .IN5(
        n11450), .Q(n11445) );
  ISOLANDX1 U25325 ( .D(n11443), .ISO(n3405), .Q(n11444) );
  INVX0 U25326 ( .IN(n11422), .QN(n2866) );
  AOI221X1 U25327 ( .IN1(n13301), .IN2(n3505), .IN3(n3339), .IN4(n13302), 
        .IN5(n13261), .QN(n13272) );
  AO221X1 U25328 ( .IN1(n13269), .IN2(n3792), .IN3(n3010), .IN4(n13276), .IN5(
        n13307), .Q(n13302) );
  ISOLANDX1 U25329 ( .D(n13300), .ISO(n3441), .Q(n13301) );
  INVX0 U25330 ( .IN(n13279), .QN(n3010) );
  AOI221X1 U25331 ( .IN1(n12992), .IN2(n3509), .IN3(n3347), .IN4(n12993), 
        .IN5(n12952), .QN(n12963) );
  AO221X1 U25332 ( .IN1(n12960), .IN2(n3747), .IN3(n3026), .IN4(n12967), .IN5(
        n12998), .Q(n12993) );
  ISOLANDX1 U25333 ( .D(n12991), .ISO(n3445), .Q(n12992) );
  INVX0 U25334 ( .IN(n12970), .QN(n3026) );
  AOI221X1 U25335 ( .IN1(n11135), .IN2(n3473), .IN3(n3275), .IN4(n11136), 
        .IN5(n11095), .QN(n11106) );
  AO221X1 U25336 ( .IN1(n11103), .IN2(n4152), .IN3(n2882), .IN4(n11110), .IN5(
        n11141), .Q(n11136) );
  ISOLANDX1 U25337 ( .D(n11134), .ISO(n3409), .Q(n11135) );
  INVX0 U25338 ( .IN(n11113), .QN(n2882) );
  AOI221X1 U25339 ( .IN1(n10825), .IN2(n3477), .IN3(n3283), .IN4(n10826), 
        .IN5(n10785), .QN(n10796) );
  AO221X1 U25340 ( .IN1(n10793), .IN2(n4107), .IN3(n2898), .IN4(n10800), .IN5(
        n10831), .Q(n10826) );
  ISOLANDX1 U25341 ( .D(n10824), .ISO(n3413), .Q(n10825) );
  INVX0 U25342 ( .IN(n10803), .QN(n2898) );
  AOI221X1 U25343 ( .IN1(n12683), .IN2(n3513), .IN3(n3355), .IN4(n12684), 
        .IN5(n12643), .QN(n12654) );
  AO221X1 U25344 ( .IN1(n12651), .IN2(n3702), .IN3(n3042), .IN4(n12658), .IN5(
        n12689), .Q(n12684) );
  ISOLANDX1 U25345 ( .D(n12682), .ISO(n3449), .Q(n12683) );
  INVX0 U25346 ( .IN(n12661), .QN(n3042) );
  AOI221X1 U25347 ( .IN1(n12374), .IN2(n3517), .IN3(n3363), .IN4(n12375), 
        .IN5(n12334), .QN(n12345) );
  AO221X1 U25348 ( .IN1(n12342), .IN2(n3657), .IN3(n3058), .IN4(n12349), .IN5(
        n12380), .Q(n12375) );
  ISOLANDX1 U25349 ( .D(n12373), .ISO(n3453), .Q(n12374) );
  INVX0 U25350 ( .IN(n12352), .QN(n3058) );
  AOI221X1 U25351 ( .IN1(n10516), .IN2(n3481), .IN3(n3291), .IN4(n10517), 
        .IN5(n10476), .QN(n10487) );
  AO221X1 U25352 ( .IN1(n10484), .IN2(n4062), .IN3(n2914), .IN4(n10491), .IN5(
        n10522), .Q(n10517) );
  ISOLANDX1 U25353 ( .D(n10515), .ISO(n3417), .Q(n10516) );
  INVX0 U25354 ( .IN(n10494), .QN(n2914) );
  AOI221X1 U25355 ( .IN1(n10206), .IN2(n3485), .IN3(n3299), .IN4(n10207), 
        .IN5(n10166), .QN(n10177) );
  AO221X1 U25356 ( .IN1(n10174), .IN2(n4017), .IN3(n2930), .IN4(n10181), .IN5(
        n10212), .Q(n10207) );
  ISOLANDX1 U25357 ( .D(n10205), .ISO(n3421), .Q(n10206) );
  INVX0 U25358 ( .IN(n10184), .QN(n2930) );
  AOI221X1 U25359 ( .IN1(n12064), .IN2(n3521), .IN3(n3371), .IN4(n12065), 
        .IN5(n12024), .QN(n12035) );
  AO221X1 U25360 ( .IN1(n12032), .IN2(n3612), .IN3(n3074), .IN4(n12039), .IN5(
        n12070), .Q(n12065) );
  ISOLANDX1 U25361 ( .D(n12063), .ISO(n3457), .Q(n12064) );
  INVX0 U25362 ( .IN(n12042), .QN(n3074) );
  AOI221X1 U25363 ( .IN1(n11754), .IN2(n3525), .IN3(n3379), .IN4(n11755), 
        .IN5(n11714), .QN(n11725) );
  AO221X1 U25364 ( .IN1(n11722), .IN2(n3567), .IN3(n3090), .IN4(n11729), .IN5(
        n11760), .Q(n11755) );
  ISOLANDX1 U25365 ( .D(n11753), .ISO(n3461), .Q(n11754) );
  INVX0 U25366 ( .IN(n11732), .QN(n3090) );
  AOI221X1 U25367 ( .IN1(n9896), .IN2(n3489), .IN3(n3307), .IN4(n9897), .IN5(
        n9856), .QN(n9867) );
  AO221X1 U25368 ( .IN1(n9864), .IN2(n3972), .IN3(n2946), .IN4(n9871), .IN5(
        n9902), .Q(n9897) );
  ISOLANDX1 U25369 ( .D(n9895), .ISO(n3425), .Q(n9896) );
  INVX0 U25370 ( .IN(n9874), .QN(n2946) );
  AOI221X1 U25371 ( .IN1(n9585), .IN2(n3493), .IN3(n3315), .IN4(n9586), .IN5(
        n9545), .QN(n9556) );
  AO221X1 U25372 ( .IN1(n9553), .IN2(n3927), .IN3(n2962), .IN4(n9560), .IN5(
        n9591), .Q(n9586) );
  ISOLANDX1 U25373 ( .D(n9584), .ISO(n3429), .Q(n9585) );
  INVX0 U25374 ( .IN(n9563), .QN(n2962) );
  AOI221X1 U25375 ( .IN1(n14193), .IN2(n3463), .IN3(n3255), .IN4(n14194), 
        .IN5(n14153), .QN(n14164) );
  AO221X1 U25376 ( .IN1(n14161), .IN2(n4242), .IN3(n2841), .IN4(n14168), .IN5(
        n14199), .Q(n14194) );
  ISOLANDX1 U25377 ( .D(n14192), .ISO(n3399), .Q(n14193) );
  INVX0 U25378 ( .IN(n14171), .QN(n2841) );
  AOI221X1 U25379 ( .IN1(n13986), .IN2(n13987), .IN3(n13950), .IN4(n13988), 
        .IN5(n13954), .QN(n13956) );
  NOR2X0 U25380 ( .IN1(n13971), .IN2(n13984), .QN(n13986) );
  AO221X1 U25381 ( .IN1(n13946), .IN2(n4226), .IN3(n2845), .IN4(n3191), .IN5(
        n13993), .Q(n13988) );
  INVX0 U25382 ( .IN(n13962), .QN(n2845) );
  AOI221X1 U25383 ( .IN1(n14126), .IN2(n14127), .IN3(n14090), .IN4(n14128), 
        .IN5(n14094), .QN(n14096) );
  NOR2X0 U25384 ( .IN1(n14111), .IN2(n14124), .QN(n14126) );
  AO221X1 U25385 ( .IN1(n14086), .IN2(n4234), .IN3(n2850), .IN4(n3192), .IN5(
        n14133), .Q(n14128) );
  INVX0 U25386 ( .IN(n14102), .QN(n2850) );
  AOI221X1 U25387 ( .IN1(n14054), .IN2(n14055), .IN3(n14018), .IN4(n14056), 
        .IN5(n14011), .QN(n14024) );
  ISOLANDX1 U25388 ( .D(n14053), .ISO(n14039), .Q(n14054) );
  AO221X1 U25389 ( .IN1(n14020), .IN2(n4218), .IN3(n2839), .IN4(n3189), .IN5(
        n14061), .Q(n14056) );
  INVX0 U25390 ( .IN(n14030), .QN(n2839) );
  NAND4X0 U25391 ( .IN1(n18163), .IN2(n13634), .IN3(n3496), .IN4(n3432), .QN(
        n13630) );
  NAND4X0 U25392 ( .IN1(n18159), .IN2(n13325), .IN3(n3500), .IN4(n3436), .QN(
        n13321) );
  NAND4X0 U25393 ( .IN1(n18160), .IN2(n11159), .IN3(n3468), .IN4(n3404), .QN(
        n11155) );
  NAND4X0 U25394 ( .IN1(n18167), .IN2(n13016), .IN3(n3504), .IN4(n3440), .QN(
        n13012) );
  NAND4X0 U25395 ( .IN1(n18169), .IN2(n12707), .IN3(n3508), .IN4(n3444), .QN(
        n12703) );
  NAND4X0 U25396 ( .IN1(n18171), .IN2(n10850), .IN3(n3472), .IN4(n3408), .QN(
        n10846) );
  NAND4X0 U25397 ( .IN1(n18173), .IN2(n10540), .IN3(n3476), .IN4(n3412), .QN(
        n10536) );
  NAND4X0 U25398 ( .IN1(n18175), .IN2(n12398), .IN3(n3512), .IN4(n3448), .QN(
        n12394) );
  NAND4X0 U25399 ( .IN1(n18161), .IN2(n12089), .IN3(n3516), .IN4(n3452), .QN(
        n12085) );
  NAND4X0 U25400 ( .IN1(n18178), .IN2(n10231), .IN3(n3480), .IN4(n3416), .QN(
        n10227) );
  NAND4X0 U25401 ( .IN1(n18180), .IN2(n9921), .IN3(n3484), .IN4(n3420), .QN(
        n9917) );
  NAND4X0 U25402 ( .IN1(n18182), .IN2(n11779), .IN3(n3520), .IN4(n3456), .QN(
        n11775) );
  NAND4X0 U25403 ( .IN1(n18184), .IN2(n11469), .IN3(n3524), .IN4(n3460), .QN(
        n11465) );
  NAND4X0 U25404 ( .IN1(n18162), .IN2(n9611), .IN3(n3488), .IN4(n3424), .QN(
        n9607) );
  NAND4X0 U25405 ( .IN1(n18187), .IN2(n9300), .IN3(n3492), .IN4(n3428), .QN(
        n9296) );
  NAND2X0 U25406 ( .IN1(n11296), .IN2(n11323), .QN(n11322) );
  NAND3X0 U25407 ( .IN1(n3403), .IN2(n11305), .IN3(n11281), .QN(n11323) );
  NAND2X0 U25408 ( .IN1(n10677), .IN2(n10704), .QN(n10703) );
  NAND3X0 U25409 ( .IN1(n3411), .IN2(n10686), .IN3(n10662), .QN(n10704) );
  NAND2X0 U25410 ( .IN1(n10058), .IN2(n10085), .QN(n10084) );
  NAND3X0 U25411 ( .IN1(n3419), .IN2(n10067), .IN3(n10043), .QN(n10085) );
  NAND2X0 U25412 ( .IN1(n9437), .IN2(n9464), .QN(n9463) );
  NAND3X0 U25413 ( .IN1(n3427), .IN2(n9446), .IN3(n9422), .QN(n9464) );
  NAND2X0 U25414 ( .IN1(n13771), .IN2(n13798), .QN(n13797) );
  NAND3X0 U25415 ( .IN1(n3431), .IN2(n13780), .IN3(n13756), .QN(n13798) );
  NAND2X0 U25416 ( .IN1(n13462), .IN2(n13489), .QN(n13488) );
  NAND3X0 U25417 ( .IN1(n3435), .IN2(n13471), .IN3(n13447), .QN(n13489) );
  NAND2X0 U25418 ( .IN1(n13153), .IN2(n13180), .QN(n13179) );
  NAND3X0 U25419 ( .IN1(n3439), .IN2(n13162), .IN3(n13138), .QN(n13180) );
  NAND2X0 U25420 ( .IN1(n12844), .IN2(n12871), .QN(n12870) );
  NAND3X0 U25421 ( .IN1(n3443), .IN2(n12853), .IN3(n12829), .QN(n12871) );
  NAND2X0 U25422 ( .IN1(n10987), .IN2(n11014), .QN(n11013) );
  NAND3X0 U25423 ( .IN1(n3407), .IN2(n10996), .IN3(n10972), .QN(n11014) );
  NAND2X0 U25424 ( .IN1(n12535), .IN2(n12562), .QN(n12561) );
  NAND3X0 U25425 ( .IN1(n3447), .IN2(n12544), .IN3(n12520), .QN(n12562) );
  NAND2X0 U25426 ( .IN1(n12226), .IN2(n12253), .QN(n12252) );
  NAND3X0 U25427 ( .IN1(n3451), .IN2(n12235), .IN3(n12211), .QN(n12253) );
  NAND2X0 U25428 ( .IN1(n10368), .IN2(n10395), .QN(n10394) );
  NAND3X0 U25429 ( .IN1(n3415), .IN2(n10377), .IN3(n10353), .QN(n10395) );
  NAND2X0 U25430 ( .IN1(n11916), .IN2(n11943), .QN(n11942) );
  NAND3X0 U25431 ( .IN1(n3455), .IN2(n11925), .IN3(n11901), .QN(n11943) );
  NAND2X0 U25432 ( .IN1(n11606), .IN2(n11633), .QN(n11632) );
  NAND3X0 U25433 ( .IN1(n3459), .IN2(n11615), .IN3(n11591), .QN(n11633) );
  NAND2X0 U25434 ( .IN1(n9748), .IN2(n9775), .QN(n9774) );
  NAND3X0 U25435 ( .IN1(n3423), .IN2(n9757), .IN3(n9733), .QN(n9775) );
  NAND2X0 U25436 ( .IN1(n14035), .IN2(n14062), .QN(n14061) );
  NAND3X0 U25437 ( .IN1(n3398), .IN2(n14044), .IN3(n14020), .QN(n14062) );
  AND3X1 U25438 ( .IN1(n2852), .IN2(s15_stb_o), .IN3(s15_addr_o[27]), .Q(
        n17086) );
  INVX0 U25439 ( .IN(n17764), .QN(n2852) );
  INVX0 U25440 ( .IN(n13913), .QN(n3390) );
  INVX0 U25441 ( .IN(n13604), .QN(n3391) );
  INVX0 U25442 ( .IN(n11438), .QN(n3383) );
  INVX0 U25443 ( .IN(n12677), .QN(n3394) );
  INVX0 U25444 ( .IN(n12368), .QN(n3395) );
  INVX0 U25445 ( .IN(n9890), .QN(n3388) );
  NAND4X0 U25446 ( .IN1(n13930), .IN2(n13931), .IN3(n13932), .IN4(n13933), 
        .QN(n13868) );
  OA22X1 U25447 ( .IN1(n13885), .IN2(n13888), .IN3(n13901), .IN4(n13894), .Q(
        n13931) );
  OA22X1 U25448 ( .IN1(n13907), .IN2(n13903), .IN3(n13902), .IN4(n13928), .Q(
        n13930) );
  OA22X1 U25449 ( .IN1(n13876), .IN2(n13927), .IN3(n13917), .IN4(n13883), .Q(
        n13933) );
  NAND4X0 U25450 ( .IN1(n13621), .IN2(n13622), .IN3(n13623), .IN4(n13624), 
        .QN(n13559) );
  OA22X1 U25451 ( .IN1(n13576), .IN2(n13579), .IN3(n13592), .IN4(n13585), .Q(
        n13622) );
  OA22X1 U25452 ( .IN1(n13598), .IN2(n13594), .IN3(n13593), .IN4(n13619), .Q(
        n13621) );
  OA22X1 U25453 ( .IN1(n13567), .IN2(n13618), .IN3(n13608), .IN4(n13574), .Q(
        n13624) );
  NAND4X0 U25454 ( .IN1(n11455), .IN2(n11456), .IN3(n11457), .IN4(n11458), 
        .QN(n11393) );
  OA22X1 U25455 ( .IN1(n11410), .IN2(n11413), .IN3(n11426), .IN4(n11419), .Q(
        n11456) );
  OA22X1 U25456 ( .IN1(n11432), .IN2(n11428), .IN3(n11427), .IN4(n11453), .Q(
        n11455) );
  OA22X1 U25457 ( .IN1(n11401), .IN2(n11452), .IN3(n11442), .IN4(n11408), .Q(
        n11458) );
  NAND4X0 U25458 ( .IN1(n13312), .IN2(n13313), .IN3(n13314), .IN4(n13315), 
        .QN(n13250) );
  OA22X1 U25459 ( .IN1(n13267), .IN2(n13270), .IN3(n13283), .IN4(n13276), .Q(
        n13313) );
  OA22X1 U25460 ( .IN1(n13289), .IN2(n13285), .IN3(n13284), .IN4(n13310), .Q(
        n13312) );
  OA22X1 U25461 ( .IN1(n13258), .IN2(n13309), .IN3(n13299), .IN4(n13265), .Q(
        n13315) );
  NAND4X0 U25462 ( .IN1(n13003), .IN2(n13004), .IN3(n13005), .IN4(n13006), 
        .QN(n12941) );
  OA22X1 U25463 ( .IN1(n12958), .IN2(n12961), .IN3(n12974), .IN4(n12967), .Q(
        n13004) );
  OA22X1 U25464 ( .IN1(n12980), .IN2(n12976), .IN3(n12975), .IN4(n13001), .Q(
        n13003) );
  OA22X1 U25465 ( .IN1(n12949), .IN2(n13000), .IN3(n12990), .IN4(n12956), .Q(
        n13006) );
  NAND4X0 U25466 ( .IN1(n11146), .IN2(n11147), .IN3(n11148), .IN4(n11149), 
        .QN(n11084) );
  OA22X1 U25467 ( .IN1(n11101), .IN2(n11104), .IN3(n11117), .IN4(n11110), .Q(
        n11147) );
  OA22X1 U25468 ( .IN1(n11123), .IN2(n11119), .IN3(n11118), .IN4(n11144), .Q(
        n11146) );
  OA22X1 U25469 ( .IN1(n11092), .IN2(n11143), .IN3(n11133), .IN4(n11099), .Q(
        n11149) );
  NAND4X0 U25470 ( .IN1(n10836), .IN2(n10837), .IN3(n10838), .IN4(n10839), 
        .QN(n10774) );
  OA22X1 U25471 ( .IN1(n10791), .IN2(n10794), .IN3(n10807), .IN4(n10800), .Q(
        n10837) );
  OA22X1 U25472 ( .IN1(n10813), .IN2(n10809), .IN3(n10808), .IN4(n10834), .Q(
        n10836) );
  OA22X1 U25473 ( .IN1(n10782), .IN2(n10833), .IN3(n10823), .IN4(n10789), .Q(
        n10839) );
  NAND4X0 U25474 ( .IN1(n12694), .IN2(n12695), .IN3(n12696), .IN4(n12697), 
        .QN(n12632) );
  OA22X1 U25475 ( .IN1(n12649), .IN2(n12652), .IN3(n12665), .IN4(n12658), .Q(
        n12695) );
  OA22X1 U25476 ( .IN1(n12671), .IN2(n12667), .IN3(n12666), .IN4(n12692), .Q(
        n12694) );
  OA22X1 U25477 ( .IN1(n12640), .IN2(n12691), .IN3(n12681), .IN4(n12647), .Q(
        n12697) );
  NAND4X0 U25478 ( .IN1(n12385), .IN2(n12386), .IN3(n12387), .IN4(n12388), 
        .QN(n12323) );
  OA22X1 U25479 ( .IN1(n12340), .IN2(n12343), .IN3(n12356), .IN4(n12349), .Q(
        n12386) );
  OA22X1 U25480 ( .IN1(n12362), .IN2(n12358), .IN3(n12357), .IN4(n12383), .Q(
        n12385) );
  OA22X1 U25481 ( .IN1(n12331), .IN2(n12382), .IN3(n12372), .IN4(n12338), .Q(
        n12388) );
  NAND4X0 U25482 ( .IN1(n10527), .IN2(n10528), .IN3(n10529), .IN4(n10530), 
        .QN(n10465) );
  OA22X1 U25483 ( .IN1(n10482), .IN2(n10485), .IN3(n10498), .IN4(n10491), .Q(
        n10528) );
  OA22X1 U25484 ( .IN1(n10504), .IN2(n10500), .IN3(n10499), .IN4(n10525), .Q(
        n10527) );
  OA22X1 U25485 ( .IN1(n10473), .IN2(n10524), .IN3(n10514), .IN4(n10480), .Q(
        n10530) );
  NAND4X0 U25486 ( .IN1(n10217), .IN2(n10218), .IN3(n10219), .IN4(n10220), 
        .QN(n10155) );
  OA22X1 U25487 ( .IN1(n10172), .IN2(n10175), .IN3(n10188), .IN4(n10181), .Q(
        n10218) );
  OA22X1 U25488 ( .IN1(n10194), .IN2(n10190), .IN3(n10189), .IN4(n10215), .Q(
        n10217) );
  OA22X1 U25489 ( .IN1(n10163), .IN2(n10214), .IN3(n10204), .IN4(n10170), .Q(
        n10220) );
  NAND4X0 U25490 ( .IN1(n12075), .IN2(n12076), .IN3(n12077), .IN4(n12078), 
        .QN(n12013) );
  OA22X1 U25491 ( .IN1(n12030), .IN2(n12033), .IN3(n12046), .IN4(n12039), .Q(
        n12076) );
  OA22X1 U25492 ( .IN1(n12052), .IN2(n12048), .IN3(n12047), .IN4(n12073), .Q(
        n12075) );
  OA22X1 U25493 ( .IN1(n12021), .IN2(n12072), .IN3(n12062), .IN4(n12028), .Q(
        n12078) );
  NAND4X0 U25494 ( .IN1(n11765), .IN2(n11766), .IN3(n11767), .IN4(n11768), 
        .QN(n11703) );
  OA22X1 U25495 ( .IN1(n11720), .IN2(n11723), .IN3(n11736), .IN4(n11729), .Q(
        n11766) );
  OA22X1 U25496 ( .IN1(n11742), .IN2(n11738), .IN3(n11737), .IN4(n11763), .Q(
        n11765) );
  OA22X1 U25497 ( .IN1(n11711), .IN2(n11762), .IN3(n11752), .IN4(n11718), .Q(
        n11768) );
  NAND4X0 U25498 ( .IN1(n9907), .IN2(n9908), .IN3(n9909), .IN4(n9910), .QN(
        n9845) );
  OA22X1 U25499 ( .IN1(n9862), .IN2(n9865), .IN3(n9878), .IN4(n9871), .Q(n9908) );
  OA22X1 U25500 ( .IN1(n9884), .IN2(n9880), .IN3(n9879), .IN4(n9905), .Q(n9907) );
  OA22X1 U25501 ( .IN1(n9853), .IN2(n9904), .IN3(n9894), .IN4(n9860), .Q(n9910) );
  NAND4X0 U25502 ( .IN1(n9596), .IN2(n9597), .IN3(n9598), .IN4(n9599), .QN(
        n9534) );
  OA22X1 U25503 ( .IN1(n9551), .IN2(n9554), .IN3(n9567), .IN4(n9560), .Q(n9597) );
  OA22X1 U25504 ( .IN1(n9573), .IN2(n9569), .IN3(n9568), .IN4(n9594), .Q(n9596) );
  OA22X1 U25505 ( .IN1(n9542), .IN2(n9593), .IN3(n9583), .IN4(n9549), .Q(n9599) );
  NAND4X0 U25506 ( .IN1(n13997), .IN2(n13998), .IN3(n13999), .IN4(n14000), 
        .QN(n13935) );
  OA22X1 U25507 ( .IN1(n3095), .IN2(n13970), .IN3(n13969), .IN4(n2844), .Q(
        n13997) );
  OA22X1 U25508 ( .IN1(n13948), .IN2(n3258), .IN3(n13967), .IN4(n3191), .Q(
        n13998) );
  OA22X1 U25509 ( .IN1(n3464), .IN2(n13995), .IN3(n13983), .IN4(n3400), .Q(
        n14000) );
  NAND4X0 U25510 ( .IN1(n14204), .IN2(n14205), .IN3(n14206), .IN4(n14207), 
        .QN(n14142) );
  OA22X1 U25511 ( .IN1(n14159), .IN2(n14162), .IN3(n14175), .IN4(n14168), .Q(
        n14205) );
  OA22X1 U25512 ( .IN1(n14181), .IN2(n14177), .IN3(n14176), .IN4(n14202), .Q(
        n14204) );
  OA22X1 U25513 ( .IN1(n14150), .IN2(n14201), .IN3(n14191), .IN4(n14157), .Q(
        n14207) );
  NAND4X0 U25514 ( .IN1(n14137), .IN2(n14138), .IN3(n14139), .IN4(n14140), 
        .QN(n14076) );
  OA22X1 U25515 ( .IN1(n3097), .IN2(n14110), .IN3(n14109), .IN4(n2849), .Q(
        n14137) );
  OA22X1 U25516 ( .IN1(n14088), .IN2(n3260), .IN3(n14107), .IN4(n3192), .Q(
        n14138) );
  OA22X1 U25517 ( .IN1(n3465), .IN2(n14135), .IN3(n14123), .IN4(n3401), .Q(
        n14140) );
  NAND4X0 U25518 ( .IN1(n3401), .IN2(n18158), .IN3(n14302), .IN4(n14303), .QN(
        n14272) );
  NOR2X0 U25519 ( .IN1(n14127), .IN2(n14120), .QN(n14302) );
  NOR4X0 U25520 ( .IN1(n14090), .IN2(n14141), .IN3(n14108), .IN4(n14105), .QN(
        n14303) );
  NOR2X0 U25521 ( .IN1(n18820), .IN2(n17764), .QN(s15_cyc_o) );
  AO21X1 U25522 ( .IN1(n13911), .IN2(n13912), .IN3(n13909), .Q(n13871) );
  NAND3X0 U25523 ( .IN1(n13913), .IN2(n13888), .IN3(n13887), .QN(n13912) );
  AO21X1 U25524 ( .IN1(n13602), .IN2(n13603), .IN3(n13600), .Q(n13562) );
  NAND3X0 U25525 ( .IN1(n13604), .IN2(n13579), .IN3(n13578), .QN(n13603) );
  AO21X1 U25526 ( .IN1(n11436), .IN2(n11437), .IN3(n11434), .Q(n11396) );
  NAND3X0 U25527 ( .IN1(n11438), .IN2(n11413), .IN3(n11412), .QN(n11437) );
  AO21X1 U25528 ( .IN1(n13293), .IN2(n13294), .IN3(n13291), .Q(n13253) );
  NAND3X0 U25529 ( .IN1(n13295), .IN2(n13270), .IN3(n13269), .QN(n13294) );
  AO21X1 U25530 ( .IN1(n12984), .IN2(n12985), .IN3(n12982), .Q(n12944) );
  NAND3X0 U25531 ( .IN1(n12986), .IN2(n12961), .IN3(n12960), .QN(n12985) );
  AO21X1 U25532 ( .IN1(n11127), .IN2(n11128), .IN3(n11125), .Q(n11087) );
  NAND3X0 U25533 ( .IN1(n11129), .IN2(n11104), .IN3(n11103), .QN(n11128) );
  AO21X1 U25534 ( .IN1(n10817), .IN2(n10818), .IN3(n10815), .Q(n10777) );
  NAND3X0 U25535 ( .IN1(n10819), .IN2(n10794), .IN3(n10793), .QN(n10818) );
  AO21X1 U25536 ( .IN1(n12675), .IN2(n12676), .IN3(n12673), .Q(n12635) );
  NAND3X0 U25537 ( .IN1(n12677), .IN2(n12652), .IN3(n12651), .QN(n12676) );
  AO21X1 U25538 ( .IN1(n12366), .IN2(n12367), .IN3(n12364), .Q(n12326) );
  NAND3X0 U25539 ( .IN1(n12368), .IN2(n12343), .IN3(n12342), .QN(n12367) );
  AO21X1 U25540 ( .IN1(n10508), .IN2(n10509), .IN3(n10506), .Q(n10468) );
  NAND3X0 U25541 ( .IN1(n10510), .IN2(n10485), .IN3(n10484), .QN(n10509) );
  AO21X1 U25542 ( .IN1(n10198), .IN2(n10199), .IN3(n10196), .Q(n10158) );
  NAND3X0 U25543 ( .IN1(n10200), .IN2(n10175), .IN3(n10174), .QN(n10199) );
  AO21X1 U25544 ( .IN1(n12056), .IN2(n12057), .IN3(n12054), .Q(n12016) );
  NAND3X0 U25545 ( .IN1(n12058), .IN2(n12033), .IN3(n12032), .QN(n12057) );
  AO21X1 U25546 ( .IN1(n11746), .IN2(n11747), .IN3(n11744), .Q(n11706) );
  NAND3X0 U25547 ( .IN1(n11748), .IN2(n11723), .IN3(n11722), .QN(n11747) );
  AO21X1 U25548 ( .IN1(n9888), .IN2(n9889), .IN3(n9886), .Q(n9848) );
  NAND3X0 U25549 ( .IN1(n9890), .IN2(n9865), .IN3(n9864), .QN(n9889) );
  AO21X1 U25550 ( .IN1(n9577), .IN2(n9578), .IN3(n9575), .Q(n9537) );
  NAND3X0 U25551 ( .IN1(n9579), .IN2(n9554), .IN3(n9553), .QN(n9578) );
  AO21X1 U25552 ( .IN1(n14185), .IN2(n14186), .IN3(n14183), .Q(n14145) );
  NAND3X0 U25553 ( .IN1(n14187), .IN2(n14162), .IN3(n14161), .QN(n14186) );
  OA22X1 U25554 ( .IN1(n13909), .IN2(n13929), .IN3(n13913), .IN4(n13911), .Q(
        n13932) );
  OA22X1 U25555 ( .IN1(n13600), .IN2(n13620), .IN3(n13604), .IN4(n13602), .Q(
        n13623) );
  OA22X1 U25556 ( .IN1(n11434), .IN2(n11454), .IN3(n11438), .IN4(n11436), .Q(
        n11457) );
  OA22X1 U25557 ( .IN1(n13291), .IN2(n13311), .IN3(n13295), .IN4(n13293), .Q(
        n13314) );
  OA22X1 U25558 ( .IN1(n12982), .IN2(n13002), .IN3(n12986), .IN4(n12984), .Q(
        n13005) );
  OA22X1 U25559 ( .IN1(n11125), .IN2(n11145), .IN3(n11129), .IN4(n11127), .Q(
        n11148) );
  OA22X1 U25560 ( .IN1(n10815), .IN2(n10835), .IN3(n10819), .IN4(n10817), .Q(
        n10838) );
  OA22X1 U25561 ( .IN1(n12673), .IN2(n12693), .IN3(n12677), .IN4(n12675), .Q(
        n12696) );
  OA22X1 U25562 ( .IN1(n12364), .IN2(n12384), .IN3(n12368), .IN4(n12366), .Q(
        n12387) );
  OA22X1 U25563 ( .IN1(n10506), .IN2(n10526), .IN3(n10510), .IN4(n10508), .Q(
        n10529) );
  OA22X1 U25564 ( .IN1(n10196), .IN2(n10216), .IN3(n10200), .IN4(n10198), .Q(
        n10219) );
  OA22X1 U25565 ( .IN1(n12054), .IN2(n12074), .IN3(n12058), .IN4(n12056), .Q(
        n12077) );
  OA22X1 U25566 ( .IN1(n11744), .IN2(n11764), .IN3(n11748), .IN4(n11746), .Q(
        n11767) );
  OA22X1 U25567 ( .IN1(n9886), .IN2(n9906), .IN3(n9890), .IN4(n9888), .Q(n9909) );
  OA22X1 U25568 ( .IN1(n9575), .IN2(n9595), .IN3(n9579), .IN4(n9577), .Q(n9598) );
  OA22X1 U25569 ( .IN1(n14183), .IN2(n14203), .IN3(n14187), .IN4(n14185), .Q(
        n14206) );
  OA22X1 U25570 ( .IN1(n18157), .IN2(n13996), .IN3(n13944), .IN4(n13977), .Q(
        n13999) );
  AO21X1 U25571 ( .IN1(n13977), .IN2(n13978), .IN3(n18157), .Q(n13945) );
  NAND3X0 U25572 ( .IN1(n13944), .IN2(n3258), .IN3(n13946), .QN(n13978) );
  AO21X1 U25573 ( .IN1(n14117), .IN2(n14118), .IN3(n18158), .Q(n14085) );
  NAND3X0 U25574 ( .IN1(n3382), .IN2(n3260), .IN3(n14086), .QN(n14118) );
  NAND4X0 U25575 ( .IN1(n18333), .IN2(n13666), .IN3(n13667), .IN4(n18247), 
        .QN(n13653) );
  NAND4X0 U25576 ( .IN1(n18332), .IN2(n13357), .IN3(n13358), .IN4(n13359), 
        .QN(n13344) );
  NAND4X0 U25577 ( .IN1(n18331), .IN2(n11191), .IN3(n11192), .IN4(n11193), 
        .QN(n11178) );
  NAND4X0 U25578 ( .IN1(n18330), .IN2(n18278), .IN3(n13049), .IN4(n18256), 
        .QN(n13035) );
  NAND4X0 U25579 ( .IN1(n18329), .IN2(n18274), .IN3(n12740), .IN4(n18252), 
        .QN(n12726) );
  NAND4X0 U25580 ( .IN1(n18328), .IN2(n18277), .IN3(n10883), .IN4(n18255), 
        .QN(n10869) );
  NAND4X0 U25581 ( .IN1(n18327), .IN2(n18264), .IN3(n10573), .IN4(n18251), 
        .QN(n10559) );
  NAND4X0 U25582 ( .IN1(n18326), .IN2(n12430), .IN3(n12431), .IN4(n18248), 
        .QN(n12417) );
  NAND4X0 U25583 ( .IN1(n18325), .IN2(n12121), .IN3(n12122), .IN4(n12123), 
        .QN(n12108) );
  NAND4X0 U25584 ( .IN1(n18324), .IN2(n18276), .IN3(n10264), .IN4(n18254), 
        .QN(n10250) );
  NAND4X0 U25585 ( .IN1(n18323), .IN2(n18263), .IN3(n9954), .IN4(n18250), .QN(
        n9940) );
  NAND4X0 U25586 ( .IN1(n18322), .IN2(n18275), .IN3(n11812), .IN4(n18253), 
        .QN(n11798) );
  NAND4X0 U25587 ( .IN1(n18321), .IN2(n18262), .IN3(n11502), .IN4(n18249), 
        .QN(n11488) );
  NAND4X0 U25588 ( .IN1(n18320), .IN2(n9643), .IN3(n9644), .IN4(n9645), .QN(
        n9630) );
  NAND4X0 U25589 ( .IN1(n18319), .IN2(n18279), .IN3(n9333), .IN4(n18257), .QN(
        n9319) );
  NAND2X0 U25590 ( .IN1(n13901), .IN2(n13926), .QN(n13925) );
  NAND3X0 U25591 ( .IN1(n13883), .IN2(n13909), .IN3(n13887), .QN(n13926) );
  NAND2X0 U25592 ( .IN1(n13592), .IN2(n13617), .QN(n13616) );
  NAND3X0 U25593 ( .IN1(n13574), .IN2(n13600), .IN3(n13578), .QN(n13617) );
  NAND2X0 U25594 ( .IN1(n11426), .IN2(n11451), .QN(n11450) );
  NAND3X0 U25595 ( .IN1(n11408), .IN2(n11434), .IN3(n11412), .QN(n11451) );
  NAND2X0 U25596 ( .IN1(n13283), .IN2(n13308), .QN(n13307) );
  NAND3X0 U25597 ( .IN1(n13265), .IN2(n13291), .IN3(n13269), .QN(n13308) );
  NAND2X0 U25598 ( .IN1(n12974), .IN2(n12999), .QN(n12998) );
  NAND3X0 U25599 ( .IN1(n12956), .IN2(n12982), .IN3(n12960), .QN(n12999) );
  NAND2X0 U25600 ( .IN1(n11117), .IN2(n11142), .QN(n11141) );
  NAND3X0 U25601 ( .IN1(n11099), .IN2(n11125), .IN3(n11103), .QN(n11142) );
  NAND2X0 U25602 ( .IN1(n10807), .IN2(n10832), .QN(n10831) );
  NAND3X0 U25603 ( .IN1(n10789), .IN2(n10815), .IN3(n10793), .QN(n10832) );
  NAND2X0 U25604 ( .IN1(n12665), .IN2(n12690), .QN(n12689) );
  NAND3X0 U25605 ( .IN1(n12647), .IN2(n12673), .IN3(n12651), .QN(n12690) );
  NAND2X0 U25606 ( .IN1(n12356), .IN2(n12381), .QN(n12380) );
  NAND3X0 U25607 ( .IN1(n12338), .IN2(n12364), .IN3(n12342), .QN(n12381) );
  NAND2X0 U25608 ( .IN1(n10498), .IN2(n10523), .QN(n10522) );
  NAND3X0 U25609 ( .IN1(n10480), .IN2(n10506), .IN3(n10484), .QN(n10523) );
  NAND2X0 U25610 ( .IN1(n10188), .IN2(n10213), .QN(n10212) );
  NAND3X0 U25611 ( .IN1(n10170), .IN2(n10196), .IN3(n10174), .QN(n10213) );
  NAND2X0 U25612 ( .IN1(n12046), .IN2(n12071), .QN(n12070) );
  NAND3X0 U25613 ( .IN1(n12028), .IN2(n12054), .IN3(n12032), .QN(n12071) );
  NAND2X0 U25614 ( .IN1(n11736), .IN2(n11761), .QN(n11760) );
  NAND3X0 U25615 ( .IN1(n11718), .IN2(n11744), .IN3(n11722), .QN(n11761) );
  NAND2X0 U25616 ( .IN1(n9878), .IN2(n9903), .QN(n9902) );
  NAND3X0 U25617 ( .IN1(n9860), .IN2(n9886), .IN3(n9864), .QN(n9903) );
  NAND2X0 U25618 ( .IN1(n9567), .IN2(n9592), .QN(n9591) );
  NAND3X0 U25619 ( .IN1(n9549), .IN2(n9575), .IN3(n9553), .QN(n9592) );
  NAND2X0 U25620 ( .IN1(n14175), .IN2(n14200), .QN(n14199) );
  NAND3X0 U25621 ( .IN1(n14157), .IN2(n14183), .IN3(n14161), .QN(n14200) );
  NAND3X0 U25622 ( .IN1(n13887), .IN2(n13883), .IN3(n3324), .QN(n13874) );
  NAND3X0 U25623 ( .IN1(n13578), .IN2(n13574), .IN3(n3332), .QN(n13565) );
  NAND3X0 U25624 ( .IN1(n11412), .IN2(n11408), .IN3(n3268), .QN(n11399) );
  NAND3X0 U25625 ( .IN1(n13269), .IN2(n13265), .IN3(n3340), .QN(n13256) );
  NAND3X0 U25626 ( .IN1(n12960), .IN2(n12956), .IN3(n3348), .QN(n12947) );
  NAND3X0 U25627 ( .IN1(n11103), .IN2(n11099), .IN3(n3276), .QN(n11090) );
  NAND3X0 U25628 ( .IN1(n10793), .IN2(n10789), .IN3(n3284), .QN(n10780) );
  NAND3X0 U25629 ( .IN1(n12651), .IN2(n12647), .IN3(n3356), .QN(n12638) );
  NAND3X0 U25630 ( .IN1(n12342), .IN2(n12338), .IN3(n3364), .QN(n12329) );
  NAND3X0 U25631 ( .IN1(n10484), .IN2(n10480), .IN3(n3292), .QN(n10471) );
  NAND3X0 U25632 ( .IN1(n10174), .IN2(n10170), .IN3(n3300), .QN(n10161) );
  NAND3X0 U25633 ( .IN1(n12032), .IN2(n12028), .IN3(n3372), .QN(n12019) );
  NAND3X0 U25634 ( .IN1(n11722), .IN2(n11718), .IN3(n3380), .QN(n11709) );
  NAND3X0 U25635 ( .IN1(n9864), .IN2(n9860), .IN3(n3308), .QN(n9851) );
  NAND3X0 U25636 ( .IN1(n9553), .IN2(n9549), .IN3(n3316), .QN(n9540) );
  NAND3X0 U25637 ( .IN1(n14161), .IN2(n14157), .IN3(n3256), .QN(n14148) );
  OA21X1 U25638 ( .IN1(n13943), .IN2(n13944), .IN3(n13945), .Q(n13942) );
  AOI21X1 U25639 ( .IN1(n3258), .IN2(n13946), .IN3(n2846), .QN(n13943) );
  OA22X1 U25640 ( .IN1(n18158), .IN2(n14136), .IN3(n3382), .IN4(n14117), .Q(
        n14139) );
  NAND3X0 U25641 ( .IN1(n13971), .IN2(n13946), .IN3(n3257), .QN(n13937) );
  NAND3X0 U25642 ( .IN1(n14111), .IN2(n14086), .IN3(n3259), .QN(n14078) );
  NOR2X0 U25643 ( .IN1(n9283), .IN2(n18816), .QN(rf_N115) );
  AND4X1 U25644 ( .IN1(n9284), .IN2(n9285), .IN3(n9286), .IN4(n9287), .Q(n9283) );
  OA221X1 U25645 ( .IN1(n18390), .IN2(n18144), .IN3(n18386), .IN4(n18022), 
        .IN5(n9291), .Q(n9284) );
  OA221X1 U25646 ( .IN1(n18374), .IN2(n18142), .IN3(n18370), .IN4(n18021), 
        .IN5(n9290), .Q(n9285) );
  NOR2X0 U25647 ( .IN1(n9274), .IN2(n18816), .QN(rf_N116) );
  AND4X1 U25648 ( .IN1(n9275), .IN2(n9276), .IN3(n9277), .IN4(n9278), .Q(n9274) );
  OA221X1 U25649 ( .IN1(n18390), .IN2(n17991), .IN3(n18386), .IN4(n18100), 
        .IN5(n9282), .Q(n9275) );
  OA221X1 U25650 ( .IN1(n18374), .IN2(n17989), .IN3(n18370), .IN4(n18099), 
        .IN5(n9281), .Q(n9276) );
  NOR2X0 U25651 ( .IN1(n9265), .IN2(n18816), .QN(rf_N117) );
  AND4X1 U25652 ( .IN1(n9266), .IN2(n9267), .IN3(n9268), .IN4(n9269), .Q(n9265) );
  OA221X1 U25653 ( .IN1(n18390), .IN2(n18110), .IN3(n18386), .IN4(n17970), 
        .IN5(n9273), .Q(n9266) );
  OA221X1 U25654 ( .IN1(n18374), .IN2(n18106), .IN3(n18370), .IN4(n17968), 
        .IN5(n9272), .Q(n9267) );
  NOR2X0 U25655 ( .IN1(n9256), .IN2(n18816), .QN(rf_N118) );
  AND4X1 U25656 ( .IN1(n9257), .IN2(n9258), .IN3(n9259), .IN4(n9260), .Q(n9256) );
  OA221X1 U25657 ( .IN1(n18390), .IN2(n17987), .IN3(n18386), .IN4(n18096), 
        .IN5(n9264), .Q(n9257) );
  OA221X1 U25658 ( .IN1(n18374), .IN2(n17985), .IN3(n18370), .IN4(n18095), 
        .IN5(n9263), .Q(n9258) );
  NOR2X0 U25659 ( .IN1(n9247), .IN2(n18816), .QN(rf_N119) );
  AND4X1 U25660 ( .IN1(n9248), .IN2(n9249), .IN3(n9250), .IN4(n9251), .Q(n9247) );
  OA221X1 U25661 ( .IN1(n18390), .IN2(n18111), .IN3(n18386), .IN4(n17971), 
        .IN5(n9255), .Q(n9248) );
  OA221X1 U25662 ( .IN1(n18374), .IN2(n18107), .IN3(n18370), .IN4(n17969), 
        .IN5(n9254), .Q(n9249) );
  NOR2X0 U25663 ( .IN1(n9238), .IN2(n18816), .QN(rf_N120) );
  AND4X1 U25664 ( .IN1(n9239), .IN2(n9240), .IN3(n9241), .IN4(n9242), .Q(n9238) );
  OA221X1 U25665 ( .IN1(n18390), .IN2(n17981), .IN3(n18386), .IN4(n18091), 
        .IN5(n9246), .Q(n9239) );
  OA221X1 U25666 ( .IN1(n18374), .IN2(n17977), .IN3(n18370), .IN4(n18089), 
        .IN5(n9245), .Q(n9240) );
  NOR2X0 U25667 ( .IN1(n9229), .IN2(n18816), .QN(rf_N121) );
  AND4X1 U25668 ( .IN1(n9230), .IN2(n9231), .IN3(n9232), .IN4(n9233), .Q(n9229) );
  OA221X1 U25669 ( .IN1(n18391), .IN2(n18104), .IN3(n18387), .IN4(n17966), 
        .IN5(n9237), .Q(n9230) );
  OA221X1 U25670 ( .IN1(n18375), .IN2(n18102), .IN3(n18371), .IN4(n17965), 
        .IN5(n9236), .Q(n9231) );
  NOR2X0 U25671 ( .IN1(n9220), .IN2(n18815), .QN(rf_N122) );
  AND4X1 U25672 ( .IN1(n9221), .IN2(n9222), .IN3(n9223), .IN4(n9224), .Q(n9220) );
  OA221X1 U25673 ( .IN1(n18391), .IN2(n17982), .IN3(n18387), .IN4(n18092), 
        .IN5(n9228), .Q(n9221) );
  OA221X1 U25674 ( .IN1(n18375), .IN2(n17978), .IN3(n18371), .IN4(n18090), 
        .IN5(n9227), .Q(n9222) );
  NOR2X0 U25675 ( .IN1(n9211), .IN2(n18815), .QN(rf_N123) );
  AND4X1 U25676 ( .IN1(n9212), .IN2(n9213), .IN3(n9214), .IN4(n9215), .Q(n9211) );
  OA221X1 U25677 ( .IN1(n18391), .IN2(n17946), .IN3(n18387), .IN4(n18151), 
        .IN5(n9219), .Q(n9212) );
  OA221X1 U25678 ( .IN1(n18375), .IN2(n17947), .IN3(n18371), .IN4(n18152), 
        .IN5(n9218), .Q(n9213) );
  NOR2X0 U25679 ( .IN1(n9202), .IN2(n18815), .QN(rf_N124) );
  AND4X1 U25680 ( .IN1(n9203), .IN2(n9204), .IN3(n9205), .IN4(n9206), .Q(n9202) );
  OA221X1 U25681 ( .IN1(n18391), .IN2(n18154), .IN3(n18387), .IN4(n17945), 
        .IN5(n9210), .Q(n9203) );
  OA221X1 U25682 ( .IN1(n18375), .IN2(n18155), .IN3(n18371), .IN4(n17964), 
        .IN5(n9209), .Q(n9204) );
  NOR2X0 U25683 ( .IN1(n9193), .IN2(n18815), .QN(rf_N125) );
  AND4X1 U25684 ( .IN1(n9194), .IN2(n9195), .IN3(n9196), .IN4(n9197), .Q(n9193) );
  OA221X1 U25685 ( .IN1(n18391), .IN2(n17943), .IN3(n18387), .IN4(n18067), 
        .IN5(n9201), .Q(n9194) );
  OA221X1 U25686 ( .IN1(n18375), .IN2(n17941), .IN3(n18371), .IN4(n18069), 
        .IN5(n9200), .Q(n9195) );
  NOR2X0 U25687 ( .IN1(n9184), .IN2(n18816), .QN(rf_N126) );
  AND4X1 U25688 ( .IN1(n9185), .IN2(n9186), .IN3(n9187), .IN4(n9188), .Q(n9184) );
  OA221X1 U25689 ( .IN1(n18391), .IN2(n18077), .IN3(n18387), .IN4(n17951), 
        .IN5(n9192), .Q(n9185) );
  OA221X1 U25690 ( .IN1(n18375), .IN2(n18075), .IN3(n18371), .IN4(n17950), 
        .IN5(n9191), .Q(n9186) );
  NOR2X0 U25691 ( .IN1(n9175), .IN2(n18817), .QN(rf_N127) );
  AND4X1 U25692 ( .IN1(n9176), .IN2(n9177), .IN3(n9178), .IN4(n9179), .Q(n9175) );
  OA221X1 U25693 ( .IN1(n18391), .IN2(n18199), .IN3(n18387), .IN4(n18030), 
        .IN5(n9183), .Q(n9176) );
  OA221X1 U25694 ( .IN1(n18375), .IN2(n18197), .IN3(n18371), .IN4(n18029), 
        .IN5(n9182), .Q(n9177) );
  NOR2X0 U25695 ( .IN1(n9166), .IN2(n18819), .QN(rf_N128) );
  AND4X1 U25696 ( .IN1(n9167), .IN2(n9168), .IN3(n9169), .IN4(n9170), .Q(n9166) );
  OA221X1 U25697 ( .IN1(n18391), .IN2(n18043), .IN3(n18387), .IN4(n18195), 
        .IN5(n9174), .Q(n9167) );
  OA221X1 U25698 ( .IN1(n18375), .IN2(n18041), .IN3(n18371), .IN4(n18194), 
        .IN5(n9173), .Q(n9168) );
  NOR2X0 U25699 ( .IN1(n9157), .IN2(n18815), .QN(rf_N129) );
  AND4X1 U25700 ( .IN1(n9158), .IN2(n9159), .IN3(n9160), .IN4(n9161), .Q(n9157) );
  OA221X1 U25701 ( .IN1(n18391), .IN2(n18203), .IN3(n18387), .IN4(n18033), 
        .IN5(n9165), .Q(n9158) );
  OA221X1 U25702 ( .IN1(n18375), .IN2(n18201), .IN3(n18371), .IN4(n18032), 
        .IN5(n9164), .Q(n9159) );
  NOR2X0 U25703 ( .IN1(n9132), .IN2(n18818), .QN(rf_N130) );
  AND4X1 U25704 ( .IN1(n9133), .IN2(n9134), .IN3(n9135), .IN4(n9136), .Q(n9132) );
  OA221X1 U25705 ( .IN1(n18391), .IN2(n18039), .IN3(n18387), .IN4(n18192), 
        .IN5(n9154), .Q(n9133) );
  OA221X1 U25706 ( .IN1(n18375), .IN2(n18037), .IN3(n18371), .IN4(n18191), 
        .IN5(n9149), .Q(n9134) );
  NAND4X0 U25707 ( .IN1(n3400), .IN2(n18157), .IN3(n2844), .IN4(n3464), .QN(
        n14273) );
  INVX0 U25708 ( .IN(n17765), .QN(s14_cyc_o) );
  INVX0 U25709 ( .IN(n17766), .QN(s13_cyc_o) );
  INVX0 U25710 ( .IN(n17767), .QN(s12_cyc_o) );
  INVX0 U25711 ( .IN(n17768), .QN(s11_cyc_o) );
  INVX0 U25712 ( .IN(n17769), .QN(s10_cyc_o) );
  INVX0 U25713 ( .IN(n17770), .QN(s9_cyc_o) );
  INVX0 U25714 ( .IN(n17771), .QN(s8_cyc_o) );
  INVX0 U25715 ( .IN(n17772), .QN(s7_cyc_o) );
  INVX0 U25716 ( .IN(n17773), .QN(s6_cyc_o) );
  INVX0 U25717 ( .IN(n17774), .QN(s5_cyc_o) );
  INVX0 U25718 ( .IN(n17775), .QN(s4_cyc_o) );
  INVX0 U25719 ( .IN(n17776), .QN(s3_cyc_o) );
  INVX0 U25720 ( .IN(n17777), .QN(s2_cyc_o) );
  INVX0 U25721 ( .IN(n17778), .QN(s1_cyc_o) );
  INVX0 U25722 ( .IN(n17779), .QN(s0_cyc_o) );
  NAND2X0 U25723 ( .IN1(n13967), .IN2(n13994), .QN(n13993) );
  NAND3X0 U25724 ( .IN1(n3400), .IN2(n18157), .IN3(n13946), .QN(n13994) );
  NAND2X0 U25725 ( .IN1(n14107), .IN2(n14134), .QN(n14133) );
  NAND3X0 U25726 ( .IN1(n3401), .IN2(n18158), .IN3(n14086), .QN(n14134) );
  NAND2X0 U25727 ( .IN1(n13834), .IN2(n13861), .QN(n13860) );
  NAND3X0 U25728 ( .IN1(n3432), .IN2(n18163), .IN3(n13814), .QN(n13861) );
  NAND2X0 U25729 ( .IN1(n13707), .IN2(n13730), .QN(n13729) );
  NAND3X0 U25730 ( .IN1(n3430), .IN2(n18164), .IN3(n13689), .QN(n13730) );
  NAND2X0 U25731 ( .IN1(n13525), .IN2(n13552), .QN(n13551) );
  NAND3X0 U25732 ( .IN1(n3436), .IN2(n18159), .IN3(n13505), .QN(n13552) );
  NAND2X0 U25733 ( .IN1(n13398), .IN2(n13421), .QN(n13420) );
  NAND3X0 U25734 ( .IN1(n3434), .IN2(n18165), .IN3(n13380), .QN(n13421) );
  NAND2X0 U25735 ( .IN1(n11359), .IN2(n11386), .QN(n11385) );
  NAND3X0 U25736 ( .IN1(n3404), .IN2(n18160), .IN3(n11339), .QN(n11386) );
  NAND2X0 U25737 ( .IN1(n11232), .IN2(n11255), .QN(n11254) );
  NAND3X0 U25738 ( .IN1(n3402), .IN2(n18166), .IN3(n11214), .QN(n11255) );
  NAND2X0 U25739 ( .IN1(n13216), .IN2(n13243), .QN(n13242) );
  NAND3X0 U25740 ( .IN1(n3440), .IN2(n18167), .IN3(n13196), .QN(n13243) );
  NAND2X0 U25741 ( .IN1(n13089), .IN2(n13112), .QN(n13111) );
  NAND3X0 U25742 ( .IN1(n3438), .IN2(n18168), .IN3(n13071), .QN(n13112) );
  NAND2X0 U25743 ( .IN1(n12907), .IN2(n12934), .QN(n12933) );
  NAND3X0 U25744 ( .IN1(n3444), .IN2(n18169), .IN3(n12887), .QN(n12934) );
  NAND2X0 U25745 ( .IN1(n12780), .IN2(n12803), .QN(n12802) );
  NAND3X0 U25746 ( .IN1(n3442), .IN2(n18170), .IN3(n12762), .QN(n12803) );
  NAND2X0 U25747 ( .IN1(n11050), .IN2(n11077), .QN(n11076) );
  NAND3X0 U25748 ( .IN1(n3408), .IN2(n18171), .IN3(n11030), .QN(n11077) );
  NAND2X0 U25749 ( .IN1(n10923), .IN2(n10946), .QN(n10945) );
  NAND3X0 U25750 ( .IN1(n3406), .IN2(n18172), .IN3(n10905), .QN(n10946) );
  NAND2X0 U25751 ( .IN1(n10740), .IN2(n10767), .QN(n10766) );
  NAND3X0 U25752 ( .IN1(n3412), .IN2(n18173), .IN3(n10720), .QN(n10767) );
  NAND2X0 U25753 ( .IN1(n10613), .IN2(n10636), .QN(n10635) );
  NAND3X0 U25754 ( .IN1(n3410), .IN2(n18174), .IN3(n10595), .QN(n10636) );
  NAND2X0 U25755 ( .IN1(n12598), .IN2(n12625), .QN(n12624) );
  NAND3X0 U25756 ( .IN1(n3448), .IN2(n18175), .IN3(n12578), .QN(n12625) );
  NAND2X0 U25757 ( .IN1(n12471), .IN2(n12494), .QN(n12493) );
  NAND3X0 U25758 ( .IN1(n3446), .IN2(n18176), .IN3(n12453), .QN(n12494) );
  NAND2X0 U25759 ( .IN1(n12289), .IN2(n12316), .QN(n12315) );
  NAND3X0 U25760 ( .IN1(n3452), .IN2(n18161), .IN3(n12269), .QN(n12316) );
  NAND2X0 U25761 ( .IN1(n12162), .IN2(n12185), .QN(n12184) );
  NAND3X0 U25762 ( .IN1(n3450), .IN2(n18177), .IN3(n12144), .QN(n12185) );
  NAND2X0 U25763 ( .IN1(n10431), .IN2(n10458), .QN(n10457) );
  NAND3X0 U25764 ( .IN1(n3416), .IN2(n18178), .IN3(n10411), .QN(n10458) );
  NAND2X0 U25765 ( .IN1(n10304), .IN2(n10327), .QN(n10326) );
  NAND3X0 U25766 ( .IN1(n3414), .IN2(n18179), .IN3(n10286), .QN(n10327) );
  NAND2X0 U25767 ( .IN1(n10121), .IN2(n10148), .QN(n10147) );
  NAND3X0 U25768 ( .IN1(n3420), .IN2(n18180), .IN3(n10101), .QN(n10148) );
  NAND2X0 U25769 ( .IN1(n9994), .IN2(n10017), .QN(n10016) );
  NAND3X0 U25770 ( .IN1(n3418), .IN2(n18181), .IN3(n9976), .QN(n10017) );
  NAND2X0 U25771 ( .IN1(n11979), .IN2(n12006), .QN(n12005) );
  NAND3X0 U25772 ( .IN1(n3456), .IN2(n18182), .IN3(n11959), .QN(n12006) );
  NAND2X0 U25773 ( .IN1(n11852), .IN2(n11875), .QN(n11874) );
  NAND3X0 U25774 ( .IN1(n3454), .IN2(n18183), .IN3(n11834), .QN(n11875) );
  NAND2X0 U25775 ( .IN1(n11669), .IN2(n11696), .QN(n11695) );
  NAND3X0 U25776 ( .IN1(n3460), .IN2(n18184), .IN3(n11649), .QN(n11696) );
  NAND2X0 U25777 ( .IN1(n11542), .IN2(n11565), .QN(n11564) );
  NAND3X0 U25778 ( .IN1(n3458), .IN2(n18185), .IN3(n11524), .QN(n11565) );
  NAND2X0 U25779 ( .IN1(n9811), .IN2(n9838), .QN(n9837) );
  NAND3X0 U25780 ( .IN1(n3424), .IN2(n18162), .IN3(n9791), .QN(n9838) );
  NAND2X0 U25781 ( .IN1(n9684), .IN2(n9707), .QN(n9706) );
  NAND3X0 U25782 ( .IN1(n3422), .IN2(n18186), .IN3(n9666), .QN(n9707) );
  NAND2X0 U25783 ( .IN1(n9500), .IN2(n9527), .QN(n9526) );
  NAND3X0 U25784 ( .IN1(n3428), .IN2(n18187), .IN3(n9480), .QN(n9527) );
  NAND2X0 U25785 ( .IN1(n9373), .IN2(n9396), .QN(n9395) );
  NAND3X0 U25786 ( .IN1(n3426), .IN2(n18188), .IN3(n9355), .QN(n9396) );
  AO22X1 U25787 ( .IN1(n14330), .IN2(n18321), .IN3(n14331), .IN4(n18625), .Q(
        n17684) );
  AO22X1 U25788 ( .IN1(n14330), .IN2(n18322), .IN3(n14331), .IN4(n17860), .Q(
        n17685) );
  AO22X1 U25789 ( .IN1(n14330), .IN2(n18325), .IN3(n14331), .IN4(n17837), .Q(
        n17686) );
  AO22X1 U25790 ( .IN1(n14330), .IN2(n18326), .IN3(n14331), .IN4(n18631), .Q(
        n17687) );
  AO22X1 U25791 ( .IN1(n14330), .IN2(n18329), .IN3(n14331), .IN4(n17839), .Q(
        n17688) );
  AO22X1 U25792 ( .IN1(n14330), .IN2(n18330), .IN3(n14331), .IN4(n17838), .Q(
        n17689) );
  AO22X1 U25793 ( .IN1(n14330), .IN2(n18332), .IN3(n14331), .IN4(n18637), .Q(
        n17690) );
  AO22X1 U25794 ( .IN1(n14330), .IN2(n18333), .IN3(n14331), .IN4(n17789), .Q(
        n17691) );
  AO22X1 U25795 ( .IN1(n14330), .IN2(n18319), .IN3(n14331), .IN4(n17866), .Q(
        n17692) );
  AO22X1 U25796 ( .IN1(n14330), .IN2(n18320), .IN3(n14331), .IN4(n17878), .Q(
        n17693) );
  AO22X1 U25797 ( .IN1(n14330), .IN2(n18323), .IN3(n14331), .IN4(n18649), .Q(
        n17694) );
  AO22X1 U25798 ( .IN1(n14330), .IN2(n18324), .IN3(n14331), .IN4(n17851), .Q(
        n17695) );
  AO22X1 U25799 ( .IN1(n14330), .IN2(n18327), .IN3(n14331), .IN4(n18661), .Q(
        n17696) );
  AO22X1 U25800 ( .IN1(n14330), .IN2(n18328), .IN3(n14331), .IN4(n17847), .Q(
        n17697) );
  AO22X1 U25801 ( .IN1(n14330), .IN2(n18331), .IN3(n14331), .IN4(n17855), .Q(
        n17698) );
  NAND2X0 U25802 ( .IN1(n2846), .IN2(n13944), .QN(n13976) );
  OA21X1 U25803 ( .IN1(n13445), .IN2(n13476), .IN3(n13443), .Q(n13440) );
  OA21X1 U25804 ( .IN1(n13460), .IN2(n13457), .IN3(n13462), .Q(n13476) );
  OA21X1 U25805 ( .IN1(n10970), .IN2(n11001), .IN3(n10968), .Q(n10965) );
  OA21X1 U25806 ( .IN1(n10985), .IN2(n10982), .IN3(n10987), .Q(n11001) );
  OA21X1 U25807 ( .IN1(n10351), .IN2(n10382), .IN3(n10349), .Q(n10346) );
  OA21X1 U25808 ( .IN1(n10366), .IN2(n10363), .IN3(n10368), .Q(n10382) );
  OA21X1 U25809 ( .IN1(n9731), .IN2(n9762), .IN3(n9729), .Q(n9726) );
  OA21X1 U25810 ( .IN1(n9746), .IN2(n9743), .IN3(n9748), .Q(n9762) );
  OA21X1 U25811 ( .IN1(n13754), .IN2(n13785), .IN3(n13752), .Q(n13749) );
  OA21X1 U25812 ( .IN1(n13769), .IN2(n13766), .IN3(n13771), .Q(n13785) );
  OA21X1 U25813 ( .IN1(n11279), .IN2(n11310), .IN3(n11277), .Q(n11274) );
  OA21X1 U25814 ( .IN1(n11294), .IN2(n11291), .IN3(n11296), .Q(n11310) );
  OA21X1 U25815 ( .IN1(n13136), .IN2(n13167), .IN3(n13134), .Q(n13131) );
  OA21X1 U25816 ( .IN1(n13151), .IN2(n13148), .IN3(n13153), .Q(n13167) );
  OA21X1 U25817 ( .IN1(n12827), .IN2(n12858), .IN3(n12825), .Q(n12822) );
  OA21X1 U25818 ( .IN1(n12842), .IN2(n12839), .IN3(n12844), .Q(n12858) );
  OA21X1 U25819 ( .IN1(n10660), .IN2(n10691), .IN3(n10658), .Q(n10655) );
  OA21X1 U25820 ( .IN1(n10675), .IN2(n10672), .IN3(n10677), .Q(n10691) );
  OA21X1 U25821 ( .IN1(n12518), .IN2(n12549), .IN3(n12516), .Q(n12513) );
  OA21X1 U25822 ( .IN1(n12533), .IN2(n12530), .IN3(n12535), .Q(n12549) );
  OA21X1 U25823 ( .IN1(n12209), .IN2(n12240), .IN3(n12207), .Q(n12204) );
  OA21X1 U25824 ( .IN1(n12224), .IN2(n12221), .IN3(n12226), .Q(n12240) );
  OA21X1 U25825 ( .IN1(n10041), .IN2(n10072), .IN3(n10039), .Q(n10036) );
  OA21X1 U25826 ( .IN1(n10056), .IN2(n10053), .IN3(n10058), .Q(n10072) );
  OA21X1 U25827 ( .IN1(n11899), .IN2(n11930), .IN3(n11897), .Q(n11894) );
  OA21X1 U25828 ( .IN1(n11914), .IN2(n11911), .IN3(n11916), .Q(n11930) );
  OA21X1 U25829 ( .IN1(n11589), .IN2(n11620), .IN3(n11587), .Q(n11584) );
  OA21X1 U25830 ( .IN1(n11604), .IN2(n11601), .IN3(n11606), .Q(n11620) );
  OA21X1 U25831 ( .IN1(n9420), .IN2(n9451), .IN3(n9418), .Q(n9415) );
  OA21X1 U25832 ( .IN1(n9435), .IN2(n9432), .IN3(n9437), .Q(n9451) );
  OA21X1 U25833 ( .IN1(n14018), .IN2(n14049), .IN3(n14016), .Q(n14013) );
  OA21X1 U25834 ( .IN1(n14033), .IN2(n14030), .IN3(n14035), .Q(n14049) );
  NAND4X0 U25835 ( .IN1(n17105), .IN2(n17106), .IN3(n17107), .IN4(n17108), 
        .QN(s15_addr_o[24]) );
  OA22X1 U25836 ( .IN1(n1765), .IN2(n19637), .IN3(n1661), .IN4(n19619), .Q(
        n17105) );
  OA22X1 U25837 ( .IN1(n1937), .IN2(n19670), .IN3(n1851), .IN4(n19652), .Q(
        n17106) );
  OA22X1 U25838 ( .IN1(n2109), .IN2(n19703), .IN3(n2023), .IN4(n19685), .Q(
        n17107) );
  NAND4X0 U25839 ( .IN1(n17109), .IN2(n17110), .IN3(n17111), .IN4(n17112), 
        .QN(s15_addr_o[26]) );
  OA22X1 U25840 ( .IN1(n1763), .IN2(n19637), .IN3(n1659), .IN4(n19619), .Q(
        n17109) );
  OA22X1 U25841 ( .IN1(n1935), .IN2(n19670), .IN3(n1849), .IN4(n19652), .Q(
        n17110) );
  OA22X1 U25842 ( .IN1(n2107), .IN2(n19703), .IN3(n2021), .IN4(n19685), .Q(
        n17111) );
  NAND4X0 U25843 ( .IN1(n17113), .IN2(n17114), .IN3(n17115), .IN4(n17116), 
        .QN(s15_addr_o[25]) );
  OA22X1 U25844 ( .IN1(n1764), .IN2(n19637), .IN3(n1660), .IN4(n19619), .Q(
        n17113) );
  OA22X1 U25845 ( .IN1(n1936), .IN2(n19670), .IN3(n1850), .IN4(n19652), .Q(
        n17114) );
  OA22X1 U25846 ( .IN1(n2108), .IN2(n19703), .IN3(n2022), .IN4(n19685), .Q(
        n17115) );
  NAND4X0 U25847 ( .IN1(n17091), .IN2(n17092), .IN3(n17093), .IN4(n17094), 
        .QN(s15_stb_o) );
  OA22X1 U25848 ( .IN1(n1795), .IN2(n16406), .IN3(n1709), .IN4(n16711), .Q(
        n17091) );
  OA22X1 U25849 ( .IN1(n1967), .IN2(n15796), .IN3(n1881), .IN4(n16101), .Q(
        n17092) );
  OA22X1 U25850 ( .IN1(n2139), .IN2(n15186), .IN3(n2053), .IN4(n15491), .Q(
        n17093) );
  NAND4X0 U25851 ( .IN1(n17087), .IN2(n17088), .IN3(n17089), .IN4(n17090), 
        .QN(s15_addr_o[27]) );
  OA22X1 U25852 ( .IN1(n1762), .IN2(n19637), .IN3(n1658), .IN4(n19620), .Q(
        n17087) );
  OA22X1 U25853 ( .IN1(n1934), .IN2(n19670), .IN3(n1848), .IN4(n19653), .Q(
        n17088) );
  OA22X1 U25854 ( .IN1(n2106), .IN2(n19703), .IN3(n2020), .IN4(n19686), .Q(
        n17089) );
  OA21X1 U25855 ( .IN1(n13788), .IN2(n13772), .IN3(n13774), .Q(n13766) );
  OA21X1 U25856 ( .IN1(n13479), .IN2(n13463), .IN3(n13465), .Q(n13457) );
  OA21X1 U25857 ( .IN1(n11313), .IN2(n11297), .IN3(n11299), .Q(n11291) );
  OA21X1 U25858 ( .IN1(n13170), .IN2(n13154), .IN3(n13156), .Q(n13148) );
  OA21X1 U25859 ( .IN1(n12861), .IN2(n12845), .IN3(n12847), .Q(n12839) );
  OA21X1 U25860 ( .IN1(n11004), .IN2(n10988), .IN3(n10990), .Q(n10982) );
  OA21X1 U25861 ( .IN1(n10694), .IN2(n10678), .IN3(n10680), .Q(n10672) );
  OA21X1 U25862 ( .IN1(n12552), .IN2(n12536), .IN3(n12538), .Q(n12530) );
  OA21X1 U25863 ( .IN1(n12243), .IN2(n12227), .IN3(n12229), .Q(n12221) );
  OA21X1 U25864 ( .IN1(n10385), .IN2(n10369), .IN3(n10371), .Q(n10363) );
  OA21X1 U25865 ( .IN1(n10075), .IN2(n10059), .IN3(n10061), .Q(n10053) );
  OA21X1 U25866 ( .IN1(n11933), .IN2(n11917), .IN3(n11919), .Q(n11911) );
  OA21X1 U25867 ( .IN1(n11623), .IN2(n11607), .IN3(n11609), .Q(n11601) );
  OA21X1 U25868 ( .IN1(n9765), .IN2(n9749), .IN3(n9751), .Q(n9743) );
  OA21X1 U25869 ( .IN1(n9454), .IN2(n9438), .IN3(n9440), .Q(n9432) );
  OA21X1 U25870 ( .IN1(n14052), .IN2(n14036), .IN3(n14038), .Q(n14030) );
  INVX0 U25871 ( .IN(n14141), .QN(n3382) );
  OA21X1 U25872 ( .IN1(n13799), .IN2(n13786), .IN3(n13773), .Q(n13788) );
  OA21X1 U25873 ( .IN1(n13490), .IN2(n13477), .IN3(n13464), .Q(n13479) );
  OA21X1 U25874 ( .IN1(n11324), .IN2(n11311), .IN3(n11298), .Q(n11313) );
  OA21X1 U25875 ( .IN1(n13181), .IN2(n13168), .IN3(n13155), .Q(n13170) );
  OA21X1 U25876 ( .IN1(n12872), .IN2(n12859), .IN3(n12846), .Q(n12861) );
  OA21X1 U25877 ( .IN1(n11015), .IN2(n11002), .IN3(n10989), .Q(n11004) );
  OA21X1 U25878 ( .IN1(n10705), .IN2(n10692), .IN3(n10679), .Q(n10694) );
  OA21X1 U25879 ( .IN1(n12563), .IN2(n12550), .IN3(n12537), .Q(n12552) );
  OA21X1 U25880 ( .IN1(n12254), .IN2(n12241), .IN3(n12228), .Q(n12243) );
  OA21X1 U25881 ( .IN1(n10396), .IN2(n10383), .IN3(n10370), .Q(n10385) );
  OA21X1 U25882 ( .IN1(n10086), .IN2(n10073), .IN3(n10060), .Q(n10075) );
  OA21X1 U25883 ( .IN1(n11944), .IN2(n11931), .IN3(n11918), .Q(n11933) );
  OA21X1 U25884 ( .IN1(n11634), .IN2(n11621), .IN3(n11608), .Q(n11623) );
  OA21X1 U25885 ( .IN1(n9776), .IN2(n9763), .IN3(n9750), .Q(n9765) );
  OA21X1 U25886 ( .IN1(n9465), .IN2(n9452), .IN3(n9439), .Q(n9454) );
  OA21X1 U25887 ( .IN1(n14063), .IN2(n14050), .IN3(n14037), .Q(n14052) );
  NAND3X0 U25888 ( .IN1(n17117), .IN2(n17118), .IN3(n4210), .QN(n7172) );
  NAND3X0 U25889 ( .IN1(n4210), .IN2(n17118), .IN3(n4205), .QN(n7174) );
  NAND3X0 U25890 ( .IN1(n4210), .IN2(n17117), .IN3(n4211), .QN(n7176) );
  OA22X1 U25891 ( .IN1(n2281), .IN2(n19736), .IN3(n2195), .IN4(n19718), .Q(
        n17108) );
  OA22X1 U25892 ( .IN1(n2280), .IN2(n19736), .IN3(n2194), .IN4(n19718), .Q(
        n17116) );
  OA22X1 U25893 ( .IN1(n2279), .IN2(n19736), .IN3(n2193), .IN4(n19718), .Q(
        n17112) );
  OA22X1 U25894 ( .IN1(n2278), .IN2(n19736), .IN3(n2192), .IN4(n19719), .Q(
        n17090) );
  OA22X1 U25895 ( .IN1(n2311), .IN2(n14496), .IN3(n2225), .IN4(n14881), .Q(
        n17094) );
  INVX0 U25896 ( .IN(n17118), .QN(n4211) );
  INVX0 U25897 ( .IN(n17119), .QN(n4210) );
  INVX0 U25898 ( .IN(n17117), .QN(n4205) );
  NAND2X0 U25899 ( .IN1(n17939), .IN2(n18150), .QN(n14070) );
  NAND2X0 U25900 ( .IN1(n18088), .IN2(n17975), .QN(n14075) );
  NAND2X0 U25901 ( .IN1(n18086), .IN2(n17974), .QN(n14072) );
  NAND2X0 U25902 ( .IN1(n18095), .IN2(n17968), .QN(n13647) );
  NAND2X0 U25903 ( .IN1(n17985), .IN2(n18106), .QN(n13338) );
  NAND2X0 U25904 ( .IN1(n17986), .IN2(n18108), .QN(n11172) );
  NAND2X0 U25905 ( .IN1(n18096), .IN2(n17970), .QN(n12411) );
  NAND2X0 U25906 ( .IN1(n17987), .IN2(n18110), .QN(n12102) );
  NAND2X0 U25907 ( .IN1(n18097), .IN2(n17972), .QN(n9624) );
  NAND2X0 U25908 ( .IN1(n17988), .IN2(n18112), .QN(n9313) );
  NAND2X0 U25909 ( .IN1(n18089), .IN2(n17969), .QN(n13644) );
  NAND2X0 U25910 ( .IN1(n17977), .IN2(n18107), .QN(n13335) );
  NAND2X0 U25911 ( .IN1(n17979), .IN2(n18109), .QN(n11169) );
  NAND2X0 U25912 ( .IN1(n18091), .IN2(n17971), .QN(n12408) );
  NAND2X0 U25913 ( .IN1(n17981), .IN2(n18111), .QN(n12099) );
  NAND2X0 U25914 ( .IN1(n18093), .IN2(n17973), .QN(n9621) );
  NAND2X0 U25915 ( .IN1(n17983), .IN2(n18113), .QN(n9310) );
  NAND2X0 U25916 ( .IN1(n18122), .IN2(n17997), .QN(n13029) );
  NAND2X0 U25917 ( .IN1(n18123), .IN2(n17999), .QN(n10863) );
  NAND2X0 U25918 ( .IN1(n18124), .IN2(n18001), .QN(n10244) );
  NAND2X0 U25919 ( .IN1(n18125), .IN2(n18003), .QN(n11792) );
  NAND2X0 U25920 ( .IN1(n18114), .IN2(n17998), .QN(n13026) );
  NAND2X0 U25921 ( .IN1(n18116), .IN2(n18000), .QN(n10860) );
  NAND2X0 U25922 ( .IN1(n18118), .IN2(n18002), .QN(n10241) );
  NAND2X0 U25923 ( .IN1(n18120), .IN2(n18004), .QN(n11789) );
  NAND2X0 U25924 ( .IN1(n18013), .IN2(n18134), .QN(n12720) );
  NAND2X0 U25925 ( .IN1(n18014), .IN2(n18136), .QN(n10553) );
  NAND2X0 U25926 ( .IN1(n18015), .IN2(n18138), .QN(n9934) );
  NAND2X0 U25927 ( .IN1(n18016), .IN2(n18140), .QN(n11482) );
  NAND2X0 U25928 ( .IN1(n18005), .IN2(n18135), .QN(n12717) );
  NAND2X0 U25929 ( .IN1(n18007), .IN2(n18137), .QN(n10550) );
  NAND2X0 U25930 ( .IN1(n18009), .IN2(n18139), .QN(n9931) );
  NAND2X0 U25931 ( .IN1(n18011), .IN2(n18141), .QN(n11479) );
  NAND2X0 U25932 ( .IN1(n18098), .IN2(n18024), .QN(n14074) );
  NAND2X0 U25933 ( .IN1(n18099), .IN2(n18021), .QN(n13650) );
  NAND2X0 U25934 ( .IN1(n17989), .IN2(n18142), .QN(n13341) );
  NAND2X0 U25935 ( .IN1(n17990), .IN2(n18143), .QN(n11175) );
  NAND2X0 U25936 ( .IN1(n18100), .IN2(n18022), .QN(n12414) );
  NAND2X0 U25937 ( .IN1(n17991), .IN2(n18144), .QN(n12105) );
  NAND2X0 U25938 ( .IN1(n18101), .IN2(n18023), .QN(n9627) );
  NAND2X0 U25939 ( .IN1(n17992), .IN2(n18145), .QN(n9316) );
  NAND2X0 U25940 ( .IN1(n18126), .IN2(n18025), .QN(n13032) );
  NAND2X0 U25941 ( .IN1(n18127), .IN2(n18026), .QN(n10866) );
  NAND2X0 U25942 ( .IN1(n18128), .IN2(n18027), .QN(n10247) );
  NAND2X0 U25943 ( .IN1(n18129), .IN2(n18028), .QN(n11795) );
  NAND2X0 U25944 ( .IN1(n18017), .IN2(n18146), .QN(n12723) );
  NAND2X0 U25945 ( .IN1(n18018), .IN2(n18147), .QN(n10556) );
  NAND2X0 U25946 ( .IN1(n18019), .IN2(n18148), .QN(n9937) );
  NAND2X0 U25947 ( .IN1(n18020), .IN2(n18149), .QN(n11485) );
  INVX0 U25948 ( .IN(n14187), .QN(n3381) );
  NAND4X0 U25949 ( .IN1(n14308), .IN2(n14309), .IN3(n14310), .IN4(n14311), 
        .QN(s15_addr_o[2]) );
  OA22X1 U25950 ( .IN1(n1787), .IN2(n19638), .IN3(n1701), .IN4(n19621), .Q(
        n14308) );
  OA22X1 U25951 ( .IN1(n1959), .IN2(n19671), .IN3(n1873), .IN4(n19654), .Q(
        n14309) );
  OA22X1 U25952 ( .IN1(n2131), .IN2(n19704), .IN3(n2045), .IN4(n19687), .Q(
        n14310) );
  NAND4X0 U25953 ( .IN1(n14316), .IN2(n14317), .IN3(n14318), .IN4(n14319), 
        .QN(s15_addr_o[3]) );
  OA22X1 U25954 ( .IN1(n1786), .IN2(n19638), .IN3(n1699), .IN4(n19620), .Q(
        n14316) );
  OA22X1 U25955 ( .IN1(n1958), .IN2(n19671), .IN3(n1872), .IN4(n19653), .Q(
        n14317) );
  OA22X1 U25956 ( .IN1(n2130), .IN2(n19704), .IN3(n2044), .IN4(n19686), .Q(
        n14318) );
  NAND4X0 U25957 ( .IN1(n14320), .IN2(n14321), .IN3(n14322), .IN4(n14323), 
        .QN(s15_addr_o[4]) );
  OA22X1 U25958 ( .IN1(n1785), .IN2(n19638), .IN3(n1697), .IN4(n19620), .Q(
        n14320) );
  OA22X1 U25959 ( .IN1(n1957), .IN2(n19671), .IN3(n1871), .IN4(n19653), .Q(
        n14321) );
  OA22X1 U25960 ( .IN1(n2129), .IN2(n19704), .IN3(n2043), .IN4(n19686), .Q(
        n14322) );
  NAND4X0 U25961 ( .IN1(n14312), .IN2(n14313), .IN3(n14314), .IN4(n14315), 
        .QN(s15_addr_o[5]) );
  OA22X1 U25962 ( .IN1(n1784), .IN2(n19638), .IN3(n1696), .IN4(n19621), .Q(
        n14312) );
  OA22X1 U25963 ( .IN1(n1956), .IN2(n19671), .IN3(n1870), .IN4(n19654), .Q(
        n14313) );
  OA22X1 U25964 ( .IN1(n2128), .IN2(n19704), .IN3(n2042), .IN4(n19687), .Q(
        n14314) );
  NOR2X0 U25965 ( .IN1(n2274), .IN2(n2277), .QN(n14831) );
  NOR2X0 U25966 ( .IN1(n2102), .IN2(n2105), .QN(n15478) );
  NOR2X0 U25967 ( .IN1(n1930), .IN2(n1933), .QN(n16088) );
  NOR2X0 U25968 ( .IN1(n1758), .IN2(n1761), .QN(n16698) );
  NOR2X0 U25969 ( .IN1(n1650), .IN2(n1657), .QN(n17024) );
  NOR2X0 U25970 ( .IN1(n2188), .IN2(n2191), .QN(n15173) );
  NOR2X0 U25971 ( .IN1(n2016), .IN2(n2019), .QN(n15783) );
  NOR2X0 U25972 ( .IN1(n1844), .IN2(n1847), .QN(n16393) );
  NOR2X0 U25973 ( .IN1(n2276), .IN2(n2275), .QN(n14822) );
  NOR2X0 U25974 ( .IN1(n2104), .IN2(n2103), .QN(n15475) );
  NOR2X0 U25975 ( .IN1(n1932), .IN2(n1931), .QN(n16085) );
  NOR2X0 U25976 ( .IN1(n1760), .IN2(n1759), .QN(n16695) );
  NOR2X0 U25977 ( .IN1(n2190), .IN2(n2189), .QN(n15170) );
  NOR2X0 U25978 ( .IN1(n2018), .IN2(n2017), .QN(n15780) );
  NOR2X0 U25979 ( .IN1(n1846), .IN2(n1845), .QN(n16390) );
  NOR2X0 U25980 ( .IN1(n1656), .IN2(n1655), .QN(n17007) );
  NAND3X0 U25981 ( .IN1(n17119), .IN2(n17118), .IN3(n4205), .QN(n7173) );
  NAND3X0 U25982 ( .IN1(n17117), .IN2(n17118), .IN3(n17119), .QN(n7171) );
  NAND3X0 U25983 ( .IN1(n17119), .IN2(n17117), .IN3(n4211), .QN(n7175) );
  NAND3X0 U25984 ( .IN1(n4205), .IN2(n17119), .IN3(n4211), .QN(n7177) );
  OA221X1 U25985 ( .IN1(n18426), .IN2(n18145), .IN3(n18422), .IN4(n18023), 
        .IN5(n9289), .Q(n9286) );
  OA22X1 U25986 ( .IN1(n18414), .IN2(n18027), .IN3(n18418), .IN4(n18148), .Q(
        n9289) );
  OA221X1 U25987 ( .IN1(n18426), .IN2(n17992), .IN3(n18422), .IN4(n18101), 
        .IN5(n9280), .Q(n9277) );
  OA22X1 U25988 ( .IN1(n18414), .IN2(n18128), .IN3(n18418), .IN4(n18019), .Q(
        n9280) );
  OA221X1 U25989 ( .IN1(n18426), .IN2(n18112), .IN3(n18422), .IN4(n17972), 
        .IN5(n9271), .Q(n9268) );
  OA22X1 U25990 ( .IN1(n18414), .IN2(n18001), .IN3(n18418), .IN4(n18138), .Q(
        n9271) );
  OA221X1 U25991 ( .IN1(n18426), .IN2(n17988), .IN3(n18422), .IN4(n18097), 
        .IN5(n9262), .Q(n9259) );
  OA22X1 U25992 ( .IN1(n18414), .IN2(n18124), .IN3(n18418), .IN4(n18015), .Q(
        n9262) );
  OA221X1 U25993 ( .IN1(n18426), .IN2(n18113), .IN3(n18422), .IN4(n17973), 
        .IN5(n9253), .Q(n9250) );
  OA22X1 U25994 ( .IN1(n18414), .IN2(n18002), .IN3(n18418), .IN4(n18139), .Q(
        n9253) );
  OA221X1 U25995 ( .IN1(n18426), .IN2(n17983), .IN3(n18422), .IN4(n18093), 
        .IN5(n9244), .Q(n9241) );
  OA22X1 U25996 ( .IN1(n18414), .IN2(n18118), .IN3(n18418), .IN4(n18009), .Q(
        n9244) );
  OA221X1 U25997 ( .IN1(n18427), .IN2(n18105), .IN3(n18423), .IN4(n17967), 
        .IN5(n9235), .Q(n9232) );
  OA22X1 U25998 ( .IN1(n18415), .IN2(n17995), .IN3(n18419), .IN4(n18132), .Q(
        n9235) );
  OA221X1 U25999 ( .IN1(n18427), .IN2(n17984), .IN3(n18423), .IN4(n18094), 
        .IN5(n9226), .Q(n9223) );
  OA22X1 U26000 ( .IN1(n18415), .IN2(n18119), .IN3(n18419), .IN4(n18010), .Q(
        n9226) );
  OA221X1 U26001 ( .IN1(n18427), .IN2(n18065), .IN3(n18423), .IN4(n17940), 
        .IN5(n9217), .Q(n9214) );
  OA22X1 U26002 ( .IN1(n18415), .IN2(n17937), .IN3(n18419), .IN4(n18084), .Q(
        n9217) );
  OA221X1 U26003 ( .IN1(n18427), .IN2(n17933), .IN3(n18423), .IN4(n18153), 
        .IN5(n9208), .Q(n9205) );
  OA22X1 U26004 ( .IN1(n18415), .IN2(n18061), .IN3(n18419), .IN4(n17957), .Q(
        n9208) );
  OA221X1 U26005 ( .IN1(n18427), .IN2(n17944), .IN3(n18423), .IN4(n18068), 
        .IN5(n9199), .Q(n9196) );
  OA22X1 U26006 ( .IN1(n18415), .IN2(n18073), .IN3(n18419), .IN4(n17955), .Q(
        n9199) );
  OA221X1 U26007 ( .IN1(n18427), .IN2(n18078), .IN3(n18423), .IN4(n17952), 
        .IN5(n9190), .Q(n9187) );
  OA22X1 U26008 ( .IN1(n18415), .IN2(n17962), .IN3(n18419), .IN4(n18081), .Q(
        n9190) );
  OA221X1 U26009 ( .IN1(n18427), .IN2(n18200), .IN3(n18423), .IN4(n18031), 
        .IN5(n9181), .Q(n9178) );
  OA22X1 U26010 ( .IN1(n18415), .IN2(n18047), .IN3(n18419), .IN4(n18215), .Q(
        n9181) );
  OA221X1 U26011 ( .IN1(n18427), .IN2(n18044), .IN3(n18423), .IN4(n18196), 
        .IN5(n9172), .Q(n9169) );
  OA22X1 U26012 ( .IN1(n18415), .IN2(n18211), .IN3(n18419), .IN4(n18059), .Q(
        n9172) );
  OA221X1 U26013 ( .IN1(n18427), .IN2(n18204), .IN3(n18423), .IN4(n18034), 
        .IN5(n9163), .Q(n9160) );
  OA22X1 U26014 ( .IN1(n18415), .IN2(n18051), .IN3(n18419), .IN4(n18219), .Q(
        n9163) );
  OA221X1 U26015 ( .IN1(n18427), .IN2(n18040), .IN3(n18423), .IN4(n18193), 
        .IN5(n9144), .Q(n9135) );
  OA22X1 U26016 ( .IN1(n18415), .IN2(n18207), .IN3(n18419), .IN4(n18055), .Q(
        n9144) );
  OA221X1 U26017 ( .IN1(n18402), .IN2(n18143), .IN3(n18334), .IN4(n18024), 
        .IN5(n9288), .Q(n9287) );
  OA22X1 U26018 ( .IN1(n18406), .IN2(n18026), .IN3(n18410), .IN4(n18147), .Q(
        n9288) );
  OA221X1 U26019 ( .IN1(n18402), .IN2(n17990), .IN3(n18334), .IN4(n18098), 
        .IN5(n9279), .Q(n9278) );
  OA22X1 U26020 ( .IN1(n18406), .IN2(n18127), .IN3(n18410), .IN4(n18018), .Q(
        n9279) );
  OA221X1 U26021 ( .IN1(n18402), .IN2(n18108), .IN3(n18334), .IN4(n17975), 
        .IN5(n9270), .Q(n9269) );
  OA22X1 U26022 ( .IN1(n18406), .IN2(n17999), .IN3(n18410), .IN4(n18136), .Q(
        n9270) );
  OA221X1 U26023 ( .IN1(n18402), .IN2(n17986), .IN3(n18334), .IN4(n18088), 
        .IN5(n9261), .Q(n9260) );
  OA22X1 U26024 ( .IN1(n18406), .IN2(n18123), .IN3(n18410), .IN4(n18014), .Q(
        n9261) );
  OA221X1 U26025 ( .IN1(n18402), .IN2(n18109), .IN3(n18334), .IN4(n17974), 
        .IN5(n9252), .Q(n9251) );
  OA22X1 U26026 ( .IN1(n18406), .IN2(n18000), .IN3(n18410), .IN4(n18137), .Q(
        n9252) );
  OA221X1 U26027 ( .IN1(n18402), .IN2(n17979), .IN3(n18334), .IN4(n18086), 
        .IN5(n9243), .Q(n9242) );
  OA22X1 U26028 ( .IN1(n18406), .IN2(n18116), .IN3(n18410), .IN4(n18007), .Q(
        n9243) );
  OA221X1 U26029 ( .IN1(n18403), .IN2(n18103), .IN3(n18335), .IN4(n17976), 
        .IN5(n9234), .Q(n9233) );
  OA22X1 U26030 ( .IN1(n18407), .IN2(n17994), .IN3(n18411), .IN4(n18131), .Q(
        n9234) );
  OA221X1 U26031 ( .IN1(n18403), .IN2(n17980), .IN3(n18335), .IN4(n18087), 
        .IN5(n9225), .Q(n9224) );
  OA22X1 U26032 ( .IN1(n18407), .IN2(n18117), .IN3(n18411), .IN4(n18008), .Q(
        n9225) );
  OA221X1 U26033 ( .IN1(n18403), .IN2(n17948), .IN3(n18335), .IN4(n18150), 
        .IN5(n9216), .Q(n9215) );
  OA22X1 U26034 ( .IN1(n18407), .IN2(n17936), .IN3(n18411), .IN4(n18083), .Q(
        n9216) );
  OA221X1 U26035 ( .IN1(n18403), .IN2(n18156), .IN3(n18335), .IN4(n17939), 
        .IN5(n9207), .Q(n9206) );
  OA22X1 U26036 ( .IN1(n18407), .IN2(n18062), .IN3(n18411), .IN4(n17958), .Q(
        n9207) );
  OA221X1 U26037 ( .IN1(n18403), .IN2(n17942), .IN3(n18335), .IN4(n18070), 
        .IN5(n9198), .Q(n9197) );
  OA22X1 U26038 ( .IN1(n18407), .IN2(n18072), .IN3(n18411), .IN4(n17954), .Q(
        n9198) );
  OA221X1 U26039 ( .IN1(n18403), .IN2(n18076), .IN3(n18335), .IN4(n17949), 
        .IN5(n9189), .Q(n9188) );
  OA22X1 U26040 ( .IN1(n18407), .IN2(n17961), .IN3(n18411), .IN4(n18080), .Q(
        n9189) );
  OA221X1 U26041 ( .IN1(n18403), .IN2(n18198), .IN3(n18335), .IN4(n18035), 
        .IN5(n9180), .Q(n9179) );
  OA22X1 U26042 ( .IN1(n18407), .IN2(n18046), .IN3(n18411), .IN4(n18214), .Q(
        n9180) );
  OA221X1 U26043 ( .IN1(n18403), .IN2(n18042), .IN3(n18335), .IN4(n18190), 
        .IN5(n9171), .Q(n9170) );
  OA22X1 U26044 ( .IN1(n18407), .IN2(n18210), .IN3(n18411), .IN4(n18058), .Q(
        n9171) );
  OA221X1 U26045 ( .IN1(n18403), .IN2(n18202), .IN3(n18335), .IN4(n18036), 
        .IN5(n9162), .Q(n9161) );
  OA22X1 U26046 ( .IN1(n18407), .IN2(n18050), .IN3(n18411), .IN4(n18218), .Q(
        n9162) );
  OA221X1 U26047 ( .IN1(n18403), .IN2(n18038), .IN3(n18335), .IN4(n18189), 
        .IN5(n9139), .Q(n9136) );
  OA22X1 U26048 ( .IN1(n18407), .IN2(n18206), .IN3(n18411), .IN4(n18054), .Q(
        n9139) );
  NOR2X0 U26049 ( .IN1(n18430), .IN2(n18334), .QN(n14208) );
  NOR2X0 U26050 ( .IN1(n18430), .IN2(n18402), .QN(n11459) );
  NOR2X0 U26051 ( .IN1(n18430), .IN2(n18406), .QN(n11150) );
  NOR2X0 U26052 ( .IN1(n18430), .IN2(n18410), .QN(n10840) );
  NOR2X0 U26053 ( .IN1(n18430), .IN2(n18414), .QN(n10531) );
  NOR2X0 U26054 ( .IN1(n18430), .IN2(n18418), .QN(n10221) );
  NOR2X0 U26055 ( .IN1(n18430), .IN2(n18422), .QN(n9911) );
  NOR2X0 U26056 ( .IN1(n18430), .IN2(n18426), .QN(n9600) );
  NOR2X0 U26057 ( .IN1(n18430), .IN2(n18370), .QN(n13934) );
  NOR2X0 U26058 ( .IN1(n18430), .IN2(n18374), .QN(n13625) );
  NOR2X0 U26059 ( .IN1(n18430), .IN2(n18378), .QN(n13316) );
  NOR2X0 U26060 ( .IN1(n18430), .IN2(n18382), .QN(n13007) );
  NOR2X0 U26061 ( .IN1(n18430), .IN2(n18386), .QN(n12698) );
  NOR2X0 U26062 ( .IN1(n18430), .IN2(n18390), .QN(n12389) );
  NOR2X0 U26063 ( .IN1(n18430), .IN2(n18394), .QN(n12079) );
  NOR2X0 U26064 ( .IN1(n18430), .IN2(n18398), .QN(n11769) );
  OA22X1 U26065 ( .IN1(n2303), .IN2(n19737), .IN3(n2217), .IN4(n19720), .Q(
        n14311) );
  OA22X1 U26066 ( .IN1(n2302), .IN2(n19737), .IN3(n2216), .IN4(n19719), .Q(
        n14319) );
  OA22X1 U26067 ( .IN1(n2301), .IN2(n19737), .IN3(n2215), .IN4(n19719), .Q(
        n14323) );
  OA22X1 U26068 ( .IN1(n2300), .IN2(n19737), .IN3(n2214), .IN4(n19720), .Q(
        n14315) );
  OA22X1 U26069 ( .IN1(n18379), .IN2(n17993), .IN3(n18383), .IN4(n18130), .Q(
        n9236) );
  OA22X1 U26070 ( .IN1(n18395), .IN2(n17996), .IN3(n18399), .IN4(n18133), .Q(
        n9237) );
  OA22X1 U26071 ( .IN1(n18379), .IN2(n18115), .IN3(n18383), .IN4(n18006), .Q(
        n9227) );
  OA22X1 U26072 ( .IN1(n18395), .IN2(n18121), .IN3(n18399), .IN4(n18012), .Q(
        n9228) );
  OA22X1 U26073 ( .IN1(n18379), .IN2(n17935), .IN3(n18383), .IN4(n18066), .Q(
        n9218) );
  OA22X1 U26074 ( .IN1(n18395), .IN2(n17938), .IN3(n18399), .IN4(n18085), .Q(
        n9219) );
  OA22X1 U26075 ( .IN1(n18379), .IN2(n18063), .IN3(n18383), .IN4(n17934), .Q(
        n9209) );
  OA22X1 U26076 ( .IN1(n18395), .IN2(n18064), .IN3(n18399), .IN4(n17959), .Q(
        n9210) );
  OA22X1 U26077 ( .IN1(n18379), .IN2(n18071), .IN3(n18383), .IN4(n17953), .Q(
        n9200) );
  OA22X1 U26078 ( .IN1(n18395), .IN2(n18074), .IN3(n18399), .IN4(n17956), .Q(
        n9201) );
  OA22X1 U26079 ( .IN1(n18379), .IN2(n17960), .IN3(n18383), .IN4(n18079), .Q(
        n9191) );
  OA22X1 U26080 ( .IN1(n18395), .IN2(n17963), .IN3(n18399), .IN4(n18082), .Q(
        n9192) );
  OA22X1 U26081 ( .IN1(n18379), .IN2(n18045), .IN3(n18383), .IN4(n18213), .Q(
        n9182) );
  OA22X1 U26082 ( .IN1(n18395), .IN2(n18048), .IN3(n18399), .IN4(n18216), .Q(
        n9183) );
  OA22X1 U26083 ( .IN1(n18379), .IN2(n18209), .IN3(n18383), .IN4(n18057), .Q(
        n9173) );
  OA22X1 U26084 ( .IN1(n18395), .IN2(n18212), .IN3(n18399), .IN4(n18060), .Q(
        n9174) );
  OA22X1 U26085 ( .IN1(n18379), .IN2(n18049), .IN3(n18383), .IN4(n18217), .Q(
        n9164) );
  OA22X1 U26086 ( .IN1(n18395), .IN2(n18052), .IN3(n18399), .IN4(n18220), .Q(
        n9165) );
  OA22X1 U26087 ( .IN1(n18379), .IN2(n18205), .IN3(n18383), .IN4(n18053), .Q(
        n9149) );
  OA22X1 U26088 ( .IN1(n18395), .IN2(n18208), .IN3(n18399), .IN4(n18056), .Q(
        n9154) );
  OA22X1 U26089 ( .IN1(n18378), .IN2(n18025), .IN3(n18382), .IN4(n18146), .Q(
        n9290) );
  OA22X1 U26090 ( .IN1(n18394), .IN2(n18028), .IN3(n18398), .IN4(n18149), .Q(
        n9291) );
  OA22X1 U26091 ( .IN1(n18378), .IN2(n18126), .IN3(n18382), .IN4(n18017), .Q(
        n9281) );
  OA22X1 U26092 ( .IN1(n18394), .IN2(n18129), .IN3(n18398), .IN4(n18020), .Q(
        n9282) );
  OA22X1 U26093 ( .IN1(n18378), .IN2(n17997), .IN3(n18382), .IN4(n18134), .Q(
        n9272) );
  OA22X1 U26094 ( .IN1(n18394), .IN2(n18003), .IN3(n18398), .IN4(n18140), .Q(
        n9273) );
  OA22X1 U26095 ( .IN1(n18378), .IN2(n18122), .IN3(n18382), .IN4(n18013), .Q(
        n9263) );
  OA22X1 U26096 ( .IN1(n18394), .IN2(n18125), .IN3(n18398), .IN4(n18016), .Q(
        n9264) );
  OA22X1 U26097 ( .IN1(n18378), .IN2(n17998), .IN3(n18382), .IN4(n18135), .Q(
        n9254) );
  OA22X1 U26098 ( .IN1(n18394), .IN2(n18004), .IN3(n18398), .IN4(n18141), .Q(
        n9255) );
  OA22X1 U26099 ( .IN1(n18378), .IN2(n18114), .IN3(n18382), .IN4(n18005), .Q(
        n9245) );
  OA22X1 U26100 ( .IN1(n18394), .IN2(n18120), .IN3(n18398), .IN4(n18011), .Q(
        n9246) );
  NAND2X0 U26101 ( .IN1(n18087), .IN2(n17976), .QN(n14073) );
  NAND2X0 U26102 ( .IN1(n18090), .IN2(n17965), .QN(n13641) );
  NAND2X0 U26103 ( .IN1(n17978), .IN2(n18102), .QN(n13332) );
  NAND2X0 U26104 ( .IN1(n17980), .IN2(n18103), .QN(n11166) );
  NAND2X0 U26105 ( .IN1(n18092), .IN2(n17966), .QN(n12405) );
  NAND2X0 U26106 ( .IN1(n17982), .IN2(n18104), .QN(n12096) );
  NAND2X0 U26107 ( .IN1(n18094), .IN2(n17967), .QN(n9618) );
  NAND2X0 U26108 ( .IN1(n17984), .IN2(n18105), .QN(n9307) );
  NAND2X0 U26109 ( .IN1(n18115), .IN2(n17993), .QN(n13023) );
  NAND2X0 U26110 ( .IN1(n18117), .IN2(n17994), .QN(n10857) );
  NAND2X0 U26111 ( .IN1(n18119), .IN2(n17995), .QN(n10238) );
  NAND2X0 U26112 ( .IN1(n18121), .IN2(n17996), .QN(n11786) );
  NAND2X0 U26113 ( .IN1(n18006), .IN2(n18130), .QN(n12714) );
  NAND2X0 U26114 ( .IN1(n18008), .IN2(n18131), .QN(n10547) );
  NAND2X0 U26115 ( .IN1(n18010), .IN2(n18132), .QN(n9928) );
  NAND2X0 U26116 ( .IN1(n18012), .IN2(n18133), .QN(n11476) );
  NAND4X0 U26117 ( .IN1(n9128), .IN2(n9129), .IN3(n9130), .IN4(n9131), .QN(
        s15_we_o) );
  OA22X1 U26118 ( .IN1(n1794), .IN2(n19639), .IN3(n1708), .IN4(n19631), .Q(
        n9128) );
  OA22X1 U26119 ( .IN1(n1966), .IN2(n19672), .IN3(n1880), .IN4(n19658), .Q(
        n9129) );
  OA22X1 U26120 ( .IN1(n2138), .IN2(n19705), .IN3(n2052), .IN4(n19691), .Q(
        n9130) );
  NAND4X0 U26121 ( .IN1(n7187), .IN2(n7188), .IN3(n7189), .IN4(n7190), .QN(
        s15_sel_o[0]) );
  OA22X1 U26122 ( .IN1(n1793), .IN2(n19644), .IN3(n1707), .IN4(n19631), .Q(
        n7187) );
  OA22X1 U26123 ( .IN1(n1965), .IN2(n19677), .IN3(n1879), .IN4(n19664), .Q(
        n7188) );
  OA22X1 U26124 ( .IN1(n2137), .IN2(n19710), .IN3(n2051), .IN4(n19697), .Q(
        n7189) );
  NAND4X0 U26125 ( .IN1(n7183), .IN2(n7184), .IN3(n7185), .IN4(n7186), .QN(
        s15_sel_o[1]) );
  OA22X1 U26126 ( .IN1(n1792), .IN2(n19644), .IN3(n1706), .IN4(n19631), .Q(
        n7183) );
  OA22X1 U26127 ( .IN1(n1964), .IN2(n19677), .IN3(n1878), .IN4(n19664), .Q(
        n7184) );
  OA22X1 U26128 ( .IN1(n2136), .IN2(n19710), .IN3(n2050), .IN4(n19697), .Q(
        n7185) );
  NAND4X0 U26129 ( .IN1(n7179), .IN2(n7180), .IN3(n7181), .IN4(n7182), .QN(
        s15_sel_o[2]) );
  OA22X1 U26130 ( .IN1(n1791), .IN2(n19644), .IN3(n1705), .IN4(n19631), .Q(
        n7179) );
  OA22X1 U26131 ( .IN1(n1963), .IN2(n19677), .IN3(n1877), .IN4(n19664), .Q(
        n7180) );
  OA22X1 U26132 ( .IN1(n2135), .IN2(n19710), .IN3(n2049), .IN4(n19697), .Q(
        n7181) );
  NAND4X0 U26133 ( .IN1(n7167), .IN2(n7168), .IN3(n7169), .IN4(n7170), .QN(
        s15_sel_o[3]) );
  OA22X1 U26134 ( .IN1(n1790), .IN2(n19639), .IN3(n1704), .IN4(n19631), .Q(
        n7167) );
  OA22X1 U26135 ( .IN1(n1962), .IN2(n19672), .IN3(n1876), .IN4(n19664), .Q(
        n7168) );
  OA22X1 U26136 ( .IN1(n2134), .IN2(n19705), .IN3(n2048), .IN4(n19697), .Q(
        n7169) );
  NAND4X0 U26137 ( .IN1(n7347), .IN2(n7348), .IN3(n7349), .IN4(n7350), .QN(
        s15_addr_o[0]) );
  OA22X1 U26138 ( .IN1(n1789), .IN2(n19641), .IN3(n1703), .IN4(n19629), .Q(
        n7347) );
  OA22X1 U26139 ( .IN1(n1961), .IN2(n19672), .IN3(n1875), .IN4(n19658), .Q(
        n7348) );
  OA22X1 U26140 ( .IN1(n2133), .IN2(n19705), .IN3(n2047), .IN4(n19691), .Q(
        n7349) );
  NAND4X0 U26141 ( .IN1(n7303), .IN2(n7304), .IN3(n7305), .IN4(n7306), .QN(
        s15_addr_o[1]) );
  OA22X1 U26142 ( .IN1(n1788), .IN2(n19642), .IN3(n1702), .IN4(n19626), .Q(
        n7303) );
  OA22X1 U26143 ( .IN1(n1960), .IN2(n19676), .IN3(n1874), .IN4(n19656), .Q(
        n7304) );
  OA22X1 U26144 ( .IN1(n2132), .IN2(n19709), .IN3(n2046), .IN4(n19689), .Q(
        n7305) );
  NAND4X0 U26145 ( .IN1(n7267), .IN2(n7268), .IN3(n7269), .IN4(n7270), .QN(
        s15_addr_o[6]) );
  OA22X1 U26146 ( .IN1(n1783), .IN2(n19640), .IN3(n1679), .IN4(n19631), .Q(
        n7267) );
  OA22X1 U26147 ( .IN1(n1955), .IN2(n19672), .IN3(n1869), .IN4(n19661), .Q(
        n7268) );
  OA22X1 U26148 ( .IN1(n2127), .IN2(n19705), .IN3(n2041), .IN4(n19694), .Q(
        n7269) );
  NAND4X0 U26149 ( .IN1(n7263), .IN2(n7264), .IN3(n7265), .IN4(n7266), .QN(
        s15_addr_o[7]) );
  OA22X1 U26150 ( .IN1(n1782), .IN2(n19642), .IN3(n1678), .IN4(n19629), .Q(
        n7263) );
  OA22X1 U26151 ( .IN1(n1954), .IN2(n19677), .IN3(n1868), .IN4(n19661), .Q(
        n7264) );
  OA22X1 U26152 ( .IN1(n2126), .IN2(n19710), .IN3(n2040), .IN4(n19694), .Q(
        n7265) );
  NAND4X0 U26153 ( .IN1(n7259), .IN2(n7260), .IN3(n7261), .IN4(n7262), .QN(
        s15_addr_o[8]) );
  OA22X1 U26154 ( .IN1(n1781), .IN2(n19642), .IN3(n1677), .IN4(n19628), .Q(
        n7259) );
  OA22X1 U26155 ( .IN1(n1953), .IN2(n19672), .IN3(n1867), .IN4(n19661), .Q(
        n7260) );
  OA22X1 U26156 ( .IN1(n2125), .IN2(n19705), .IN3(n2039), .IN4(n19694), .Q(
        n7261) );
  NAND4X0 U26157 ( .IN1(n7255), .IN2(n7256), .IN3(n7257), .IN4(n7258), .QN(
        s15_addr_o[9]) );
  OA22X1 U26158 ( .IN1(n1780), .IN2(n19642), .IN3(n1676), .IN4(n19628), .Q(
        n7255) );
  OA22X1 U26159 ( .IN1(n1952), .IN2(n19675), .IN3(n1866), .IN4(n19662), .Q(
        n7256) );
  OA22X1 U26160 ( .IN1(n2124), .IN2(n19708), .IN3(n2038), .IN4(n19695), .Q(
        n7257) );
  NAND4X0 U26161 ( .IN1(n7343), .IN2(n7344), .IN3(n7345), .IN4(n7346), .QN(
        s15_addr_o[10]) );
  OA22X1 U26162 ( .IN1(n1779), .IN2(n19639), .IN3(n1675), .IN4(n19623), .Q(
        n7343) );
  OA22X1 U26163 ( .IN1(n1951), .IN2(n19675), .IN3(n1865), .IN4(n19658), .Q(
        n7344) );
  OA22X1 U26164 ( .IN1(n2123), .IN2(n19708), .IN3(n2037), .IN4(n19691), .Q(
        n7345) );
  NAND4X0 U26165 ( .IN1(n7339), .IN2(n7340), .IN3(n7341), .IN4(n7342), .QN(
        s15_addr_o[11]) );
  OA22X1 U26166 ( .IN1(n1778), .IN2(n19643), .IN3(n1674), .IN4(n19624), .Q(
        n7339) );
  OA22X1 U26167 ( .IN1(n1950), .IN2(n19676), .IN3(n1864), .IN4(n19659), .Q(
        n7340) );
  OA22X1 U26168 ( .IN1(n2122), .IN2(n19709), .IN3(n2036), .IN4(n19692), .Q(
        n7341) );
  NAND4X0 U26169 ( .IN1(n7335), .IN2(n7336), .IN3(n7337), .IN4(n7338), .QN(
        s15_addr_o[12]) );
  OA22X1 U26170 ( .IN1(n1777), .IN2(n19640), .IN3(n1673), .IN4(n19624), .Q(
        n7335) );
  OA22X1 U26171 ( .IN1(n1949), .IN2(n19674), .IN3(n1863), .IN4(n19659), .Q(
        n7336) );
  OA22X1 U26172 ( .IN1(n2121), .IN2(n19707), .IN3(n2035), .IN4(n19692), .Q(
        n7337) );
  NAND4X0 U26173 ( .IN1(n7331), .IN2(n7332), .IN3(n7333), .IN4(n7334), .QN(
        s15_addr_o[13]) );
  OA22X1 U26174 ( .IN1(n1776), .IN2(n19640), .IN3(n1672), .IN4(n19624), .Q(
        n7331) );
  OA22X1 U26175 ( .IN1(n1948), .IN2(n19674), .IN3(n1862), .IN4(n19659), .Q(
        n7332) );
  OA22X1 U26176 ( .IN1(n2120), .IN2(n19707), .IN3(n2034), .IN4(n19692), .Q(
        n7333) );
  NAND4X0 U26177 ( .IN1(n7327), .IN2(n7328), .IN3(n7329), .IN4(n7330), .QN(
        s15_addr_o[14]) );
  OA22X1 U26178 ( .IN1(n1775), .IN2(n19640), .IN3(n1671), .IN4(n19631), .Q(
        n7327) );
  OA22X1 U26179 ( .IN1(n1947), .IN2(n19674), .IN3(n1861), .IN4(n19660), .Q(
        n7328) );
  OA22X1 U26180 ( .IN1(n2119), .IN2(n19707), .IN3(n2033), .IN4(n19693), .Q(
        n7329) );
  NAND4X0 U26181 ( .IN1(n7323), .IN2(n7324), .IN3(n7325), .IN4(n7326), .QN(
        s15_addr_o[15]) );
  OA22X1 U26182 ( .IN1(n1774), .IN2(n19640), .IN3(n1670), .IN4(n19631), .Q(
        n7323) );
  OA22X1 U26183 ( .IN1(n1946), .IN2(n19674), .IN3(n1860), .IN4(n19660), .Q(
        n7324) );
  OA22X1 U26184 ( .IN1(n2118), .IN2(n19707), .IN3(n2032), .IN4(n19693), .Q(
        n7325) );
  NAND4X0 U26185 ( .IN1(n7319), .IN2(n7320), .IN3(n7321), .IN4(n7322), .QN(
        s15_addr_o[16]) );
  OA22X1 U26186 ( .IN1(n1773), .IN2(n19641), .IN3(n1669), .IN4(n19631), .Q(
        n7319) );
  OA22X1 U26187 ( .IN1(n1945), .IN2(n19676), .IN3(n1859), .IN4(n19660), .Q(
        n7320) );
  OA22X1 U26188 ( .IN1(n2117), .IN2(n19709), .IN3(n2031), .IN4(n19693), .Q(
        n7321) );
  NAND4X0 U26189 ( .IN1(n7315), .IN2(n7316), .IN3(n7317), .IN4(n7318), .QN(
        s15_addr_o[17]) );
  OA22X1 U26190 ( .IN1(n1772), .IN2(n19641), .IN3(n1668), .IN4(n19625), .Q(
        n7315) );
  OA22X1 U26191 ( .IN1(n1944), .IN2(n19673), .IN3(n1858), .IN4(n19660), .Q(
        n7316) );
  OA22X1 U26192 ( .IN1(n2116), .IN2(n19706), .IN3(n2030), .IN4(n19693), .Q(
        n7317) );
  NAND4X0 U26193 ( .IN1(n7311), .IN2(n7312), .IN3(n7313), .IN4(n7314), .QN(
        s15_addr_o[18]) );
  OA22X1 U26194 ( .IN1(n1771), .IN2(n19641), .IN3(n1667), .IN4(n19625), .Q(
        n7311) );
  OA22X1 U26195 ( .IN1(n1943), .IN2(n19675), .IN3(n1857), .IN4(n19660), .Q(
        n7312) );
  OA22X1 U26196 ( .IN1(n2115), .IN2(n19708), .IN3(n2029), .IN4(n19693), .Q(
        n7313) );
  NAND4X0 U26197 ( .IN1(n7307), .IN2(n7308), .IN3(n7309), .IN4(n7310), .QN(
        s15_addr_o[19]) );
  OA22X1 U26198 ( .IN1(n1770), .IN2(n19641), .IN3(n1666), .IN4(n19625), .Q(
        n7307) );
  OA22X1 U26199 ( .IN1(n1942), .IN2(n19674), .IN3(n1856), .IN4(n19663), .Q(
        n7308) );
  OA22X1 U26200 ( .IN1(n2114), .IN2(n19707), .IN3(n2028), .IN4(n19696), .Q(
        n7309) );
  NAND4X0 U26201 ( .IN1(n7299), .IN2(n7300), .IN3(n7301), .IN4(n7302), .QN(
        s15_addr_o[20]) );
  OA22X1 U26202 ( .IN1(n1769), .IN2(n19642), .IN3(n1665), .IN4(n19626), .Q(
        n7299) );
  OA22X1 U26203 ( .IN1(n1941), .IN2(n19674), .IN3(n1855), .IN4(n19656), .Q(
        n7300) );
  OA22X1 U26204 ( .IN1(n2113), .IN2(n19707), .IN3(n2027), .IN4(n19689), .Q(
        n7301) );
  NAND4X0 U26205 ( .IN1(n7295), .IN2(n7296), .IN3(n7297), .IN4(n7298), .QN(
        s15_addr_o[21]) );
  OA22X1 U26206 ( .IN1(n1768), .IN2(n19642), .IN3(n1664), .IN4(n19626), .Q(
        n7295) );
  OA22X1 U26207 ( .IN1(n1940), .IN2(n19675), .IN3(n1854), .IN4(n19656), .Q(
        n7296) );
  OA22X1 U26208 ( .IN1(n2112), .IN2(n19708), .IN3(n2026), .IN4(n19689), .Q(
        n7297) );
  NAND4X0 U26209 ( .IN1(n7291), .IN2(n7292), .IN3(n7293), .IN4(n7294), .QN(
        s15_addr_o[22]) );
  OA22X1 U26210 ( .IN1(n1767), .IN2(n19642), .IN3(n1663), .IN4(n19627), .Q(
        n7291) );
  OA22X1 U26211 ( .IN1(n1939), .IN2(n19677), .IN3(n1853), .IN4(n19655), .Q(
        n7292) );
  OA22X1 U26212 ( .IN1(n2111), .IN2(n19710), .IN3(n2025), .IN4(n19688), .Q(
        n7293) );
  NAND4X0 U26213 ( .IN1(n7287), .IN2(n7288), .IN3(n7289), .IN4(n7290), .QN(
        s15_addr_o[23]) );
  OA22X1 U26214 ( .IN1(n1766), .IN2(n19643), .IN3(n1662), .IN4(n19627), .Q(
        n7287) );
  OA22X1 U26215 ( .IN1(n1938), .IN2(n19676), .IN3(n1852), .IN4(n19655), .Q(
        n7288) );
  OA22X1 U26216 ( .IN1(n2110), .IN2(n19709), .IN3(n2024), .IN4(n19688), .Q(
        n7289) );
  NAND4X0 U26217 ( .IN1(n7283), .IN2(n7284), .IN3(n7285), .IN4(n7286), .QN(
        s15_addr_o[28]) );
  OA22X1 U26218 ( .IN1(n1761), .IN2(n19643), .IN3(n1657), .IN4(n19627), .Q(
        n7283) );
  OA22X1 U26219 ( .IN1(n1933), .IN2(n19674), .IN3(n1847), .IN4(n19655), .Q(
        n7284) );
  OA22X1 U26220 ( .IN1(n2105), .IN2(n19707), .IN3(n2019), .IN4(n19688), .Q(
        n7285) );
  NAND4X0 U26221 ( .IN1(n7279), .IN2(n7280), .IN3(n7281), .IN4(n7282), .QN(
        s15_addr_o[29]) );
  OA22X1 U26222 ( .IN1(n1760), .IN2(n19643), .IN3(n1656), .IN4(n19626), .Q(
        n7279) );
  OA22X1 U26223 ( .IN1(n1932), .IN2(n19674), .IN3(n1846), .IN4(n19656), .Q(
        n7280) );
  OA22X1 U26224 ( .IN1(n2104), .IN2(n19707), .IN3(n2018), .IN4(n19689), .Q(
        n7281) );
  NAND4X0 U26225 ( .IN1(n7275), .IN2(n7276), .IN3(n7277), .IN4(n7278), .QN(
        s15_addr_o[30]) );
  OA22X1 U26226 ( .IN1(n1759), .IN2(n19643), .IN3(n1655), .IN4(n19627), .Q(
        n7275) );
  OA22X1 U26227 ( .IN1(n1931), .IN2(n19675), .IN3(n1845), .IN4(n19655), .Q(
        n7276) );
  OA22X1 U26228 ( .IN1(n2103), .IN2(n19708), .IN3(n2017), .IN4(n19688), .Q(
        n7277) );
  NAND4X0 U26229 ( .IN1(n7271), .IN2(n7272), .IN3(n7273), .IN4(n7274), .QN(
        s15_addr_o[31]) );
  OA22X1 U26230 ( .IN1(n1758), .IN2(n19643), .IN3(n1650), .IN4(n19630), .Q(
        n7271) );
  OA22X1 U26231 ( .IN1(n1930), .IN2(n19677), .IN3(n1844), .IN4(n19658), .Q(
        n7272) );
  OA22X1 U26232 ( .IN1(n2102), .IN2(n19710), .IN3(n2016), .IN4(n19691), .Q(
        n7273) );
  NAND4X0 U26233 ( .IN1(n7251), .IN2(n7252), .IN3(n7253), .IN4(n7254), .QN(
        s15_data_o[16]) );
  OA22X1 U26234 ( .IN1(n1725), .IN2(n19641), .IN3(n1620), .IN4(n19628), .Q(
        n7251) );
  OA22X1 U26235 ( .IN1(n1897), .IN2(n19675), .IN3(n1811), .IN4(n19662), .Q(
        n7252) );
  OA22X1 U26236 ( .IN1(n2069), .IN2(n19708), .IN3(n1983), .IN4(n19695), .Q(
        n7253) );
  NAND4X0 U26237 ( .IN1(n7247), .IN2(n7248), .IN3(n7249), .IN4(n7250), .QN(
        s15_data_o[17]) );
  OA22X1 U26238 ( .IN1(n1724), .IN2(n19643), .IN3(n1619), .IN4(n19628), .Q(
        n7247) );
  OA22X1 U26239 ( .IN1(n1896), .IN2(n19675), .IN3(n1810), .IN4(n19662), .Q(
        n7248) );
  OA22X1 U26240 ( .IN1(n2068), .IN2(n19708), .IN3(n1982), .IN4(n19695), .Q(
        n7249) );
  NAND4X0 U26241 ( .IN1(n7243), .IN2(n7244), .IN3(n7245), .IN4(n7246), .QN(
        s15_data_o[18]) );
  OA22X1 U26242 ( .IN1(n1723), .IN2(n19640), .IN3(n1618), .IN4(n19628), .Q(
        n7243) );
  OA22X1 U26243 ( .IN1(n1895), .IN2(n19675), .IN3(n1809), .IN4(n19657), .Q(
        n7244) );
  OA22X1 U26244 ( .IN1(n2067), .IN2(n19708), .IN3(n1981), .IN4(n19690), .Q(
        n7245) );
  NAND4X0 U26245 ( .IN1(n7239), .IN2(n7240), .IN3(n7241), .IN4(n7242), .QN(
        s15_data_o[19]) );
  OA22X1 U26246 ( .IN1(n1722), .IN2(n19639), .IN3(n1617), .IN4(n19628), .Q(
        n7239) );
  OA22X1 U26247 ( .IN1(n1894), .IN2(n19676), .IN3(n1808), .IN4(n19661), .Q(
        n7240) );
  OA22X1 U26248 ( .IN1(n2066), .IN2(n19709), .IN3(n1980), .IN4(n19694), .Q(
        n7241) );
  NAND4X0 U26249 ( .IN1(n7235), .IN2(n7236), .IN3(n7237), .IN4(n7238), .QN(
        s15_data_o[20]) );
  OA22X1 U26250 ( .IN1(n1721), .IN2(n19644), .IN3(n1616), .IN4(n19629), .Q(
        n7235) );
  OA22X1 U26251 ( .IN1(n1893), .IN2(n19676), .IN3(n1807), .IN4(n19662), .Q(
        n7236) );
  OA22X1 U26252 ( .IN1(n2065), .IN2(n19709), .IN3(n1979), .IN4(n19695), .Q(
        n7237) );
  NAND4X0 U26253 ( .IN1(n7231), .IN2(n7232), .IN3(n7233), .IN4(n7234), .QN(
        s15_data_o[21]) );
  OA22X1 U26254 ( .IN1(n1720), .IN2(n19641), .IN3(n1615), .IN4(n19629), .Q(
        n7231) );
  OA22X1 U26255 ( .IN1(n1892), .IN2(n19676), .IN3(n1806), .IN4(n19663), .Q(
        n7232) );
  OA22X1 U26256 ( .IN1(n2064), .IN2(n19709), .IN3(n1978), .IN4(n19696), .Q(
        n7233) );
  NAND4X0 U26257 ( .IN1(n7227), .IN2(n7228), .IN3(n7229), .IN4(n7230), .QN(
        s15_data_o[22]) );
  OA22X1 U26258 ( .IN1(n1719), .IN2(n19640), .IN3(n1614), .IN4(n19629), .Q(
        n7227) );
  OA22X1 U26259 ( .IN1(n1891), .IN2(n19676), .IN3(n1805), .IN4(n19663), .Q(
        n7228) );
  OA22X1 U26260 ( .IN1(n2063), .IN2(n19709), .IN3(n1977), .IN4(n19696), .Q(
        n7229) );
  NAND4X0 U26261 ( .IN1(n7223), .IN2(n7224), .IN3(n7225), .IN4(n7226), .QN(
        s15_data_o[23]) );
  OA22X1 U26262 ( .IN1(n1718), .IN2(n19639), .IN3(n1613), .IN4(n19629), .Q(
        n7223) );
  OA22X1 U26263 ( .IN1(n1890), .IN2(n19674), .IN3(n1804), .IN4(n19663), .Q(
        n7224) );
  OA22X1 U26264 ( .IN1(n2062), .IN2(n19707), .IN3(n1976), .IN4(n19696), .Q(
        n7225) );
  NAND4X0 U26265 ( .IN1(n7219), .IN2(n7220), .IN3(n7221), .IN4(n7222), .QN(
        s15_data_o[24]) );
  OA22X1 U26266 ( .IN1(n1717), .IN2(n19644), .IN3(n1612), .IN4(n19630), .Q(
        n7219) );
  OA22X1 U26267 ( .IN1(n1889), .IN2(n19675), .IN3(n1803), .IN4(n19659), .Q(
        n7220) );
  OA22X1 U26268 ( .IN1(n2061), .IN2(n19708), .IN3(n1975), .IN4(n19692), .Q(
        n7221) );
  NAND4X0 U26269 ( .IN1(n7215), .IN2(n7216), .IN3(n7217), .IN4(n7218), .QN(
        s15_data_o[25]) );
  OA22X1 U26270 ( .IN1(n1716), .IN2(n19639), .IN3(n1611), .IN4(n19630), .Q(
        n7215) );
  OA22X1 U26271 ( .IN1(n1888), .IN2(n19676), .IN3(n1802), .IN4(n19661), .Q(
        n7216) );
  OA22X1 U26272 ( .IN1(n2060), .IN2(n19709), .IN3(n1974), .IN4(n19694), .Q(
        n7217) );
  NAND4X0 U26273 ( .IN1(n7211), .IN2(n7212), .IN3(n7213), .IN4(n7214), .QN(
        s15_data_o[26]) );
  OA22X1 U26274 ( .IN1(n1715), .IN2(n19644), .IN3(n1610), .IN4(n19630), .Q(
        n7211) );
  OA22X1 U26275 ( .IN1(n1887), .IN2(n19672), .IN3(n1801), .IN4(n19662), .Q(
        n7212) );
  OA22X1 U26276 ( .IN1(n2059), .IN2(n19705), .IN3(n1973), .IN4(n19695), .Q(
        n7213) );
  NAND4X0 U26277 ( .IN1(n7207), .IN2(n7208), .IN3(n7209), .IN4(n7210), .QN(
        s15_data_o[27]) );
  OA22X1 U26278 ( .IN1(n1714), .IN2(n19644), .IN3(n1609), .IN4(n19622), .Q(
        n7207) );
  OA22X1 U26279 ( .IN1(n1886), .IN2(n19677), .IN3(n1800), .IN4(n19656), .Q(
        n7208) );
  OA22X1 U26280 ( .IN1(n2058), .IN2(n19710), .IN3(n1972), .IN4(n19689), .Q(
        n7209) );
  NAND4X0 U26281 ( .IN1(n7203), .IN2(n7204), .IN3(n7205), .IN4(n7206), .QN(
        s15_data_o[28]) );
  OA22X1 U26282 ( .IN1(n1713), .IN2(n19644), .IN3(n1608), .IN4(n19631), .Q(
        n7203) );
  OA22X1 U26283 ( .IN1(n1885), .IN2(n19677), .IN3(n1799), .IN4(n19664), .Q(
        n7204) );
  OA22X1 U26284 ( .IN1(n2057), .IN2(n19710), .IN3(n1971), .IN4(n19697), .Q(
        n7205) );
  NAND4X0 U26285 ( .IN1(n7199), .IN2(n7200), .IN3(n7201), .IN4(n7202), .QN(
        s15_data_o[29]) );
  OA22X1 U26286 ( .IN1(n1712), .IN2(n19644), .IN3(n1607), .IN4(n19622), .Q(
        n7199) );
  OA22X1 U26287 ( .IN1(n1884), .IN2(n19677), .IN3(n1798), .IN4(n19656), .Q(
        n7200) );
  OA22X1 U26288 ( .IN1(n2056), .IN2(n19710), .IN3(n1970), .IN4(n19689), .Q(
        n7201) );
  NAND4X0 U26289 ( .IN1(n7195), .IN2(n7196), .IN3(n7197), .IN4(n7198), .QN(
        s15_data_o[30]) );
  OA22X1 U26290 ( .IN1(n1711), .IN2(n19644), .IN3(n1606), .IN4(n19631), .Q(
        n7195) );
  OA22X1 U26291 ( .IN1(n1883), .IN2(n19677), .IN3(n1797), .IN4(n19664), .Q(
        n7196) );
  OA22X1 U26292 ( .IN1(n2055), .IN2(n19710), .IN3(n1969), .IN4(n19697), .Q(
        n7197) );
  NAND4X0 U26293 ( .IN1(n7191), .IN2(n7192), .IN3(n7193), .IN4(n7194), .QN(
        s15_data_o[31]) );
  OA22X1 U26294 ( .IN1(n1710), .IN2(n19639), .IN3(n1605), .IN4(n19624), .Q(
        n7191) );
  OA22X1 U26295 ( .IN1(n1882), .IN2(n19676), .IN3(n1796), .IN4(n19656), .Q(
        n7192) );
  OA22X1 U26296 ( .IN1(n2054), .IN2(n19709), .IN3(n1968), .IN4(n19689), .Q(
        n7193) );
  NAND4X0 U26297 ( .IN1(n7363), .IN2(n7364), .IN3(n7365), .IN4(n7366), .QN(
        s14_stb_o) );
  OA22X1 U26298 ( .IN1(n1795), .IN2(n7373), .IN3(n1709), .IN4(n7374), .Q(n7363) );
  OA22X1 U26299 ( .IN1(n1967), .IN2(n7371), .IN3(n1881), .IN4(n7372), .Q(n7364) );
  OA22X1 U26300 ( .IN1(n2139), .IN2(n7369), .IN3(n2053), .IN4(n7370), .Q(n7365) );
  NAND4X0 U26301 ( .IN1(n7351), .IN2(n7352), .IN3(n7353), .IN4(n7354), .QN(
        s14_we_o) );
  OA22X1 U26302 ( .IN1(n1794), .IN2(n19505), .IN3(n1708), .IN4(n19499), .Q(
        n7351) );
  OA22X1 U26303 ( .IN1(n1966), .IN2(n19538), .IN3(n1880), .IN4(n19532), .Q(
        n7352) );
  OA22X1 U26304 ( .IN1(n2138), .IN2(n19571), .IN3(n2052), .IN4(n19566), .Q(
        n7353) );
  NAND4X0 U26305 ( .IN1(n7387), .IN2(n7388), .IN3(n7389), .IN4(n7390), .QN(
        s14_sel_o[0]) );
  OA22X1 U26306 ( .IN1(n1793), .IN2(n19512), .IN3(n1707), .IN4(n19498), .Q(
        n7387) );
  OA22X1 U26307 ( .IN1(n1965), .IN2(n19545), .IN3(n1879), .IN4(n19531), .Q(
        n7388) );
  OA22X1 U26308 ( .IN1(n2137), .IN2(n19578), .IN3(n2051), .IN4(n19565), .Q(
        n7389) );
  NAND4X0 U26309 ( .IN1(n7383), .IN2(n7384), .IN3(n7385), .IN4(n7386), .QN(
        s14_sel_o[1]) );
  OA22X1 U26310 ( .IN1(n1792), .IN2(n19512), .IN3(n1706), .IN4(n19498), .Q(
        n7383) );
  OA22X1 U26311 ( .IN1(n1964), .IN2(n19545), .IN3(n1878), .IN4(n19531), .Q(
        n7384) );
  OA22X1 U26312 ( .IN1(n2136), .IN2(n19578), .IN3(n2050), .IN4(n19565), .Q(
        n7385) );
  NAND4X0 U26313 ( .IN1(n7379), .IN2(n7380), .IN3(n7381), .IN4(n7382), .QN(
        s14_sel_o[2]) );
  OA22X1 U26314 ( .IN1(n1791), .IN2(n19512), .IN3(n1705), .IN4(n19499), .Q(
        n7379) );
  OA22X1 U26315 ( .IN1(n1963), .IN2(n19545), .IN3(n1877), .IN4(n19532), .Q(
        n7380) );
  OA22X1 U26316 ( .IN1(n2135), .IN2(n19578), .IN3(n2049), .IN4(n19566), .Q(
        n7381) );
  NAND4X0 U26317 ( .IN1(n7375), .IN2(n7376), .IN3(n7377), .IN4(n7378), .QN(
        s14_sel_o[3]) );
  OA22X1 U26318 ( .IN1(n1790), .IN2(n19512), .IN3(n1704), .IN4(n19499), .Q(
        n7375) );
  OA22X1 U26319 ( .IN1(n1962), .IN2(n19545), .IN3(n1876), .IN4(n19532), .Q(
        n7376) );
  OA22X1 U26320 ( .IN1(n2134), .IN2(n19578), .IN3(n2048), .IN4(n19566), .Q(
        n7377) );
  NAND4X0 U26321 ( .IN1(n7643), .IN2(n7644), .IN3(n7645), .IN4(n7646), .QN(
        s14_addr_o[0]) );
  OA22X1 U26322 ( .IN1(n1789), .IN2(n19505), .IN3(n1703), .IN4(n19482), .Q(
        n7643) );
  OA22X1 U26323 ( .IN1(n1961), .IN2(n19538), .IN3(n1875), .IN4(n19515), .Q(
        n7644) );
  OA22X1 U26324 ( .IN1(n2133), .IN2(n19571), .IN3(n2047), .IN4(n19548), .Q(
        n7645) );
  NAND4X0 U26325 ( .IN1(n7599), .IN2(n7600), .IN3(n7601), .IN4(n7602), .QN(
        s14_addr_o[1]) );
  OA22X1 U26326 ( .IN1(n1788), .IN2(n19507), .IN3(n1702), .IN4(n19485), .Q(
        n7599) );
  OA22X1 U26327 ( .IN1(n1960), .IN2(n19540), .IN3(n1874), .IN4(n19518), .Q(
        n7600) );
  OA22X1 U26328 ( .IN1(n2132), .IN2(n19573), .IN3(n2046), .IN4(n19551), .Q(
        n7601) );
  NAND4X0 U26329 ( .IN1(n7555), .IN2(n7556), .IN3(n7557), .IN4(n7558), .QN(
        s14_addr_o[2]) );
  OA22X1 U26330 ( .IN1(n1787), .IN2(n19507), .IN3(n1701), .IN4(n19489), .Q(
        n7555) );
  OA22X1 U26331 ( .IN1(n1959), .IN2(n19540), .IN3(n1873), .IN4(n19522), .Q(
        n7556) );
  OA22X1 U26332 ( .IN1(n2131), .IN2(n19573), .IN3(n2045), .IN4(n19555), .Q(
        n7557) );
  NAND4X0 U26333 ( .IN1(n7543), .IN2(n7544), .IN3(n7545), .IN4(n7546), .QN(
        s14_addr_o[3]) );
  OA22X1 U26334 ( .IN1(n1786), .IN2(n19512), .IN3(n1699), .IN4(n19490), .Q(
        n7543) );
  OA22X1 U26335 ( .IN1(n1958), .IN2(n19545), .IN3(n1872), .IN4(n19523), .Q(
        n7544) );
  OA22X1 U26336 ( .IN1(n2130), .IN2(n19578), .IN3(n2044), .IN4(n19562), .Q(
        n7545) );
  NAND4X0 U26337 ( .IN1(n7539), .IN2(n7540), .IN3(n7541), .IN4(n7542), .QN(
        s14_addr_o[4]) );
  OA22X1 U26338 ( .IN1(n1785), .IN2(n19505), .IN3(n1697), .IN4(n19490), .Q(
        n7539) );
  OA22X1 U26339 ( .IN1(n1957), .IN2(n19538), .IN3(n1871), .IN4(n19523), .Q(
        n7540) );
  OA22X1 U26340 ( .IN1(n2129), .IN2(n19571), .IN3(n2043), .IN4(n19564), .Q(
        n7541) );
  NAND4X0 U26341 ( .IN1(n7535), .IN2(n7536), .IN3(n7537), .IN4(n7538), .QN(
        s14_addr_o[5]) );
  OA22X1 U26342 ( .IN1(n1784), .IN2(n19512), .IN3(n1696), .IN4(n19489), .Q(
        n7535) );
  OA22X1 U26343 ( .IN1(n1956), .IN2(n19545), .IN3(n1870), .IN4(n19522), .Q(
        n7536) );
  OA22X1 U26344 ( .IN1(n2128), .IN2(n19578), .IN3(n2042), .IN4(n19556), .Q(
        n7537) );
  NAND4X0 U26345 ( .IN1(n7531), .IN2(n7532), .IN3(n7533), .IN4(n7534), .QN(
        s14_addr_o[6]) );
  OA22X1 U26346 ( .IN1(n1783), .IN2(n19508), .IN3(n1679), .IN4(n19490), .Q(
        n7531) );
  OA22X1 U26347 ( .IN1(n1955), .IN2(n19541), .IN3(n1869), .IN4(n19523), .Q(
        n7532) );
  OA22X1 U26348 ( .IN1(n2127), .IN2(n19574), .IN3(n2041), .IN4(n19556), .Q(
        n7533) );
  NAND4X0 U26349 ( .IN1(n7527), .IN2(n7528), .IN3(n7529), .IN4(n7530), .QN(
        s14_addr_o[7]) );
  OA22X1 U26350 ( .IN1(n1782), .IN2(n19508), .IN3(n1678), .IN4(n19482), .Q(
        n7527) );
  OA22X1 U26351 ( .IN1(n1954), .IN2(n19541), .IN3(n1868), .IN4(n19515), .Q(
        n7528) );
  OA22X1 U26352 ( .IN1(n2126), .IN2(n19574), .IN3(n2040), .IN4(n19556), .Q(
        n7529) );
  NAND4X0 U26353 ( .IN1(n7523), .IN2(n7524), .IN3(n7525), .IN4(n7526), .QN(
        s14_addr_o[8]) );
  OA22X1 U26354 ( .IN1(n1781), .IN2(n19508), .IN3(n1677), .IN4(n19491), .Q(
        n7523) );
  OA22X1 U26355 ( .IN1(n1953), .IN2(n19541), .IN3(n1867), .IN4(n19524), .Q(
        n7524) );
  OA22X1 U26356 ( .IN1(n2125), .IN2(n19574), .IN3(n2039), .IN4(n19557), .Q(
        n7525) );
  NAND4X0 U26357 ( .IN1(n7519), .IN2(n7520), .IN3(n7521), .IN4(n7522), .QN(
        s14_addr_o[9]) );
  OA22X1 U26358 ( .IN1(n1780), .IN2(n19508), .IN3(n1676), .IN4(n19491), .Q(
        n7519) );
  OA22X1 U26359 ( .IN1(n1952), .IN2(n19541), .IN3(n1866), .IN4(n19524), .Q(
        n7520) );
  OA22X1 U26360 ( .IN1(n2124), .IN2(n19574), .IN3(n2038), .IN4(n19557), .Q(
        n7521) );
  NAND4X0 U26361 ( .IN1(n7639), .IN2(n7640), .IN3(n7641), .IN4(n7642), .QN(
        s14_addr_o[10]) );
  OA22X1 U26362 ( .IN1(n1779), .IN2(n19505), .IN3(n1675), .IN4(n19482), .Q(
        n7639) );
  OA22X1 U26363 ( .IN1(n1951), .IN2(n19538), .IN3(n1865), .IN4(n19515), .Q(
        n7640) );
  OA22X1 U26364 ( .IN1(n2123), .IN2(n19571), .IN3(n2037), .IN4(n19548), .Q(
        n7641) );
  NAND4X0 U26365 ( .IN1(n7635), .IN2(n7636), .IN3(n7637), .IN4(n7638), .QN(
        s14_addr_o[11]) );
  OA22X1 U26366 ( .IN1(n1778), .IN2(n19505), .IN3(n1674), .IN4(n19482), .Q(
        n7635) );
  OA22X1 U26367 ( .IN1(n1950), .IN2(n19538), .IN3(n1864), .IN4(n19515), .Q(
        n7636) );
  OA22X1 U26368 ( .IN1(n2122), .IN2(n19571), .IN3(n2036), .IN4(n19548), .Q(
        n7637) );
  NAND4X0 U26369 ( .IN1(n7631), .IN2(n7632), .IN3(n7633), .IN4(n7634), .QN(
        s14_addr_o[12]) );
  OA22X1 U26370 ( .IN1(n1777), .IN2(n19505), .IN3(n1673), .IN4(n19483), .Q(
        n7631) );
  OA22X1 U26371 ( .IN1(n1949), .IN2(n19538), .IN3(n1863), .IN4(n19516), .Q(
        n7632) );
  OA22X1 U26372 ( .IN1(n2121), .IN2(n19571), .IN3(n2035), .IN4(n19549), .Q(
        n7633) );
  NAND4X0 U26373 ( .IN1(n7627), .IN2(n7628), .IN3(n7629), .IN4(n7630), .QN(
        s14_addr_o[13]) );
  OA22X1 U26374 ( .IN1(n1776), .IN2(n19506), .IN3(n1672), .IN4(n19483), .Q(
        n7627) );
  OA22X1 U26375 ( .IN1(n1948), .IN2(n19539), .IN3(n1862), .IN4(n19516), .Q(
        n7628) );
  OA22X1 U26376 ( .IN1(n2120), .IN2(n19572), .IN3(n2034), .IN4(n19549), .Q(
        n7629) );
  NAND4X0 U26377 ( .IN1(n7623), .IN2(n7624), .IN3(n7625), .IN4(n7626), .QN(
        s14_addr_o[14]) );
  OA22X1 U26378 ( .IN1(n1775), .IN2(n19506), .IN3(n1671), .IN4(n19483), .Q(
        n7623) );
  OA22X1 U26379 ( .IN1(n1947), .IN2(n19539), .IN3(n1861), .IN4(n19516), .Q(
        n7624) );
  OA22X1 U26380 ( .IN1(n2119), .IN2(n19572), .IN3(n2033), .IN4(n19549), .Q(
        n7625) );
  NAND4X0 U26381 ( .IN1(n7619), .IN2(n7620), .IN3(n7621), .IN4(n7622), .QN(
        s14_addr_o[15]) );
  OA22X1 U26382 ( .IN1(n1774), .IN2(n19506), .IN3(n1670), .IN4(n19484), .Q(
        n7619) );
  OA22X1 U26383 ( .IN1(n1946), .IN2(n19539), .IN3(n1860), .IN4(n19517), .Q(
        n7620) );
  OA22X1 U26384 ( .IN1(n2118), .IN2(n19572), .IN3(n2032), .IN4(n19550), .Q(
        n7621) );
  NAND4X0 U26385 ( .IN1(n7615), .IN2(n7616), .IN3(n7617), .IN4(n7618), .QN(
        s14_addr_o[16]) );
  OA22X1 U26386 ( .IN1(n1773), .IN2(n19506), .IN3(n1669), .IN4(n19484), .Q(
        n7615) );
  OA22X1 U26387 ( .IN1(n1945), .IN2(n19539), .IN3(n1859), .IN4(n19517), .Q(
        n7616) );
  OA22X1 U26388 ( .IN1(n2117), .IN2(n19572), .IN3(n2031), .IN4(n19550), .Q(
        n7617) );
  NAND4X0 U26389 ( .IN1(n7611), .IN2(n7612), .IN3(n7613), .IN4(n7614), .QN(
        s14_addr_o[17]) );
  OA22X1 U26390 ( .IN1(n1772), .IN2(n19507), .IN3(n1668), .IN4(n19484), .Q(
        n7611) );
  OA22X1 U26391 ( .IN1(n1944), .IN2(n19540), .IN3(n1858), .IN4(n19517), .Q(
        n7612) );
  OA22X1 U26392 ( .IN1(n2116), .IN2(n19573), .IN3(n2030), .IN4(n19550), .Q(
        n7613) );
  NAND4X0 U26393 ( .IN1(n7607), .IN2(n7608), .IN3(n7609), .IN4(n7610), .QN(
        s14_addr_o[18]) );
  OA22X1 U26394 ( .IN1(n1771), .IN2(n19507), .IN3(n1667), .IN4(n19485), .Q(
        n7607) );
  OA22X1 U26395 ( .IN1(n1943), .IN2(n19540), .IN3(n1857), .IN4(n19518), .Q(
        n7608) );
  OA22X1 U26396 ( .IN1(n2115), .IN2(n19573), .IN3(n2029), .IN4(n19551), .Q(
        n7609) );
  NAND4X0 U26397 ( .IN1(n7603), .IN2(n7604), .IN3(n7605), .IN4(n7606), .QN(
        s14_addr_o[19]) );
  OA22X1 U26398 ( .IN1(n1770), .IN2(n19507), .IN3(n1666), .IN4(n19485), .Q(
        n7603) );
  OA22X1 U26399 ( .IN1(n1942), .IN2(n19540), .IN3(n1856), .IN4(n19518), .Q(
        n7604) );
  OA22X1 U26400 ( .IN1(n2114), .IN2(n19573), .IN3(n2028), .IN4(n19551), .Q(
        n7605) );
  NAND4X0 U26401 ( .IN1(n7595), .IN2(n7596), .IN3(n7597), .IN4(n7598), .QN(
        s14_addr_o[20]) );
  OA22X1 U26402 ( .IN1(n1769), .IN2(n19506), .IN3(n1665), .IN4(n19486), .Q(
        n7595) );
  OA22X1 U26403 ( .IN1(n1941), .IN2(n19539), .IN3(n1855), .IN4(n19519), .Q(
        n7596) );
  OA22X1 U26404 ( .IN1(n2113), .IN2(n19572), .IN3(n2027), .IN4(n19552), .Q(
        n7597) );
  NAND4X0 U26405 ( .IN1(n7591), .IN2(n7592), .IN3(n7593), .IN4(n7594), .QN(
        s14_addr_o[21]) );
  OA22X1 U26406 ( .IN1(n1768), .IN2(n19506), .IN3(n1664), .IN4(n19486), .Q(
        n7591) );
  OA22X1 U26407 ( .IN1(n1940), .IN2(n19539), .IN3(n1854), .IN4(n19519), .Q(
        n7592) );
  OA22X1 U26408 ( .IN1(n2112), .IN2(n19572), .IN3(n2026), .IN4(n19552), .Q(
        n7593) );
  NAND4X0 U26409 ( .IN1(n7587), .IN2(n7588), .IN3(n7589), .IN4(n7590), .QN(
        s14_addr_o[22]) );
  OA22X1 U26410 ( .IN1(n1767), .IN2(n19505), .IN3(n1663), .IN4(n19486), .Q(
        n7587) );
  OA22X1 U26411 ( .IN1(n1939), .IN2(n19538), .IN3(n1853), .IN4(n19519), .Q(
        n7588) );
  OA22X1 U26412 ( .IN1(n2111), .IN2(n19571), .IN3(n2025), .IN4(n19552), .Q(
        n7589) );
  NAND4X0 U26413 ( .IN1(n7583), .IN2(n7584), .IN3(n7585), .IN4(n7586), .QN(
        s14_addr_o[23]) );
  OA22X1 U26414 ( .IN1(n1766), .IN2(n19506), .IN3(n1662), .IN4(n19487), .Q(
        n7583) );
  OA22X1 U26415 ( .IN1(n1938), .IN2(n19539), .IN3(n1852), .IN4(n19520), .Q(
        n7584) );
  OA22X1 U26416 ( .IN1(n2110), .IN2(n19572), .IN3(n2024), .IN4(n19553), .Q(
        n7585) );
  NAND4X0 U26417 ( .IN1(n7579), .IN2(n7580), .IN3(n7581), .IN4(n7582), .QN(
        s14_addr_o[24]) );
  OA22X1 U26418 ( .IN1(n1765), .IN2(n19512), .IN3(n1661), .IN4(n19487), .Q(
        n7579) );
  OA22X1 U26419 ( .IN1(n1937), .IN2(n19545), .IN3(n1851), .IN4(n19520), .Q(
        n7580) );
  OA22X1 U26420 ( .IN1(n2109), .IN2(n19578), .IN3(n2023), .IN4(n19553), .Q(
        n7581) );
  NAND4X0 U26421 ( .IN1(n7575), .IN2(n7576), .IN3(n7577), .IN4(n7578), .QN(
        s14_addr_o[25]) );
  OA22X1 U26422 ( .IN1(n1764), .IN2(n19508), .IN3(n1660), .IN4(n19487), .Q(
        n7575) );
  OA22X1 U26423 ( .IN1(n1936), .IN2(n19541), .IN3(n1850), .IN4(n19520), .Q(
        n7576) );
  OA22X1 U26424 ( .IN1(n2108), .IN2(n19574), .IN3(n2022), .IN4(n19553), .Q(
        n7577) );
  NAND4X0 U26425 ( .IN1(n7571), .IN2(n7572), .IN3(n7573), .IN4(n7574), .QN(
        s14_addr_o[26]) );
  OA22X1 U26426 ( .IN1(n1763), .IN2(n19507), .IN3(n1659), .IN4(n19488), .Q(
        n7571) );
  OA22X1 U26427 ( .IN1(n1935), .IN2(n19540), .IN3(n1849), .IN4(n19521), .Q(
        n7572) );
  OA22X1 U26428 ( .IN1(n2107), .IN2(n19573), .IN3(n2021), .IN4(n19554), .Q(
        n7573) );
  NAND4X0 U26429 ( .IN1(n7567), .IN2(n7568), .IN3(n7569), .IN4(n7570), .QN(
        s14_addr_o[27]) );
  OA22X1 U26430 ( .IN1(n1762), .IN2(n19506), .IN3(n1658), .IN4(n19488), .Q(
        n7567) );
  OA22X1 U26431 ( .IN1(n1934), .IN2(n19539), .IN3(n1848), .IN4(n19521), .Q(
        n7568) );
  OA22X1 U26432 ( .IN1(n2106), .IN2(n19572), .IN3(n2020), .IN4(n19554), .Q(
        n7569) );
  NAND4X0 U26433 ( .IN1(n7563), .IN2(n7564), .IN3(n7565), .IN4(n7566), .QN(
        s14_addr_o[28]) );
  OA22X1 U26434 ( .IN1(n1761), .IN2(n19506), .IN3(n1657), .IN4(n19488), .Q(
        n7563) );
  OA22X1 U26435 ( .IN1(n1933), .IN2(n19539), .IN3(n1847), .IN4(n19521), .Q(
        n7564) );
  OA22X1 U26436 ( .IN1(n2105), .IN2(n19572), .IN3(n2019), .IN4(n19554), .Q(
        n7565) );
  NAND4X0 U26437 ( .IN1(n7559), .IN2(n7560), .IN3(n7561), .IN4(n7562), .QN(
        s14_addr_o[29]) );
  OA22X1 U26438 ( .IN1(n1760), .IN2(n19510), .IN3(n1656), .IN4(n19489), .Q(
        n7559) );
  OA22X1 U26439 ( .IN1(n1932), .IN2(n19543), .IN3(n1846), .IN4(n19522), .Q(
        n7560) );
  OA22X1 U26440 ( .IN1(n2104), .IN2(n19577), .IN3(n2018), .IN4(n19555), .Q(
        n7561) );
  NAND4X0 U26441 ( .IN1(n7551), .IN2(n7552), .IN3(n7553), .IN4(n7554), .QN(
        s14_addr_o[30]) );
  OA22X1 U26442 ( .IN1(n1759), .IN2(n19511), .IN3(n1655), .IN4(n19489), .Q(
        n7551) );
  OA22X1 U26443 ( .IN1(n1931), .IN2(n19544), .IN3(n1845), .IN4(n19522), .Q(
        n7552) );
  OA22X1 U26444 ( .IN1(n2103), .IN2(n19575), .IN3(n2017), .IN4(n19555), .Q(
        n7553) );
  NAND4X0 U26445 ( .IN1(n7547), .IN2(n7548), .IN3(n7549), .IN4(n7550), .QN(
        s14_addr_o[31]) );
  OA22X1 U26446 ( .IN1(n1758), .IN2(n19509), .IN3(n1650), .IN4(n19490), .Q(
        n7547) );
  OA22X1 U26447 ( .IN1(n1930), .IN2(n19542), .IN3(n1844), .IN4(n19523), .Q(
        n7548) );
  OA22X1 U26448 ( .IN1(n2102), .IN2(n19576), .IN3(n2016), .IN4(n19562), .Q(
        n7549) );
  NAND4X0 U26449 ( .IN1(n7515), .IN2(n7516), .IN3(n7517), .IN4(n7518), .QN(
        s14_data_o[0]) );
  OA22X1 U26450 ( .IN1(n1741), .IN2(n19508), .IN3(n1636), .IN4(n19491), .Q(
        n7515) );
  OA22X1 U26451 ( .IN1(n1913), .IN2(n19541), .IN3(n1827), .IN4(n19524), .Q(
        n7516) );
  OA22X1 U26452 ( .IN1(n2085), .IN2(n19574), .IN3(n1999), .IN4(n19557), .Q(
        n7517) );
  NAND4X0 U26453 ( .IN1(n7471), .IN2(n7472), .IN3(n7473), .IN4(n7474), .QN(
        s14_data_o[1]) );
  OA22X1 U26454 ( .IN1(n1740), .IN2(n19510), .IN3(n1635), .IN4(n19489), .Q(
        n7471) );
  OA22X1 U26455 ( .IN1(n1912), .IN2(n19543), .IN3(n1826), .IN4(n19522), .Q(
        n7472) );
  OA22X1 U26456 ( .IN1(n2084), .IN2(n19576), .IN3(n1998), .IN4(n19560), .Q(
        n7473) );
  NAND4X0 U26457 ( .IN1(n7427), .IN2(n7428), .IN3(n7429), .IN4(n7430), .QN(
        s14_data_o[2]) );
  OA22X1 U26458 ( .IN1(n1739), .IN2(n19511), .IN3(n1634), .IN4(n19482), .Q(
        n7427) );
  OA22X1 U26459 ( .IN1(n1911), .IN2(n19544), .IN3(n1825), .IN4(n19515), .Q(
        n7428) );
  OA22X1 U26460 ( .IN1(n2083), .IN2(n19576), .IN3(n1997), .IN4(n19564), .Q(
        n7429) );
  NAND4X0 U26461 ( .IN1(n7415), .IN2(n7416), .IN3(n7417), .IN4(n7418), .QN(
        s14_data_o[3]) );
  OA22X1 U26462 ( .IN1(n1738), .IN2(n19509), .IN3(n1633), .IN4(n19484), .Q(
        n7415) );
  OA22X1 U26463 ( .IN1(n1910), .IN2(n19542), .IN3(n1824), .IN4(n19517), .Q(
        n7416) );
  OA22X1 U26464 ( .IN1(n2082), .IN2(n19575), .IN3(n1996), .IN4(n19563), .Q(
        n7417) );
  NAND4X0 U26465 ( .IN1(n7411), .IN2(n7412), .IN3(n7413), .IN4(n7414), .QN(
        s14_data_o[4]) );
  OA22X1 U26466 ( .IN1(n1737), .IN2(n19510), .IN3(n1632), .IN4(n19499), .Q(
        n7411) );
  OA22X1 U26467 ( .IN1(n1909), .IN2(n19543), .IN3(n1823), .IN4(n19532), .Q(
        n7412) );
  OA22X1 U26468 ( .IN1(n2081), .IN2(n19575), .IN3(n1995), .IN4(n19563), .Q(
        n7413) );
  NAND4X0 U26469 ( .IN1(n7407), .IN2(n7408), .IN3(n7409), .IN4(n7410), .QN(
        s14_data_o[5]) );
  OA22X1 U26470 ( .IN1(n1736), .IN2(n19511), .IN3(n1631), .IN4(n19497), .Q(
        n7407) );
  OA22X1 U26471 ( .IN1(n1908), .IN2(n19544), .IN3(n1822), .IN4(n19530), .Q(
        n7408) );
  OA22X1 U26472 ( .IN1(n2080), .IN2(n19576), .IN3(n1994), .IN4(n19563), .Q(
        n7409) );
  NAND4X0 U26473 ( .IN1(n7403), .IN2(n7404), .IN3(n7405), .IN4(n7406), .QN(
        s14_data_o[6]) );
  OA22X1 U26474 ( .IN1(n1735), .IN2(n19507), .IN3(n1630), .IN4(n19497), .Q(
        n7403) );
  OA22X1 U26475 ( .IN1(n1907), .IN2(n19540), .IN3(n1821), .IN4(n19530), .Q(
        n7404) );
  OA22X1 U26476 ( .IN1(n2079), .IN2(n19573), .IN3(n1993), .IN4(n19564), .Q(
        n7405) );
  NAND4X0 U26477 ( .IN1(n7399), .IN2(n7400), .IN3(n7401), .IN4(n7402), .QN(
        s14_data_o[7]) );
  OA22X1 U26478 ( .IN1(n1734), .IN2(n19505), .IN3(n1629), .IN4(n19497), .Q(
        n7399) );
  OA22X1 U26479 ( .IN1(n1906), .IN2(n19538), .IN3(n1820), .IN4(n19530), .Q(
        n7400) );
  OA22X1 U26480 ( .IN1(n2078), .IN2(n19571), .IN3(n1992), .IN4(n19564), .Q(
        n7401) );
  NAND4X0 U26481 ( .IN1(n7395), .IN2(n7396), .IN3(n7397), .IN4(n7398), .QN(
        s14_data_o[8]) );
  OA22X1 U26482 ( .IN1(n1733), .IN2(n19512), .IN3(n1628), .IN4(n19497), .Q(
        n7395) );
  OA22X1 U26483 ( .IN1(n1905), .IN2(n19545), .IN3(n1819), .IN4(n19530), .Q(
        n7396) );
  OA22X1 U26484 ( .IN1(n2077), .IN2(n19578), .IN3(n1991), .IN4(n19564), .Q(
        n7397) );
  NAND4X0 U26485 ( .IN1(n7391), .IN2(n7392), .IN3(n7393), .IN4(n7394), .QN(
        s14_data_o[9]) );
  OA22X1 U26486 ( .IN1(n1732), .IN2(n19505), .IN3(n1627), .IN4(n19498), .Q(
        n7391) );
  OA22X1 U26487 ( .IN1(n1904), .IN2(n19538), .IN3(n1818), .IN4(n19531), .Q(
        n7392) );
  OA22X1 U26488 ( .IN1(n2076), .IN2(n19571), .IN3(n1990), .IN4(n19565), .Q(
        n7393) );
  NAND4X0 U26489 ( .IN1(n7511), .IN2(n7512), .IN3(n7513), .IN4(n7514), .QN(
        s14_data_o[10]) );
  OA22X1 U26490 ( .IN1(n1731), .IN2(n19507), .IN3(n1626), .IN4(n19492), .Q(
        n7511) );
  OA22X1 U26491 ( .IN1(n1903), .IN2(n19540), .IN3(n1817), .IN4(n19525), .Q(
        n7512) );
  OA22X1 U26492 ( .IN1(n2075), .IN2(n19573), .IN3(n1989), .IN4(n19558), .Q(
        n7513) );
  NAND4X0 U26493 ( .IN1(n7507), .IN2(n7508), .IN3(n7509), .IN4(n7510), .QN(
        s14_data_o[11]) );
  OA22X1 U26494 ( .IN1(n1730), .IN2(n19512), .IN3(n1625), .IN4(n19492), .Q(
        n7507) );
  OA22X1 U26495 ( .IN1(n1902), .IN2(n19545), .IN3(n1816), .IN4(n19525), .Q(
        n7508) );
  OA22X1 U26496 ( .IN1(n2074), .IN2(n19578), .IN3(n1988), .IN4(n19558), .Q(
        n7509) );
  NAND4X0 U26497 ( .IN1(n7503), .IN2(n7504), .IN3(n7505), .IN4(n7506), .QN(
        s14_data_o[12]) );
  OA22X1 U26498 ( .IN1(n1729), .IN2(n19508), .IN3(n1624), .IN4(n19492), .Q(
        n7503) );
  OA22X1 U26499 ( .IN1(n1901), .IN2(n19541), .IN3(n1815), .IN4(n19525), .Q(
        n7504) );
  OA22X1 U26500 ( .IN1(n2073), .IN2(n19574), .IN3(n1987), .IN4(n19558), .Q(
        n7505) );
  NAND4X0 U26501 ( .IN1(n7499), .IN2(n7500), .IN3(n7501), .IN4(n7502), .QN(
        s14_data_o[13]) );
  OA22X1 U26502 ( .IN1(n1728), .IN2(n19509), .IN3(n1623), .IN4(n19486), .Q(
        n7499) );
  OA22X1 U26503 ( .IN1(n1900), .IN2(n19542), .IN3(n1814), .IN4(n19519), .Q(
        n7500) );
  OA22X1 U26504 ( .IN1(n2072), .IN2(n19575), .IN3(n1986), .IN4(n19559), .Q(
        n7501) );
  NAND4X0 U26505 ( .IN1(n7495), .IN2(n7496), .IN3(n7497), .IN4(n7498), .QN(
        s14_data_o[14]) );
  OA22X1 U26506 ( .IN1(n1727), .IN2(n19509), .IN3(n1622), .IN4(n19491), .Q(
        n7495) );
  OA22X1 U26507 ( .IN1(n1899), .IN2(n19542), .IN3(n1813), .IN4(n19524), .Q(
        n7496) );
  OA22X1 U26508 ( .IN1(n2071), .IN2(n19575), .IN3(n1985), .IN4(n19559), .Q(
        n7497) );
  NAND4X0 U26509 ( .IN1(n7491), .IN2(n7492), .IN3(n7493), .IN4(n7494), .QN(
        s14_data_o[15]) );
  OA22X1 U26510 ( .IN1(n1726), .IN2(n19509), .IN3(n1621), .IN4(n19492), .Q(
        n7491) );
  OA22X1 U26511 ( .IN1(n1898), .IN2(n19542), .IN3(n1812), .IN4(n19525), .Q(
        n7492) );
  OA22X1 U26512 ( .IN1(n2070), .IN2(n19575), .IN3(n1984), .IN4(n19559), .Q(
        n7493) );
  NAND4X0 U26513 ( .IN1(n7487), .IN2(n7488), .IN3(n7489), .IN4(n7490), .QN(
        s14_data_o[16]) );
  OA22X1 U26514 ( .IN1(n1725), .IN2(n19509), .IN3(n1620), .IN4(n19493), .Q(
        n7487) );
  OA22X1 U26515 ( .IN1(n1897), .IN2(n19542), .IN3(n1811), .IN4(n19526), .Q(
        n7488) );
  OA22X1 U26516 ( .IN1(n2069), .IN2(n19575), .IN3(n1983), .IN4(n19548), .Q(
        n7489) );
  NAND4X0 U26517 ( .IN1(n7483), .IN2(n7484), .IN3(n7485), .IN4(n7486), .QN(
        s14_data_o[17]) );
  OA22X1 U26518 ( .IN1(n1724), .IN2(n19510), .IN3(n1619), .IN4(n19493), .Q(
        n7483) );
  OA22X1 U26519 ( .IN1(n1896), .IN2(n19543), .IN3(n1810), .IN4(n19526), .Q(
        n7484) );
  OA22X1 U26520 ( .IN1(n2068), .IN2(n19576), .IN3(n1982), .IN4(n19549), .Q(
        n7485) );
  NAND4X0 U26521 ( .IN1(n7479), .IN2(n7480), .IN3(n7481), .IN4(n7482), .QN(
        s14_data_o[18]) );
  OA22X1 U26522 ( .IN1(n1723), .IN2(n19510), .IN3(n1618), .IN4(n19493), .Q(
        n7479) );
  OA22X1 U26523 ( .IN1(n1895), .IN2(n19543), .IN3(n1809), .IN4(n19526), .Q(
        n7480) );
  OA22X1 U26524 ( .IN1(n2067), .IN2(n19576), .IN3(n1981), .IN4(n19550), .Q(
        n7481) );
  NAND4X0 U26525 ( .IN1(n7475), .IN2(n7476), .IN3(n7477), .IN4(n7478), .QN(
        s14_data_o[19]) );
  OA22X1 U26526 ( .IN1(n1722), .IN2(n19510), .IN3(n1617), .IN4(n19493), .Q(
        n7475) );
  OA22X1 U26527 ( .IN1(n1894), .IN2(n19543), .IN3(n1808), .IN4(n19526), .Q(
        n7476) );
  OA22X1 U26528 ( .IN1(n2066), .IN2(n19576), .IN3(n1980), .IN4(n19561), .Q(
        n7477) );
  NAND4X0 U26529 ( .IN1(n7467), .IN2(n7468), .IN3(n7469), .IN4(n7470), .QN(
        s14_data_o[20]) );
  OA22X1 U26530 ( .IN1(n1721), .IN2(n19511), .IN3(n1616), .IN4(n19490), .Q(
        n7467) );
  OA22X1 U26531 ( .IN1(n1893), .IN2(n19544), .IN3(n1807), .IN4(n19523), .Q(
        n7468) );
  OA22X1 U26532 ( .IN1(n2065), .IN2(n19577), .IN3(n1979), .IN4(n19566), .Q(
        n7469) );
  NAND4X0 U26533 ( .IN1(n7463), .IN2(n7464), .IN3(n7465), .IN4(n7466), .QN(
        s14_data_o[21]) );
  OA22X1 U26534 ( .IN1(n1720), .IN2(n19511), .IN3(n1615), .IN4(n19494), .Q(
        n7463) );
  OA22X1 U26535 ( .IN1(n1892), .IN2(n19544), .IN3(n1806), .IN4(n19527), .Q(
        n7464) );
  OA22X1 U26536 ( .IN1(n2064), .IN2(n19577), .IN3(n1978), .IN4(n19560), .Q(
        n7465) );
  NAND4X0 U26537 ( .IN1(n7459), .IN2(n7460), .IN3(n7461), .IN4(n7462), .QN(
        s14_data_o[22]) );
  OA22X1 U26538 ( .IN1(n1719), .IN2(n19509), .IN3(n1614), .IN4(n19494), .Q(
        n7459) );
  OA22X1 U26539 ( .IN1(n1891), .IN2(n19542), .IN3(n1805), .IN4(n19527), .Q(
        n7460) );
  OA22X1 U26540 ( .IN1(n2063), .IN2(n19577), .IN3(n1977), .IN4(n19560), .Q(
        n7461) );
  NAND4X0 U26541 ( .IN1(n7455), .IN2(n7456), .IN3(n7457), .IN4(n7458), .QN(
        s14_data_o[23]) );
  OA22X1 U26542 ( .IN1(n1718), .IN2(n19510), .IN3(n1613), .IN4(n19494), .Q(
        n7455) );
  OA22X1 U26543 ( .IN1(n1890), .IN2(n19543), .IN3(n1804), .IN4(n19527), .Q(
        n7456) );
  OA22X1 U26544 ( .IN1(n2062), .IN2(n19577), .IN3(n1976), .IN4(n19560), .Q(
        n7457) );
  NAND4X0 U26545 ( .IN1(n7451), .IN2(n7452), .IN3(n7453), .IN4(n7454), .QN(
        s14_data_o[24]) );
  OA22X1 U26546 ( .IN1(n1717), .IN2(n19508), .IN3(n1612), .IN4(n19495), .Q(
        n7451) );
  OA22X1 U26547 ( .IN1(n1889), .IN2(n19541), .IN3(n1803), .IN4(n19528), .Q(
        n7452) );
  OA22X1 U26548 ( .IN1(n2061), .IN2(n19574), .IN3(n1975), .IN4(n19561), .Q(
        n7453) );
  NAND4X0 U26549 ( .IN1(n7447), .IN2(n7448), .IN3(n7449), .IN4(n7450), .QN(
        s14_data_o[25]) );
  OA22X1 U26550 ( .IN1(n1716), .IN2(n19508), .IN3(n1611), .IN4(n19495), .Q(
        n7447) );
  OA22X1 U26551 ( .IN1(n1888), .IN2(n19541), .IN3(n1802), .IN4(n19528), .Q(
        n7448) );
  OA22X1 U26552 ( .IN1(n2060), .IN2(n19574), .IN3(n1974), .IN4(n19561), .Q(
        n7449) );
  NAND4X0 U26553 ( .IN1(n7443), .IN2(n7444), .IN3(n7445), .IN4(n7446), .QN(
        s14_data_o[26]) );
  OA22X1 U26554 ( .IN1(n1715), .IN2(n19507), .IN3(n1610), .IN4(n19495), .Q(
        n7443) );
  OA22X1 U26555 ( .IN1(n1887), .IN2(n19540), .IN3(n1801), .IN4(n19528), .Q(
        n7444) );
  OA22X1 U26556 ( .IN1(n2059), .IN2(n19573), .IN3(n1973), .IN4(n19561), .Q(
        n7445) );
  NAND4X0 U26557 ( .IN1(n7439), .IN2(n7440), .IN3(n7441), .IN4(n7442), .QN(
        s14_data_o[27]) );
  OA22X1 U26558 ( .IN1(n1714), .IN2(n19510), .IN3(n1609), .IN4(n19496), .Q(
        n7439) );
  OA22X1 U26559 ( .IN1(n1886), .IN2(n19543), .IN3(n1800), .IN4(n19529), .Q(
        n7440) );
  OA22X1 U26560 ( .IN1(n2058), .IN2(n19577), .IN3(n1972), .IN4(n19562), .Q(
        n7441) );
  NAND4X0 U26561 ( .IN1(n7435), .IN2(n7436), .IN3(n7437), .IN4(n7438), .QN(
        s14_data_o[28]) );
  OA22X1 U26562 ( .IN1(n1713), .IN2(n19511), .IN3(n1608), .IN4(n19496), .Q(
        n7435) );
  OA22X1 U26563 ( .IN1(n1885), .IN2(n19544), .IN3(n1799), .IN4(n19529), .Q(
        n7436) );
  OA22X1 U26564 ( .IN1(n2057), .IN2(n19577), .IN3(n1971), .IN4(n19562), .Q(
        n7437) );
  NAND4X0 U26565 ( .IN1(n7431), .IN2(n7432), .IN3(n7433), .IN4(n7434), .QN(
        s14_data_o[29]) );
  OA22X1 U26566 ( .IN1(n1712), .IN2(n19511), .IN3(n1607), .IN4(n19496), .Q(
        n7431) );
  OA22X1 U26567 ( .IN1(n1884), .IN2(n19544), .IN3(n1798), .IN4(n19529), .Q(
        n7432) );
  OA22X1 U26568 ( .IN1(n2056), .IN2(n19575), .IN3(n1970), .IN4(n19562), .Q(
        n7433) );
  NAND4X0 U26569 ( .IN1(n7423), .IN2(n7424), .IN3(n7425), .IN4(n7426), .QN(
        s14_data_o[30]) );
  OA22X1 U26570 ( .IN1(n1711), .IN2(n19511), .IN3(n1606), .IN4(n19498), .Q(
        n7423) );
  OA22X1 U26571 ( .IN1(n1883), .IN2(n19544), .IN3(n1797), .IN4(n19531), .Q(
        n7424) );
  OA22X1 U26572 ( .IN1(n2055), .IN2(n19576), .IN3(n1969), .IN4(n19560), .Q(
        n7425) );
  NAND4X0 U26573 ( .IN1(n7419), .IN2(n7420), .IN3(n7421), .IN4(n7422), .QN(
        s14_data_o[31]) );
  OA22X1 U26574 ( .IN1(n1710), .IN2(n19509), .IN3(n1605), .IN4(n19483), .Q(
        n7419) );
  OA22X1 U26575 ( .IN1(n1882), .IN2(n19542), .IN3(n1796), .IN4(n19516), .Q(
        n7420) );
  OA22X1 U26576 ( .IN1(n2054), .IN2(n19577), .IN3(n1968), .IN4(n19561), .Q(
        n7421) );
  NAND4X0 U26577 ( .IN1(n7659), .IN2(n7660), .IN3(n7661), .IN4(n7662), .QN(
        s13_stb_o) );
  OA22X1 U26578 ( .IN1(n1795), .IN2(n7669), .IN3(n1709), .IN4(n7670), .Q(n7659) );
  OA22X1 U26579 ( .IN1(n1967), .IN2(n7667), .IN3(n1881), .IN4(n7668), .Q(n7660) );
  OA22X1 U26580 ( .IN1(n2139), .IN2(n7665), .IN3(n2053), .IN4(n7666), .Q(n7661) );
  NAND4X0 U26581 ( .IN1(n7647), .IN2(n7648), .IN3(n7649), .IN4(n7650), .QN(
        s13_we_o) );
  OA22X1 U26582 ( .IN1(n1794), .IN2(n19373), .IN3(n1708), .IN4(n19367), .Q(
        n7647) );
  OA22X1 U26583 ( .IN1(n1966), .IN2(n19406), .IN3(n1880), .IN4(n19400), .Q(
        n7648) );
  OA22X1 U26584 ( .IN1(n2138), .IN2(n19439), .IN3(n2052), .IN4(n19433), .Q(
        n7649) );
  NAND4X0 U26585 ( .IN1(n7683), .IN2(n7684), .IN3(n7685), .IN4(n7686), .QN(
        s13_sel_o[0]) );
  OA22X1 U26586 ( .IN1(n1793), .IN2(n19380), .IN3(n1707), .IN4(n19366), .Q(
        n7683) );
  OA22X1 U26587 ( .IN1(n1965), .IN2(n19413), .IN3(n1879), .IN4(n19399), .Q(
        n7684) );
  OA22X1 U26588 ( .IN1(n2137), .IN2(n19446), .IN3(n2051), .IN4(n19432), .Q(
        n7685) );
  NAND4X0 U26589 ( .IN1(n7679), .IN2(n7680), .IN3(n7681), .IN4(n7682), .QN(
        s13_sel_o[1]) );
  OA22X1 U26590 ( .IN1(n1792), .IN2(n19380), .IN3(n1706), .IN4(n19366), .Q(
        n7679) );
  OA22X1 U26591 ( .IN1(n1964), .IN2(n19413), .IN3(n1878), .IN4(n19399), .Q(
        n7680) );
  OA22X1 U26592 ( .IN1(n2136), .IN2(n19446), .IN3(n2050), .IN4(n19432), .Q(
        n7681) );
  NAND4X0 U26593 ( .IN1(n7675), .IN2(n7676), .IN3(n7677), .IN4(n7678), .QN(
        s13_sel_o[2]) );
  OA22X1 U26594 ( .IN1(n1791), .IN2(n19380), .IN3(n1705), .IN4(n19367), .Q(
        n7675) );
  OA22X1 U26595 ( .IN1(n1963), .IN2(n19413), .IN3(n1877), .IN4(n19400), .Q(
        n7676) );
  OA22X1 U26596 ( .IN1(n2135), .IN2(n19446), .IN3(n2049), .IN4(n19433), .Q(
        n7677) );
  NAND4X0 U26597 ( .IN1(n7671), .IN2(n7672), .IN3(n7673), .IN4(n7674), .QN(
        s13_sel_o[3]) );
  OA22X1 U26598 ( .IN1(n1790), .IN2(n19380), .IN3(n1704), .IN4(n19367), .Q(
        n7671) );
  OA22X1 U26599 ( .IN1(n1962), .IN2(n19413), .IN3(n1876), .IN4(n19400), .Q(
        n7672) );
  OA22X1 U26600 ( .IN1(n2134), .IN2(n19446), .IN3(n2048), .IN4(n19433), .Q(
        n7673) );
  NAND4X0 U26601 ( .IN1(n7939), .IN2(n7940), .IN3(n7941), .IN4(n7942), .QN(
        s13_addr_o[0]) );
  OA22X1 U26602 ( .IN1(n1789), .IN2(n19373), .IN3(n1703), .IN4(n19350), .Q(
        n7939) );
  OA22X1 U26603 ( .IN1(n1961), .IN2(n19406), .IN3(n1875), .IN4(n19383), .Q(
        n7940) );
  OA22X1 U26604 ( .IN1(n2133), .IN2(n19439), .IN3(n2047), .IN4(n19416), .Q(
        n7941) );
  NAND4X0 U26605 ( .IN1(n7895), .IN2(n7896), .IN3(n7897), .IN4(n7898), .QN(
        s13_addr_o[1]) );
  OA22X1 U26606 ( .IN1(n1788), .IN2(n19375), .IN3(n1702), .IN4(n19353), .Q(
        n7895) );
  OA22X1 U26607 ( .IN1(n1960), .IN2(n19408), .IN3(n1874), .IN4(n19386), .Q(
        n7896) );
  OA22X1 U26608 ( .IN1(n2132), .IN2(n19441), .IN3(n2046), .IN4(n19419), .Q(
        n7897) );
  NAND4X0 U26609 ( .IN1(n7851), .IN2(n7852), .IN3(n7853), .IN4(n7854), .QN(
        s13_addr_o[2]) );
  OA22X1 U26610 ( .IN1(n1787), .IN2(n19375), .IN3(n1701), .IN4(n19357), .Q(
        n7851) );
  OA22X1 U26611 ( .IN1(n1959), .IN2(n19408), .IN3(n1873), .IN4(n19390), .Q(
        n7852) );
  OA22X1 U26612 ( .IN1(n2131), .IN2(n19441), .IN3(n2045), .IN4(n19423), .Q(
        n7853) );
  NAND4X0 U26613 ( .IN1(n7839), .IN2(n7840), .IN3(n7841), .IN4(n7842), .QN(
        s13_addr_o[3]) );
  OA22X1 U26614 ( .IN1(n1786), .IN2(n19380), .IN3(n1699), .IN4(n19358), .Q(
        n7839) );
  OA22X1 U26615 ( .IN1(n1958), .IN2(n19413), .IN3(n1872), .IN4(n19391), .Q(
        n7840) );
  OA22X1 U26616 ( .IN1(n2130), .IN2(n19446), .IN3(n2044), .IN4(n19424), .Q(
        n7841) );
  NAND4X0 U26617 ( .IN1(n7835), .IN2(n7836), .IN3(n7837), .IN4(n7838), .QN(
        s13_addr_o[4]) );
  OA22X1 U26618 ( .IN1(n1785), .IN2(n19373), .IN3(n1697), .IN4(n19358), .Q(
        n7835) );
  OA22X1 U26619 ( .IN1(n1957), .IN2(n19406), .IN3(n1871), .IN4(n19391), .Q(
        n7836) );
  OA22X1 U26620 ( .IN1(n2129), .IN2(n19439), .IN3(n2043), .IN4(n19424), .Q(
        n7837) );
  NAND4X0 U26621 ( .IN1(n7831), .IN2(n7832), .IN3(n7833), .IN4(n7834), .QN(
        s13_addr_o[5]) );
  OA22X1 U26622 ( .IN1(n1784), .IN2(n19380), .IN3(n1696), .IN4(n19357), .Q(
        n7831) );
  OA22X1 U26623 ( .IN1(n1956), .IN2(n19413), .IN3(n1870), .IN4(n19390), .Q(
        n7832) );
  OA22X1 U26624 ( .IN1(n2128), .IN2(n19446), .IN3(n2042), .IN4(n19423), .Q(
        n7833) );
  NAND4X0 U26625 ( .IN1(n7827), .IN2(n7828), .IN3(n7829), .IN4(n7830), .QN(
        s13_addr_o[6]) );
  OA22X1 U26626 ( .IN1(n1783), .IN2(n19376), .IN3(n1679), .IN4(n19358), .Q(
        n7827) );
  OA22X1 U26627 ( .IN1(n1955), .IN2(n19409), .IN3(n1869), .IN4(n19391), .Q(
        n7828) );
  OA22X1 U26628 ( .IN1(n2127), .IN2(n19442), .IN3(n2041), .IN4(n19424), .Q(
        n7829) );
  NAND4X0 U26629 ( .IN1(n7823), .IN2(n7824), .IN3(n7825), .IN4(n7826), .QN(
        s13_addr_o[7]) );
  OA22X1 U26630 ( .IN1(n1782), .IN2(n19376), .IN3(n1678), .IN4(n19350), .Q(
        n7823) );
  OA22X1 U26631 ( .IN1(n1954), .IN2(n19409), .IN3(n1868), .IN4(n19383), .Q(
        n7824) );
  OA22X1 U26632 ( .IN1(n2126), .IN2(n19442), .IN3(n2040), .IN4(n19423), .Q(
        n7825) );
  NAND4X0 U26633 ( .IN1(n7819), .IN2(n7820), .IN3(n7821), .IN4(n7822), .QN(
        s13_addr_o[8]) );
  OA22X1 U26634 ( .IN1(n1781), .IN2(n19376), .IN3(n1677), .IN4(n19359), .Q(
        n7819) );
  OA22X1 U26635 ( .IN1(n1953), .IN2(n19409), .IN3(n1867), .IN4(n19392), .Q(
        n7820) );
  OA22X1 U26636 ( .IN1(n2125), .IN2(n19442), .IN3(n2039), .IN4(n19425), .Q(
        n7821) );
  NAND4X0 U26637 ( .IN1(n7815), .IN2(n7816), .IN3(n7817), .IN4(n7818), .QN(
        s13_addr_o[9]) );
  OA22X1 U26638 ( .IN1(n1780), .IN2(n19376), .IN3(n1676), .IN4(n19359), .Q(
        n7815) );
  OA22X1 U26639 ( .IN1(n1952), .IN2(n19409), .IN3(n1866), .IN4(n19392), .Q(
        n7816) );
  OA22X1 U26640 ( .IN1(n2124), .IN2(n19442), .IN3(n2038), .IN4(n19425), .Q(
        n7817) );
  NAND4X0 U26641 ( .IN1(n7935), .IN2(n7936), .IN3(n7937), .IN4(n7938), .QN(
        s13_addr_o[10]) );
  OA22X1 U26642 ( .IN1(n1779), .IN2(n19373), .IN3(n1675), .IN4(n19350), .Q(
        n7935) );
  OA22X1 U26643 ( .IN1(n1951), .IN2(n19406), .IN3(n1865), .IN4(n19383), .Q(
        n7936) );
  OA22X1 U26644 ( .IN1(n2123), .IN2(n19439), .IN3(n2037), .IN4(n19416), .Q(
        n7937) );
  NAND4X0 U26645 ( .IN1(n7931), .IN2(n7932), .IN3(n7933), .IN4(n7934), .QN(
        s13_addr_o[11]) );
  OA22X1 U26646 ( .IN1(n1778), .IN2(n19373), .IN3(n1674), .IN4(n19350), .Q(
        n7931) );
  OA22X1 U26647 ( .IN1(n1950), .IN2(n19406), .IN3(n1864), .IN4(n19383), .Q(
        n7932) );
  OA22X1 U26648 ( .IN1(n2122), .IN2(n19439), .IN3(n2036), .IN4(n19416), .Q(
        n7933) );
  NAND4X0 U26649 ( .IN1(n7927), .IN2(n7928), .IN3(n7929), .IN4(n7930), .QN(
        s13_addr_o[12]) );
  OA22X1 U26650 ( .IN1(n1777), .IN2(n19373), .IN3(n1673), .IN4(n19351), .Q(
        n7927) );
  OA22X1 U26651 ( .IN1(n1949), .IN2(n19406), .IN3(n1863), .IN4(n19384), .Q(
        n7928) );
  OA22X1 U26652 ( .IN1(n2121), .IN2(n19439), .IN3(n2035), .IN4(n19417), .Q(
        n7929) );
  NAND4X0 U26653 ( .IN1(n7923), .IN2(n7924), .IN3(n7925), .IN4(n7926), .QN(
        s13_addr_o[13]) );
  OA22X1 U26654 ( .IN1(n1776), .IN2(n19374), .IN3(n1672), .IN4(n19351), .Q(
        n7923) );
  OA22X1 U26655 ( .IN1(n1948), .IN2(n19407), .IN3(n1862), .IN4(n19384), .Q(
        n7924) );
  OA22X1 U26656 ( .IN1(n2120), .IN2(n19440), .IN3(n2034), .IN4(n19417), .Q(
        n7925) );
  NAND4X0 U26657 ( .IN1(n7919), .IN2(n7920), .IN3(n7921), .IN4(n7922), .QN(
        s13_addr_o[14]) );
  OA22X1 U26658 ( .IN1(n1775), .IN2(n19374), .IN3(n1671), .IN4(n19351), .Q(
        n7919) );
  OA22X1 U26659 ( .IN1(n1947), .IN2(n19407), .IN3(n1861), .IN4(n19384), .Q(
        n7920) );
  OA22X1 U26660 ( .IN1(n2119), .IN2(n19440), .IN3(n2033), .IN4(n19417), .Q(
        n7921) );
  NAND4X0 U26661 ( .IN1(n7915), .IN2(n7916), .IN3(n7917), .IN4(n7918), .QN(
        s13_addr_o[15]) );
  OA22X1 U26662 ( .IN1(n1774), .IN2(n19374), .IN3(n1670), .IN4(n19352), .Q(
        n7915) );
  OA22X1 U26663 ( .IN1(n1946), .IN2(n19407), .IN3(n1860), .IN4(n19385), .Q(
        n7916) );
  OA22X1 U26664 ( .IN1(n2118), .IN2(n19440), .IN3(n2032), .IN4(n19418), .Q(
        n7917) );
  NAND4X0 U26665 ( .IN1(n7911), .IN2(n7912), .IN3(n7913), .IN4(n7914), .QN(
        s13_addr_o[16]) );
  OA22X1 U26666 ( .IN1(n1773), .IN2(n19374), .IN3(n1669), .IN4(n19352), .Q(
        n7911) );
  OA22X1 U26667 ( .IN1(n1945), .IN2(n19407), .IN3(n1859), .IN4(n19385), .Q(
        n7912) );
  OA22X1 U26668 ( .IN1(n2117), .IN2(n19440), .IN3(n2031), .IN4(n19418), .Q(
        n7913) );
  NAND4X0 U26669 ( .IN1(n7907), .IN2(n7908), .IN3(n7909), .IN4(n7910), .QN(
        s13_addr_o[17]) );
  OA22X1 U26670 ( .IN1(n1772), .IN2(n19375), .IN3(n1668), .IN4(n19352), .Q(
        n7907) );
  OA22X1 U26671 ( .IN1(n1944), .IN2(n19408), .IN3(n1858), .IN4(n19385), .Q(
        n7908) );
  OA22X1 U26672 ( .IN1(n2116), .IN2(n19441), .IN3(n2030), .IN4(n19418), .Q(
        n7909) );
  NAND4X0 U26673 ( .IN1(n7903), .IN2(n7904), .IN3(n7905), .IN4(n7906), .QN(
        s13_addr_o[18]) );
  OA22X1 U26674 ( .IN1(n1771), .IN2(n19375), .IN3(n1667), .IN4(n19353), .Q(
        n7903) );
  OA22X1 U26675 ( .IN1(n1943), .IN2(n19408), .IN3(n1857), .IN4(n19386), .Q(
        n7904) );
  OA22X1 U26676 ( .IN1(n2115), .IN2(n19441), .IN3(n2029), .IN4(n19419), .Q(
        n7905) );
  NAND4X0 U26677 ( .IN1(n7899), .IN2(n7900), .IN3(n7901), .IN4(n7902), .QN(
        s13_addr_o[19]) );
  OA22X1 U26678 ( .IN1(n1770), .IN2(n19375), .IN3(n1666), .IN4(n19353), .Q(
        n7899) );
  OA22X1 U26679 ( .IN1(n1942), .IN2(n19408), .IN3(n1856), .IN4(n19386), .Q(
        n7900) );
  OA22X1 U26680 ( .IN1(n2114), .IN2(n19441), .IN3(n2028), .IN4(n19419), .Q(
        n7901) );
  NAND4X0 U26681 ( .IN1(n7891), .IN2(n7892), .IN3(n7893), .IN4(n7894), .QN(
        s13_addr_o[20]) );
  OA22X1 U26682 ( .IN1(n1769), .IN2(n19374), .IN3(n1665), .IN4(n19354), .Q(
        n7891) );
  OA22X1 U26683 ( .IN1(n1941), .IN2(n19407), .IN3(n1855), .IN4(n19387), .Q(
        n7892) );
  OA22X1 U26684 ( .IN1(n2113), .IN2(n19440), .IN3(n2027), .IN4(n19420), .Q(
        n7893) );
  NAND4X0 U26685 ( .IN1(n7887), .IN2(n7888), .IN3(n7889), .IN4(n7890), .QN(
        s13_addr_o[21]) );
  OA22X1 U26686 ( .IN1(n1768), .IN2(n19374), .IN3(n1664), .IN4(n19354), .Q(
        n7887) );
  OA22X1 U26687 ( .IN1(n1940), .IN2(n19407), .IN3(n1854), .IN4(n19387), .Q(
        n7888) );
  OA22X1 U26688 ( .IN1(n2112), .IN2(n19440), .IN3(n2026), .IN4(n19420), .Q(
        n7889) );
  NAND4X0 U26689 ( .IN1(n7883), .IN2(n7884), .IN3(n7885), .IN4(n7886), .QN(
        s13_addr_o[22]) );
  OA22X1 U26690 ( .IN1(n1767), .IN2(n19373), .IN3(n1663), .IN4(n19354), .Q(
        n7883) );
  OA22X1 U26691 ( .IN1(n1939), .IN2(n19406), .IN3(n1853), .IN4(n19387), .Q(
        n7884) );
  OA22X1 U26692 ( .IN1(n2111), .IN2(n19439), .IN3(n2025), .IN4(n19420), .Q(
        n7885) );
  NAND4X0 U26693 ( .IN1(n7879), .IN2(n7880), .IN3(n7881), .IN4(n7882), .QN(
        s13_addr_o[23]) );
  OA22X1 U26694 ( .IN1(n1766), .IN2(n19374), .IN3(n1662), .IN4(n19355), .Q(
        n7879) );
  OA22X1 U26695 ( .IN1(n1938), .IN2(n19407), .IN3(n1852), .IN4(n19388), .Q(
        n7880) );
  OA22X1 U26696 ( .IN1(n2110), .IN2(n19440), .IN3(n2024), .IN4(n19421), .Q(
        n7881) );
  NAND4X0 U26697 ( .IN1(n7875), .IN2(n7876), .IN3(n7877), .IN4(n7878), .QN(
        s13_addr_o[24]) );
  OA22X1 U26698 ( .IN1(n1765), .IN2(n19380), .IN3(n1661), .IN4(n19355), .Q(
        n7875) );
  OA22X1 U26699 ( .IN1(n1937), .IN2(n19413), .IN3(n1851), .IN4(n19388), .Q(
        n7876) );
  OA22X1 U26700 ( .IN1(n2109), .IN2(n19446), .IN3(n2023), .IN4(n19421), .Q(
        n7877) );
  NAND4X0 U26701 ( .IN1(n7871), .IN2(n7872), .IN3(n7873), .IN4(n7874), .QN(
        s13_addr_o[25]) );
  OA22X1 U26702 ( .IN1(n1764), .IN2(n19376), .IN3(n1660), .IN4(n19355), .Q(
        n7871) );
  OA22X1 U26703 ( .IN1(n1936), .IN2(n19409), .IN3(n1850), .IN4(n19388), .Q(
        n7872) );
  OA22X1 U26704 ( .IN1(n2108), .IN2(n19442), .IN3(n2022), .IN4(n19421), .Q(
        n7873) );
  NAND4X0 U26705 ( .IN1(n7867), .IN2(n7868), .IN3(n7869), .IN4(n7870), .QN(
        s13_addr_o[26]) );
  OA22X1 U26706 ( .IN1(n1763), .IN2(n19375), .IN3(n1659), .IN4(n19356), .Q(
        n7867) );
  OA22X1 U26707 ( .IN1(n1935), .IN2(n19408), .IN3(n1849), .IN4(n19389), .Q(
        n7868) );
  OA22X1 U26708 ( .IN1(n2107), .IN2(n19441), .IN3(n2021), .IN4(n19422), .Q(
        n7869) );
  NAND4X0 U26709 ( .IN1(n7863), .IN2(n7864), .IN3(n7865), .IN4(n7866), .QN(
        s13_addr_o[27]) );
  OA22X1 U26710 ( .IN1(n1762), .IN2(n19374), .IN3(n1658), .IN4(n19356), .Q(
        n7863) );
  OA22X1 U26711 ( .IN1(n1934), .IN2(n19407), .IN3(n1848), .IN4(n19389), .Q(
        n7864) );
  OA22X1 U26712 ( .IN1(n2106), .IN2(n19440), .IN3(n2020), .IN4(n19422), .Q(
        n7865) );
  NAND4X0 U26713 ( .IN1(n7859), .IN2(n7860), .IN3(n7861), .IN4(n7862), .QN(
        s13_addr_o[28]) );
  OA22X1 U26714 ( .IN1(n1761), .IN2(n19374), .IN3(n1657), .IN4(n19356), .Q(
        n7859) );
  OA22X1 U26715 ( .IN1(n1933), .IN2(n19407), .IN3(n1847), .IN4(n19389), .Q(
        n7860) );
  OA22X1 U26716 ( .IN1(n2105), .IN2(n19440), .IN3(n2019), .IN4(n19422), .Q(
        n7861) );
  NAND4X0 U26717 ( .IN1(n7855), .IN2(n7856), .IN3(n7857), .IN4(n7858), .QN(
        s13_addr_o[29]) );
  OA22X1 U26718 ( .IN1(n1760), .IN2(n19378), .IN3(n1656), .IN4(n19357), .Q(
        n7855) );
  OA22X1 U26719 ( .IN1(n1932), .IN2(n19411), .IN3(n1846), .IN4(n19390), .Q(
        n7856) );
  OA22X1 U26720 ( .IN1(n2104), .IN2(n19444), .IN3(n2018), .IN4(n19423), .Q(
        n7857) );
  NAND4X0 U26721 ( .IN1(n7847), .IN2(n7848), .IN3(n7849), .IN4(n7850), .QN(
        s13_addr_o[30]) );
  OA22X1 U26722 ( .IN1(n1759), .IN2(n19379), .IN3(n1655), .IN4(n19357), .Q(
        n7847) );
  OA22X1 U26723 ( .IN1(n1931), .IN2(n19412), .IN3(n1845), .IN4(n19390), .Q(
        n7848) );
  OA22X1 U26724 ( .IN1(n2103), .IN2(n19445), .IN3(n2017), .IN4(n19423), .Q(
        n7849) );
  NAND4X0 U26725 ( .IN1(n7843), .IN2(n7844), .IN3(n7845), .IN4(n7846), .QN(
        s13_addr_o[31]) );
  OA22X1 U26726 ( .IN1(n1758), .IN2(n19377), .IN3(n1650), .IN4(n19358), .Q(
        n7843) );
  OA22X1 U26727 ( .IN1(n1930), .IN2(n19410), .IN3(n1844), .IN4(n19391), .Q(
        n7844) );
  OA22X1 U26728 ( .IN1(n2102), .IN2(n19443), .IN3(n2016), .IN4(n19424), .Q(
        n7845) );
  NAND4X0 U26729 ( .IN1(n7811), .IN2(n7812), .IN3(n7813), .IN4(n7814), .QN(
        s13_data_o[0]) );
  OA22X1 U26730 ( .IN1(n1741), .IN2(n19376), .IN3(n1636), .IN4(n19359), .Q(
        n7811) );
  OA22X1 U26731 ( .IN1(n1913), .IN2(n19409), .IN3(n1827), .IN4(n19392), .Q(
        n7812) );
  OA22X1 U26732 ( .IN1(n2085), .IN2(n19442), .IN3(n1999), .IN4(n19425), .Q(
        n7813) );
  NAND4X0 U26733 ( .IN1(n7767), .IN2(n7768), .IN3(n7769), .IN4(n7770), .QN(
        s13_data_o[1]) );
  OA22X1 U26734 ( .IN1(n1740), .IN2(n19378), .IN3(n1635), .IN4(n19357), .Q(
        n7767) );
  OA22X1 U26735 ( .IN1(n1912), .IN2(n19411), .IN3(n1826), .IN4(n19390), .Q(
        n7768) );
  OA22X1 U26736 ( .IN1(n2084), .IN2(n19444), .IN3(n1998), .IN4(n19423), .Q(
        n7769) );
  NAND4X0 U26737 ( .IN1(n7723), .IN2(n7724), .IN3(n7725), .IN4(n7726), .QN(
        s13_data_o[2]) );
  OA22X1 U26738 ( .IN1(n1739), .IN2(n19379), .IN3(n1634), .IN4(n19350), .Q(
        n7723) );
  OA22X1 U26739 ( .IN1(n1911), .IN2(n19412), .IN3(n1825), .IN4(n19383), .Q(
        n7724) );
  OA22X1 U26740 ( .IN1(n2083), .IN2(n19445), .IN3(n1997), .IN4(n19416), .Q(
        n7725) );
  NAND4X0 U26741 ( .IN1(n7711), .IN2(n7712), .IN3(n7713), .IN4(n7714), .QN(
        s13_data_o[3]) );
  OA22X1 U26742 ( .IN1(n1738), .IN2(n19377), .IN3(n1633), .IN4(n19352), .Q(
        n7711) );
  OA22X1 U26743 ( .IN1(n1910), .IN2(n19410), .IN3(n1824), .IN4(n19385), .Q(
        n7712) );
  OA22X1 U26744 ( .IN1(n2082), .IN2(n19443), .IN3(n1996), .IN4(n19418), .Q(
        n7713) );
  NAND4X0 U26745 ( .IN1(n7707), .IN2(n7708), .IN3(n7709), .IN4(n7710), .QN(
        s13_data_o[4]) );
  OA22X1 U26746 ( .IN1(n1737), .IN2(n19378), .IN3(n1632), .IN4(n19367), .Q(
        n7707) );
  OA22X1 U26747 ( .IN1(n1909), .IN2(n19411), .IN3(n1823), .IN4(n19400), .Q(
        n7708) );
  OA22X1 U26748 ( .IN1(n2081), .IN2(n19444), .IN3(n1995), .IN4(n19433), .Q(
        n7709) );
  NAND4X0 U26749 ( .IN1(n7703), .IN2(n7704), .IN3(n7705), .IN4(n7706), .QN(
        s13_data_o[5]) );
  OA22X1 U26750 ( .IN1(n1736), .IN2(n19379), .IN3(n1631), .IN4(n19365), .Q(
        n7703) );
  OA22X1 U26751 ( .IN1(n1908), .IN2(n19412), .IN3(n1822), .IN4(n19398), .Q(
        n7704) );
  OA22X1 U26752 ( .IN1(n2080), .IN2(n19445), .IN3(n1994), .IN4(n19431), .Q(
        n7705) );
  NAND4X0 U26753 ( .IN1(n7699), .IN2(n7700), .IN3(n7701), .IN4(n7702), .QN(
        s13_data_o[6]) );
  OA22X1 U26754 ( .IN1(n1735), .IN2(n19375), .IN3(n1630), .IN4(n19365), .Q(
        n7699) );
  OA22X1 U26755 ( .IN1(n1907), .IN2(n19408), .IN3(n1821), .IN4(n19398), .Q(
        n7700) );
  OA22X1 U26756 ( .IN1(n2079), .IN2(n19441), .IN3(n1993), .IN4(n19431), .Q(
        n7701) );
  NAND4X0 U26757 ( .IN1(n7695), .IN2(n7696), .IN3(n7697), .IN4(n7698), .QN(
        s13_data_o[7]) );
  OA22X1 U26758 ( .IN1(n1734), .IN2(n19373), .IN3(n1629), .IN4(n19365), .Q(
        n7695) );
  OA22X1 U26759 ( .IN1(n1906), .IN2(n19406), .IN3(n1820), .IN4(n19398), .Q(
        n7696) );
  OA22X1 U26760 ( .IN1(n2078), .IN2(n19439), .IN3(n1992), .IN4(n19431), .Q(
        n7697) );
  NAND4X0 U26761 ( .IN1(n7691), .IN2(n7692), .IN3(n7693), .IN4(n7694), .QN(
        s13_data_o[8]) );
  OA22X1 U26762 ( .IN1(n1733), .IN2(n19380), .IN3(n1628), .IN4(n19365), .Q(
        n7691) );
  OA22X1 U26763 ( .IN1(n1905), .IN2(n19413), .IN3(n1819), .IN4(n19398), .Q(
        n7692) );
  OA22X1 U26764 ( .IN1(n2077), .IN2(n19446), .IN3(n1991), .IN4(n19431), .Q(
        n7693) );
  NAND4X0 U26765 ( .IN1(n7687), .IN2(n7688), .IN3(n7689), .IN4(n7690), .QN(
        s13_data_o[9]) );
  OA22X1 U26766 ( .IN1(n1732), .IN2(n19373), .IN3(n1627), .IN4(n19366), .Q(
        n7687) );
  OA22X1 U26767 ( .IN1(n1904), .IN2(n19406), .IN3(n1818), .IN4(n19399), .Q(
        n7688) );
  OA22X1 U26768 ( .IN1(n2076), .IN2(n19439), .IN3(n1990), .IN4(n19432), .Q(
        n7689) );
  NAND4X0 U26769 ( .IN1(n7807), .IN2(n7808), .IN3(n7809), .IN4(n7810), .QN(
        s13_data_o[10]) );
  OA22X1 U26770 ( .IN1(n1731), .IN2(n19375), .IN3(n1626), .IN4(n19360), .Q(
        n7807) );
  OA22X1 U26771 ( .IN1(n1903), .IN2(n19408), .IN3(n1817), .IN4(n19393), .Q(
        n7808) );
  OA22X1 U26772 ( .IN1(n2075), .IN2(n19441), .IN3(n1989), .IN4(n19426), .Q(
        n7809) );
  NAND4X0 U26773 ( .IN1(n7803), .IN2(n7804), .IN3(n7805), .IN4(n7806), .QN(
        s13_data_o[11]) );
  OA22X1 U26774 ( .IN1(n1730), .IN2(n19380), .IN3(n1625), .IN4(n19360), .Q(
        n7803) );
  OA22X1 U26775 ( .IN1(n1902), .IN2(n19413), .IN3(n1816), .IN4(n19393), .Q(
        n7804) );
  OA22X1 U26776 ( .IN1(n2074), .IN2(n19446), .IN3(n1988), .IN4(n19426), .Q(
        n7805) );
  NAND4X0 U26777 ( .IN1(n7799), .IN2(n7800), .IN3(n7801), .IN4(n7802), .QN(
        s13_data_o[12]) );
  OA22X1 U26778 ( .IN1(n1729), .IN2(n19376), .IN3(n1624), .IN4(n19360), .Q(
        n7799) );
  OA22X1 U26779 ( .IN1(n1901), .IN2(n19409), .IN3(n1815), .IN4(n19393), .Q(
        n7800) );
  OA22X1 U26780 ( .IN1(n2073), .IN2(n19442), .IN3(n1987), .IN4(n19426), .Q(
        n7801) );
  NAND4X0 U26781 ( .IN1(n7795), .IN2(n7796), .IN3(n7797), .IN4(n7798), .QN(
        s13_data_o[13]) );
  OA22X1 U26782 ( .IN1(n1728), .IN2(n19377), .IN3(n1623), .IN4(n19354), .Q(
        n7795) );
  OA22X1 U26783 ( .IN1(n1900), .IN2(n19410), .IN3(n1814), .IN4(n19387), .Q(
        n7796) );
  OA22X1 U26784 ( .IN1(n2072), .IN2(n19443), .IN3(n1986), .IN4(n19420), .Q(
        n7797) );
  NAND4X0 U26785 ( .IN1(n7791), .IN2(n7792), .IN3(n7793), .IN4(n7794), .QN(
        s13_data_o[14]) );
  OA22X1 U26786 ( .IN1(n1727), .IN2(n19377), .IN3(n1622), .IN4(n19359), .Q(
        n7791) );
  OA22X1 U26787 ( .IN1(n1899), .IN2(n19410), .IN3(n1813), .IN4(n19392), .Q(
        n7792) );
  OA22X1 U26788 ( .IN1(n2071), .IN2(n19443), .IN3(n1985), .IN4(n19425), .Q(
        n7793) );
  NAND4X0 U26789 ( .IN1(n7787), .IN2(n7788), .IN3(n7789), .IN4(n7790), .QN(
        s13_data_o[15]) );
  OA22X1 U26790 ( .IN1(n1726), .IN2(n19377), .IN3(n1621), .IN4(n19360), .Q(
        n7787) );
  OA22X1 U26791 ( .IN1(n1898), .IN2(n19410), .IN3(n1812), .IN4(n19393), .Q(
        n7788) );
  OA22X1 U26792 ( .IN1(n2070), .IN2(n19443), .IN3(n1984), .IN4(n19426), .Q(
        n7789) );
  NAND4X0 U26793 ( .IN1(n7783), .IN2(n7784), .IN3(n7785), .IN4(n7786), .QN(
        s13_data_o[16]) );
  OA22X1 U26794 ( .IN1(n1725), .IN2(n19377), .IN3(n1620), .IN4(n19361), .Q(
        n7783) );
  OA22X1 U26795 ( .IN1(n1897), .IN2(n19410), .IN3(n1811), .IN4(n19394), .Q(
        n7784) );
  OA22X1 U26796 ( .IN1(n2069), .IN2(n19443), .IN3(n1983), .IN4(n19427), .Q(
        n7785) );
  NAND4X0 U26797 ( .IN1(n7779), .IN2(n7780), .IN3(n7781), .IN4(n7782), .QN(
        s13_data_o[17]) );
  OA22X1 U26798 ( .IN1(n1724), .IN2(n19378), .IN3(n1619), .IN4(n19361), .Q(
        n7779) );
  OA22X1 U26799 ( .IN1(n1896), .IN2(n19411), .IN3(n1810), .IN4(n19394), .Q(
        n7780) );
  OA22X1 U26800 ( .IN1(n2068), .IN2(n19444), .IN3(n1982), .IN4(n19427), .Q(
        n7781) );
  NAND4X0 U26801 ( .IN1(n7775), .IN2(n7776), .IN3(n7777), .IN4(n7778), .QN(
        s13_data_o[18]) );
  OA22X1 U26802 ( .IN1(n1723), .IN2(n19378), .IN3(n1618), .IN4(n19361), .Q(
        n7775) );
  OA22X1 U26803 ( .IN1(n1895), .IN2(n19411), .IN3(n1809), .IN4(n19394), .Q(
        n7776) );
  OA22X1 U26804 ( .IN1(n2067), .IN2(n19444), .IN3(n1981), .IN4(n19427), .Q(
        n7777) );
  NAND4X0 U26805 ( .IN1(n7771), .IN2(n7772), .IN3(n7773), .IN4(n7774), .QN(
        s13_data_o[19]) );
  OA22X1 U26806 ( .IN1(n1722), .IN2(n19378), .IN3(n1617), .IN4(n19361), .Q(
        n7771) );
  OA22X1 U26807 ( .IN1(n1894), .IN2(n19411), .IN3(n1808), .IN4(n19394), .Q(
        n7772) );
  OA22X1 U26808 ( .IN1(n2066), .IN2(n19444), .IN3(n1980), .IN4(n19427), .Q(
        n7773) );
  NAND4X0 U26809 ( .IN1(n7763), .IN2(n7764), .IN3(n7765), .IN4(n7766), .QN(
        s13_data_o[20]) );
  OA22X1 U26810 ( .IN1(n1721), .IN2(n19379), .IN3(n1616), .IN4(n19358), .Q(
        n7763) );
  OA22X1 U26811 ( .IN1(n1893), .IN2(n19412), .IN3(n1807), .IN4(n19391), .Q(
        n7764) );
  OA22X1 U26812 ( .IN1(n2065), .IN2(n19445), .IN3(n1979), .IN4(n19424), .Q(
        n7765) );
  NAND4X0 U26813 ( .IN1(n7759), .IN2(n7760), .IN3(n7761), .IN4(n7762), .QN(
        s13_data_o[21]) );
  OA22X1 U26814 ( .IN1(n1720), .IN2(n19379), .IN3(n1615), .IN4(n19362), .Q(
        n7759) );
  OA22X1 U26815 ( .IN1(n1892), .IN2(n19412), .IN3(n1806), .IN4(n19395), .Q(
        n7760) );
  OA22X1 U26816 ( .IN1(n2064), .IN2(n19445), .IN3(n1978), .IN4(n19428), .Q(
        n7761) );
  NAND4X0 U26817 ( .IN1(n7755), .IN2(n7756), .IN3(n7757), .IN4(n7758), .QN(
        s13_data_o[22]) );
  OA22X1 U26818 ( .IN1(n1719), .IN2(n19377), .IN3(n1614), .IN4(n19362), .Q(
        n7755) );
  OA22X1 U26819 ( .IN1(n1891), .IN2(n19410), .IN3(n1805), .IN4(n19395), .Q(
        n7756) );
  OA22X1 U26820 ( .IN1(n2063), .IN2(n19443), .IN3(n1977), .IN4(n19428), .Q(
        n7757) );
  NAND4X0 U26821 ( .IN1(n7751), .IN2(n7752), .IN3(n7753), .IN4(n7754), .QN(
        s13_data_o[23]) );
  OA22X1 U26822 ( .IN1(n1718), .IN2(n19378), .IN3(n1613), .IN4(n19362), .Q(
        n7751) );
  OA22X1 U26823 ( .IN1(n1890), .IN2(n19411), .IN3(n1804), .IN4(n19395), .Q(
        n7752) );
  OA22X1 U26824 ( .IN1(n2062), .IN2(n19444), .IN3(n1976), .IN4(n19428), .Q(
        n7753) );
  NAND4X0 U26825 ( .IN1(n7747), .IN2(n7748), .IN3(n7749), .IN4(n7750), .QN(
        s13_data_o[24]) );
  OA22X1 U26826 ( .IN1(n1717), .IN2(n19376), .IN3(n1612), .IN4(n19363), .Q(
        n7747) );
  OA22X1 U26827 ( .IN1(n1889), .IN2(n19409), .IN3(n1803), .IN4(n19396), .Q(
        n7748) );
  OA22X1 U26828 ( .IN1(n2061), .IN2(n19442), .IN3(n1975), .IN4(n19429), .Q(
        n7749) );
  NAND4X0 U26829 ( .IN1(n7743), .IN2(n7744), .IN3(n7745), .IN4(n7746), .QN(
        s13_data_o[25]) );
  OA22X1 U26830 ( .IN1(n1716), .IN2(n19376), .IN3(n1611), .IN4(n19363), .Q(
        n7743) );
  OA22X1 U26831 ( .IN1(n1888), .IN2(n19409), .IN3(n1802), .IN4(n19396), .Q(
        n7744) );
  OA22X1 U26832 ( .IN1(n2060), .IN2(n19442), .IN3(n1974), .IN4(n19429), .Q(
        n7745) );
  NAND4X0 U26833 ( .IN1(n7739), .IN2(n7740), .IN3(n7741), .IN4(n7742), .QN(
        s13_data_o[26]) );
  OA22X1 U26834 ( .IN1(n1715), .IN2(n19375), .IN3(n1610), .IN4(n19363), .Q(
        n7739) );
  OA22X1 U26835 ( .IN1(n1887), .IN2(n19408), .IN3(n1801), .IN4(n19396), .Q(
        n7740) );
  OA22X1 U26836 ( .IN1(n2059), .IN2(n19441), .IN3(n1973), .IN4(n19429), .Q(
        n7741) );
  NAND4X0 U26837 ( .IN1(n7735), .IN2(n7736), .IN3(n7737), .IN4(n7738), .QN(
        s13_data_o[27]) );
  OA22X1 U26838 ( .IN1(n1714), .IN2(n19378), .IN3(n1609), .IN4(n19364), .Q(
        n7735) );
  OA22X1 U26839 ( .IN1(n1886), .IN2(n19411), .IN3(n1800), .IN4(n19397), .Q(
        n7736) );
  OA22X1 U26840 ( .IN1(n2058), .IN2(n19444), .IN3(n1972), .IN4(n19430), .Q(
        n7737) );
  NAND4X0 U26841 ( .IN1(n7731), .IN2(n7732), .IN3(n7733), .IN4(n7734), .QN(
        s13_data_o[28]) );
  OA22X1 U26842 ( .IN1(n1713), .IN2(n19379), .IN3(n1608), .IN4(n19364), .Q(
        n7731) );
  OA22X1 U26843 ( .IN1(n1885), .IN2(n19412), .IN3(n1799), .IN4(n19397), .Q(
        n7732) );
  OA22X1 U26844 ( .IN1(n2057), .IN2(n19445), .IN3(n1971), .IN4(n19430), .Q(
        n7733) );
  NAND4X0 U26845 ( .IN1(n7727), .IN2(n7728), .IN3(n7729), .IN4(n7730), .QN(
        s13_data_o[29]) );
  OA22X1 U26846 ( .IN1(n1712), .IN2(n19379), .IN3(n1607), .IN4(n19364), .Q(
        n7727) );
  OA22X1 U26847 ( .IN1(n1884), .IN2(n19412), .IN3(n1798), .IN4(n19397), .Q(
        n7728) );
  OA22X1 U26848 ( .IN1(n2056), .IN2(n19445), .IN3(n1970), .IN4(n19430), .Q(
        n7729) );
  NAND4X0 U26849 ( .IN1(n7719), .IN2(n7720), .IN3(n7721), .IN4(n7722), .QN(
        s13_data_o[30]) );
  OA22X1 U26850 ( .IN1(n1711), .IN2(n19379), .IN3(n1606), .IN4(n19366), .Q(
        n7719) );
  OA22X1 U26851 ( .IN1(n1883), .IN2(n19412), .IN3(n1797), .IN4(n19399), .Q(
        n7720) );
  OA22X1 U26852 ( .IN1(n2055), .IN2(n19445), .IN3(n1969), .IN4(n19432), .Q(
        n7721) );
  NAND4X0 U26853 ( .IN1(n7715), .IN2(n7716), .IN3(n7717), .IN4(n7718), .QN(
        s13_data_o[31]) );
  OA22X1 U26854 ( .IN1(n1710), .IN2(n19377), .IN3(n1605), .IN4(n19351), .Q(
        n7715) );
  OA22X1 U26855 ( .IN1(n1882), .IN2(n19410), .IN3(n1796), .IN4(n19384), .Q(
        n7716) );
  OA22X1 U26856 ( .IN1(n2054), .IN2(n19443), .IN3(n1968), .IN4(n19417), .Q(
        n7717) );
  NAND4X0 U26857 ( .IN1(n7955), .IN2(n7956), .IN3(n7957), .IN4(n7958), .QN(
        s12_stb_o) );
  OA22X1 U26858 ( .IN1(n1795), .IN2(n7965), .IN3(n1709), .IN4(n7966), .Q(n7955) );
  OA22X1 U26859 ( .IN1(n1967), .IN2(n7963), .IN3(n1881), .IN4(n7964), .Q(n7956) );
  OA22X1 U26860 ( .IN1(n2139), .IN2(n7961), .IN3(n2053), .IN4(n7962), .Q(n7957) );
  NAND4X0 U26861 ( .IN1(n7943), .IN2(n7944), .IN3(n7945), .IN4(n7946), .QN(
        s12_we_o) );
  OA22X1 U26862 ( .IN1(n1794), .IN2(n19241), .IN3(n1708), .IN4(n19235), .Q(
        n7943) );
  OA22X1 U26863 ( .IN1(n1966), .IN2(n19274), .IN3(n1880), .IN4(n19268), .Q(
        n7944) );
  OA22X1 U26864 ( .IN1(n2138), .IN2(n19307), .IN3(n2052), .IN4(n19301), .Q(
        n7945) );
  NAND4X0 U26865 ( .IN1(n7979), .IN2(n7980), .IN3(n7981), .IN4(n7982), .QN(
        s12_sel_o[0]) );
  OA22X1 U26866 ( .IN1(n1793), .IN2(n19248), .IN3(n1707), .IN4(n19234), .Q(
        n7979) );
  OA22X1 U26867 ( .IN1(n1965), .IN2(n19281), .IN3(n1879), .IN4(n19267), .Q(
        n7980) );
  OA22X1 U26868 ( .IN1(n2137), .IN2(n19314), .IN3(n2051), .IN4(n19300), .Q(
        n7981) );
  NAND4X0 U26869 ( .IN1(n7975), .IN2(n7976), .IN3(n7977), .IN4(n7978), .QN(
        s12_sel_o[1]) );
  OA22X1 U26870 ( .IN1(n1792), .IN2(n19248), .IN3(n1706), .IN4(n19234), .Q(
        n7975) );
  OA22X1 U26871 ( .IN1(n1964), .IN2(n19281), .IN3(n1878), .IN4(n19267), .Q(
        n7976) );
  OA22X1 U26872 ( .IN1(n2136), .IN2(n19314), .IN3(n2050), .IN4(n19300), .Q(
        n7977) );
  NAND4X0 U26873 ( .IN1(n7971), .IN2(n7972), .IN3(n7973), .IN4(n7974), .QN(
        s12_sel_o[2]) );
  OA22X1 U26874 ( .IN1(n1791), .IN2(n19248), .IN3(n1705), .IN4(n19235), .Q(
        n7971) );
  OA22X1 U26875 ( .IN1(n1963), .IN2(n19281), .IN3(n1877), .IN4(n19268), .Q(
        n7972) );
  OA22X1 U26876 ( .IN1(n2135), .IN2(n19314), .IN3(n2049), .IN4(n19301), .Q(
        n7973) );
  NAND4X0 U26877 ( .IN1(n7967), .IN2(n7968), .IN3(n7969), .IN4(n7970), .QN(
        s12_sel_o[3]) );
  OA22X1 U26878 ( .IN1(n1790), .IN2(n19248), .IN3(n1704), .IN4(n19235), .Q(
        n7967) );
  OA22X1 U26879 ( .IN1(n1962), .IN2(n19281), .IN3(n1876), .IN4(n19268), .Q(
        n7968) );
  OA22X1 U26880 ( .IN1(n2134), .IN2(n19314), .IN3(n2048), .IN4(n19301), .Q(
        n7969) );
  NAND4X0 U26881 ( .IN1(n8235), .IN2(n8236), .IN3(n8237), .IN4(n8238), .QN(
        s12_addr_o[0]) );
  OA22X1 U26882 ( .IN1(n1789), .IN2(n19241), .IN3(n1703), .IN4(n19218), .Q(
        n8235) );
  OA22X1 U26883 ( .IN1(n1961), .IN2(n19274), .IN3(n1875), .IN4(n19251), .Q(
        n8236) );
  OA22X1 U26884 ( .IN1(n2133), .IN2(n19307), .IN3(n2047), .IN4(n19284), .Q(
        n8237) );
  NAND4X0 U26885 ( .IN1(n8191), .IN2(n8192), .IN3(n8193), .IN4(n8194), .QN(
        s12_addr_o[1]) );
  OA22X1 U26886 ( .IN1(n1788), .IN2(n19243), .IN3(n1702), .IN4(n19221), .Q(
        n8191) );
  OA22X1 U26887 ( .IN1(n1960), .IN2(n19276), .IN3(n1874), .IN4(n19254), .Q(
        n8192) );
  OA22X1 U26888 ( .IN1(n2132), .IN2(n19309), .IN3(n2046), .IN4(n19287), .Q(
        n8193) );
  NAND4X0 U26889 ( .IN1(n8147), .IN2(n8148), .IN3(n8149), .IN4(n8150), .QN(
        s12_addr_o[2]) );
  OA22X1 U26890 ( .IN1(n1787), .IN2(n19243), .IN3(n1701), .IN4(n19225), .Q(
        n8147) );
  OA22X1 U26891 ( .IN1(n1959), .IN2(n19276), .IN3(n1873), .IN4(n19258), .Q(
        n8148) );
  OA22X1 U26892 ( .IN1(n2131), .IN2(n19309), .IN3(n2045), .IN4(n19291), .Q(
        n8149) );
  NAND4X0 U26893 ( .IN1(n8135), .IN2(n8136), .IN3(n8137), .IN4(n8138), .QN(
        s12_addr_o[3]) );
  OA22X1 U26894 ( .IN1(n1786), .IN2(n19248), .IN3(n1699), .IN4(n19226), .Q(
        n8135) );
  OA22X1 U26895 ( .IN1(n1958), .IN2(n19281), .IN3(n1872), .IN4(n19259), .Q(
        n8136) );
  OA22X1 U26896 ( .IN1(n2130), .IN2(n19314), .IN3(n2044), .IN4(n19292), .Q(
        n8137) );
  NAND4X0 U26897 ( .IN1(n8131), .IN2(n8132), .IN3(n8133), .IN4(n8134), .QN(
        s12_addr_o[4]) );
  OA22X1 U26898 ( .IN1(n1785), .IN2(n19241), .IN3(n1697), .IN4(n19226), .Q(
        n8131) );
  OA22X1 U26899 ( .IN1(n1957), .IN2(n19274), .IN3(n1871), .IN4(n19259), .Q(
        n8132) );
  OA22X1 U26900 ( .IN1(n2129), .IN2(n19307), .IN3(n2043), .IN4(n19292), .Q(
        n8133) );
  NAND4X0 U26901 ( .IN1(n8127), .IN2(n8128), .IN3(n8129), .IN4(n8130), .QN(
        s12_addr_o[5]) );
  OA22X1 U26902 ( .IN1(n1784), .IN2(n19248), .IN3(n1696), .IN4(n19225), .Q(
        n8127) );
  OA22X1 U26903 ( .IN1(n1956), .IN2(n19281), .IN3(n1870), .IN4(n19258), .Q(
        n8128) );
  OA22X1 U26904 ( .IN1(n2128), .IN2(n19314), .IN3(n2042), .IN4(n19291), .Q(
        n8129) );
  NAND4X0 U26905 ( .IN1(n8123), .IN2(n8124), .IN3(n8125), .IN4(n8126), .QN(
        s12_addr_o[6]) );
  OA22X1 U26906 ( .IN1(n1783), .IN2(n19244), .IN3(n1679), .IN4(n19226), .Q(
        n8123) );
  OA22X1 U26907 ( .IN1(n1955), .IN2(n19277), .IN3(n1869), .IN4(n19259), .Q(
        n8124) );
  OA22X1 U26908 ( .IN1(n2127), .IN2(n19310), .IN3(n2041), .IN4(n19292), .Q(
        n8125) );
  NAND4X0 U26909 ( .IN1(n8119), .IN2(n8120), .IN3(n8121), .IN4(n8122), .QN(
        s12_addr_o[7]) );
  OA22X1 U26910 ( .IN1(n1782), .IN2(n19244), .IN3(n1678), .IN4(n19218), .Q(
        n8119) );
  OA22X1 U26911 ( .IN1(n1954), .IN2(n19277), .IN3(n1868), .IN4(n19251), .Q(
        n8120) );
  OA22X1 U26912 ( .IN1(n2126), .IN2(n19310), .IN3(n2040), .IN4(n19291), .Q(
        n8121) );
  NAND4X0 U26913 ( .IN1(n8115), .IN2(n8116), .IN3(n8117), .IN4(n8118), .QN(
        s12_addr_o[8]) );
  OA22X1 U26914 ( .IN1(n1781), .IN2(n19244), .IN3(n1677), .IN4(n19227), .Q(
        n8115) );
  OA22X1 U26915 ( .IN1(n1953), .IN2(n19277), .IN3(n1867), .IN4(n19260), .Q(
        n8116) );
  OA22X1 U26916 ( .IN1(n2125), .IN2(n19310), .IN3(n2039), .IN4(n19293), .Q(
        n8117) );
  NAND4X0 U26917 ( .IN1(n8111), .IN2(n8112), .IN3(n8113), .IN4(n8114), .QN(
        s12_addr_o[9]) );
  OA22X1 U26918 ( .IN1(n1780), .IN2(n19244), .IN3(n1676), .IN4(n19227), .Q(
        n8111) );
  OA22X1 U26919 ( .IN1(n1952), .IN2(n19277), .IN3(n1866), .IN4(n19260), .Q(
        n8112) );
  OA22X1 U26920 ( .IN1(n2124), .IN2(n19310), .IN3(n2038), .IN4(n19293), .Q(
        n8113) );
  NAND4X0 U26921 ( .IN1(n8231), .IN2(n8232), .IN3(n8233), .IN4(n8234), .QN(
        s12_addr_o[10]) );
  OA22X1 U26922 ( .IN1(n1779), .IN2(n19241), .IN3(n1675), .IN4(n19218), .Q(
        n8231) );
  OA22X1 U26923 ( .IN1(n1951), .IN2(n19274), .IN3(n1865), .IN4(n19251), .Q(
        n8232) );
  OA22X1 U26924 ( .IN1(n2123), .IN2(n19307), .IN3(n2037), .IN4(n19284), .Q(
        n8233) );
  NAND4X0 U26925 ( .IN1(n8227), .IN2(n8228), .IN3(n8229), .IN4(n8230), .QN(
        s12_addr_o[11]) );
  OA22X1 U26926 ( .IN1(n1778), .IN2(n19241), .IN3(n1674), .IN4(n19218), .Q(
        n8227) );
  OA22X1 U26927 ( .IN1(n1950), .IN2(n19274), .IN3(n1864), .IN4(n19251), .Q(
        n8228) );
  OA22X1 U26928 ( .IN1(n2122), .IN2(n19307), .IN3(n2036), .IN4(n19284), .Q(
        n8229) );
  NAND4X0 U26929 ( .IN1(n8223), .IN2(n8224), .IN3(n8225), .IN4(n8226), .QN(
        s12_addr_o[12]) );
  OA22X1 U26930 ( .IN1(n1777), .IN2(n19241), .IN3(n1673), .IN4(n19219), .Q(
        n8223) );
  OA22X1 U26931 ( .IN1(n1949), .IN2(n19274), .IN3(n1863), .IN4(n19252), .Q(
        n8224) );
  OA22X1 U26932 ( .IN1(n2121), .IN2(n19307), .IN3(n2035), .IN4(n19285), .Q(
        n8225) );
  NAND4X0 U26933 ( .IN1(n8219), .IN2(n8220), .IN3(n8221), .IN4(n8222), .QN(
        s12_addr_o[13]) );
  OA22X1 U26934 ( .IN1(n1776), .IN2(n19242), .IN3(n1672), .IN4(n19219), .Q(
        n8219) );
  OA22X1 U26935 ( .IN1(n1948), .IN2(n19275), .IN3(n1862), .IN4(n19252), .Q(
        n8220) );
  OA22X1 U26936 ( .IN1(n2120), .IN2(n19308), .IN3(n2034), .IN4(n19285), .Q(
        n8221) );
  NAND4X0 U26937 ( .IN1(n8215), .IN2(n8216), .IN3(n8217), .IN4(n8218), .QN(
        s12_addr_o[14]) );
  OA22X1 U26938 ( .IN1(n1775), .IN2(n19242), .IN3(n1671), .IN4(n19219), .Q(
        n8215) );
  OA22X1 U26939 ( .IN1(n1947), .IN2(n19275), .IN3(n1861), .IN4(n19252), .Q(
        n8216) );
  OA22X1 U26940 ( .IN1(n2119), .IN2(n19308), .IN3(n2033), .IN4(n19285), .Q(
        n8217) );
  NAND4X0 U26941 ( .IN1(n8211), .IN2(n8212), .IN3(n8213), .IN4(n8214), .QN(
        s12_addr_o[15]) );
  OA22X1 U26942 ( .IN1(n1774), .IN2(n19242), .IN3(n1670), .IN4(n19220), .Q(
        n8211) );
  OA22X1 U26943 ( .IN1(n1946), .IN2(n19275), .IN3(n1860), .IN4(n19253), .Q(
        n8212) );
  OA22X1 U26944 ( .IN1(n2118), .IN2(n19308), .IN3(n2032), .IN4(n19286), .Q(
        n8213) );
  NAND4X0 U26945 ( .IN1(n8207), .IN2(n8208), .IN3(n8209), .IN4(n8210), .QN(
        s12_addr_o[16]) );
  OA22X1 U26946 ( .IN1(n1773), .IN2(n19242), .IN3(n1669), .IN4(n19220), .Q(
        n8207) );
  OA22X1 U26947 ( .IN1(n1945), .IN2(n19275), .IN3(n1859), .IN4(n19253), .Q(
        n8208) );
  OA22X1 U26948 ( .IN1(n2117), .IN2(n19308), .IN3(n2031), .IN4(n19286), .Q(
        n8209) );
  NAND4X0 U26949 ( .IN1(n8203), .IN2(n8204), .IN3(n8205), .IN4(n8206), .QN(
        s12_addr_o[17]) );
  OA22X1 U26950 ( .IN1(n1772), .IN2(n19243), .IN3(n1668), .IN4(n19220), .Q(
        n8203) );
  OA22X1 U26951 ( .IN1(n1944), .IN2(n19276), .IN3(n1858), .IN4(n19253), .Q(
        n8204) );
  OA22X1 U26952 ( .IN1(n2116), .IN2(n19309), .IN3(n2030), .IN4(n19286), .Q(
        n8205) );
  NAND4X0 U26953 ( .IN1(n8199), .IN2(n8200), .IN3(n8201), .IN4(n8202), .QN(
        s12_addr_o[18]) );
  OA22X1 U26954 ( .IN1(n1771), .IN2(n19243), .IN3(n1667), .IN4(n19221), .Q(
        n8199) );
  OA22X1 U26955 ( .IN1(n1943), .IN2(n19276), .IN3(n1857), .IN4(n19254), .Q(
        n8200) );
  OA22X1 U26956 ( .IN1(n2115), .IN2(n19309), .IN3(n2029), .IN4(n19287), .Q(
        n8201) );
  NAND4X0 U26957 ( .IN1(n8195), .IN2(n8196), .IN3(n8197), .IN4(n8198), .QN(
        s12_addr_o[19]) );
  OA22X1 U26958 ( .IN1(n1770), .IN2(n19243), .IN3(n1666), .IN4(n19221), .Q(
        n8195) );
  OA22X1 U26959 ( .IN1(n1942), .IN2(n19276), .IN3(n1856), .IN4(n19254), .Q(
        n8196) );
  OA22X1 U26960 ( .IN1(n2114), .IN2(n19309), .IN3(n2028), .IN4(n19287), .Q(
        n8197) );
  NAND4X0 U26961 ( .IN1(n8187), .IN2(n8188), .IN3(n8189), .IN4(n8190), .QN(
        s12_addr_o[20]) );
  OA22X1 U26962 ( .IN1(n1769), .IN2(n19242), .IN3(n1665), .IN4(n19222), .Q(
        n8187) );
  OA22X1 U26963 ( .IN1(n1941), .IN2(n19275), .IN3(n1855), .IN4(n19255), .Q(
        n8188) );
  OA22X1 U26964 ( .IN1(n2113), .IN2(n19308), .IN3(n2027), .IN4(n19288), .Q(
        n8189) );
  NAND4X0 U26965 ( .IN1(n8183), .IN2(n8184), .IN3(n8185), .IN4(n8186), .QN(
        s12_addr_o[21]) );
  OA22X1 U26966 ( .IN1(n1768), .IN2(n19242), .IN3(n1664), .IN4(n19222), .Q(
        n8183) );
  OA22X1 U26967 ( .IN1(n1940), .IN2(n19275), .IN3(n1854), .IN4(n19255), .Q(
        n8184) );
  OA22X1 U26968 ( .IN1(n2112), .IN2(n19308), .IN3(n2026), .IN4(n19288), .Q(
        n8185) );
  NAND4X0 U26969 ( .IN1(n8179), .IN2(n8180), .IN3(n8181), .IN4(n8182), .QN(
        s12_addr_o[22]) );
  OA22X1 U26970 ( .IN1(n1767), .IN2(n19241), .IN3(n1663), .IN4(n19222), .Q(
        n8179) );
  OA22X1 U26971 ( .IN1(n1939), .IN2(n19274), .IN3(n1853), .IN4(n19255), .Q(
        n8180) );
  OA22X1 U26972 ( .IN1(n2111), .IN2(n19307), .IN3(n2025), .IN4(n19288), .Q(
        n8181) );
  NAND4X0 U26973 ( .IN1(n8175), .IN2(n8176), .IN3(n8177), .IN4(n8178), .QN(
        s12_addr_o[23]) );
  OA22X1 U26974 ( .IN1(n1766), .IN2(n19242), .IN3(n1662), .IN4(n19223), .Q(
        n8175) );
  OA22X1 U26975 ( .IN1(n1938), .IN2(n19275), .IN3(n1852), .IN4(n19256), .Q(
        n8176) );
  OA22X1 U26976 ( .IN1(n2110), .IN2(n19308), .IN3(n2024), .IN4(n19289), .Q(
        n8177) );
  NAND4X0 U26977 ( .IN1(n8171), .IN2(n8172), .IN3(n8173), .IN4(n8174), .QN(
        s12_addr_o[24]) );
  OA22X1 U26978 ( .IN1(n1765), .IN2(n19248), .IN3(n1661), .IN4(n19223), .Q(
        n8171) );
  OA22X1 U26979 ( .IN1(n1937), .IN2(n19281), .IN3(n1851), .IN4(n19256), .Q(
        n8172) );
  OA22X1 U26980 ( .IN1(n2109), .IN2(n19314), .IN3(n2023), .IN4(n19289), .Q(
        n8173) );
  NAND4X0 U26981 ( .IN1(n8167), .IN2(n8168), .IN3(n8169), .IN4(n8170), .QN(
        s12_addr_o[25]) );
  OA22X1 U26982 ( .IN1(n1764), .IN2(n19244), .IN3(n1660), .IN4(n19223), .Q(
        n8167) );
  OA22X1 U26983 ( .IN1(n1936), .IN2(n19277), .IN3(n1850), .IN4(n19256), .Q(
        n8168) );
  OA22X1 U26984 ( .IN1(n2108), .IN2(n19310), .IN3(n2022), .IN4(n19289), .Q(
        n8169) );
  NAND4X0 U26985 ( .IN1(n8163), .IN2(n8164), .IN3(n8165), .IN4(n8166), .QN(
        s12_addr_o[26]) );
  OA22X1 U26986 ( .IN1(n1763), .IN2(n19243), .IN3(n1659), .IN4(n19224), .Q(
        n8163) );
  OA22X1 U26987 ( .IN1(n1935), .IN2(n19276), .IN3(n1849), .IN4(n19257), .Q(
        n8164) );
  OA22X1 U26988 ( .IN1(n2107), .IN2(n19309), .IN3(n2021), .IN4(n19290), .Q(
        n8165) );
  NAND4X0 U26989 ( .IN1(n8159), .IN2(n8160), .IN3(n8161), .IN4(n8162), .QN(
        s12_addr_o[27]) );
  OA22X1 U26990 ( .IN1(n1762), .IN2(n19242), .IN3(n1658), .IN4(n19224), .Q(
        n8159) );
  OA22X1 U26991 ( .IN1(n1934), .IN2(n19275), .IN3(n1848), .IN4(n19257), .Q(
        n8160) );
  OA22X1 U26992 ( .IN1(n2106), .IN2(n19308), .IN3(n2020), .IN4(n19290), .Q(
        n8161) );
  NAND4X0 U26993 ( .IN1(n8155), .IN2(n8156), .IN3(n8157), .IN4(n8158), .QN(
        s12_addr_o[28]) );
  OA22X1 U26994 ( .IN1(n1761), .IN2(n19242), .IN3(n1657), .IN4(n19224), .Q(
        n8155) );
  OA22X1 U26995 ( .IN1(n1933), .IN2(n19275), .IN3(n1847), .IN4(n19257), .Q(
        n8156) );
  OA22X1 U26996 ( .IN1(n2105), .IN2(n19308), .IN3(n2019), .IN4(n19290), .Q(
        n8157) );
  NAND4X0 U26997 ( .IN1(n8151), .IN2(n8152), .IN3(n8153), .IN4(n8154), .QN(
        s12_addr_o[29]) );
  OA22X1 U26998 ( .IN1(n1760), .IN2(n19246), .IN3(n1656), .IN4(n19225), .Q(
        n8151) );
  OA22X1 U26999 ( .IN1(n1932), .IN2(n19279), .IN3(n1846), .IN4(n19258), .Q(
        n8152) );
  OA22X1 U27000 ( .IN1(n2104), .IN2(n19312), .IN3(n2018), .IN4(n19291), .Q(
        n8153) );
  NAND4X0 U27001 ( .IN1(n8143), .IN2(n8144), .IN3(n8145), .IN4(n8146), .QN(
        s12_addr_o[30]) );
  OA22X1 U27002 ( .IN1(n1759), .IN2(n19247), .IN3(n1655), .IN4(n19225), .Q(
        n8143) );
  OA22X1 U27003 ( .IN1(n1931), .IN2(n19280), .IN3(n1845), .IN4(n19258), .Q(
        n8144) );
  OA22X1 U27004 ( .IN1(n2103), .IN2(n19313), .IN3(n2017), .IN4(n19291), .Q(
        n8145) );
  NAND4X0 U27005 ( .IN1(n8139), .IN2(n8140), .IN3(n8141), .IN4(n8142), .QN(
        s12_addr_o[31]) );
  OA22X1 U27006 ( .IN1(n1758), .IN2(n19245), .IN3(n1650), .IN4(n19226), .Q(
        n8139) );
  OA22X1 U27007 ( .IN1(n1930), .IN2(n19278), .IN3(n1844), .IN4(n19259), .Q(
        n8140) );
  OA22X1 U27008 ( .IN1(n2102), .IN2(n19311), .IN3(n2016), .IN4(n19292), .Q(
        n8141) );
  NAND4X0 U27009 ( .IN1(n8107), .IN2(n8108), .IN3(n8109), .IN4(n8110), .QN(
        s12_data_o[0]) );
  OA22X1 U27010 ( .IN1(n1741), .IN2(n19244), .IN3(n1636), .IN4(n19227), .Q(
        n8107) );
  OA22X1 U27011 ( .IN1(n1913), .IN2(n19277), .IN3(n1827), .IN4(n19260), .Q(
        n8108) );
  OA22X1 U27012 ( .IN1(n2085), .IN2(n19310), .IN3(n1999), .IN4(n19293), .Q(
        n8109) );
  NAND4X0 U27013 ( .IN1(n8063), .IN2(n8064), .IN3(n8065), .IN4(n8066), .QN(
        s12_data_o[1]) );
  OA22X1 U27014 ( .IN1(n1740), .IN2(n19246), .IN3(n1635), .IN4(n19225), .Q(
        n8063) );
  OA22X1 U27015 ( .IN1(n1912), .IN2(n19279), .IN3(n1826), .IN4(n19258), .Q(
        n8064) );
  OA22X1 U27016 ( .IN1(n2084), .IN2(n19312), .IN3(n1998), .IN4(n19291), .Q(
        n8065) );
  NAND4X0 U27017 ( .IN1(n8019), .IN2(n8020), .IN3(n8021), .IN4(n8022), .QN(
        s12_data_o[2]) );
  OA22X1 U27018 ( .IN1(n1739), .IN2(n19247), .IN3(n1634), .IN4(n19218), .Q(
        n8019) );
  OA22X1 U27019 ( .IN1(n1911), .IN2(n19280), .IN3(n1825), .IN4(n19251), .Q(
        n8020) );
  OA22X1 U27020 ( .IN1(n2083), .IN2(n19313), .IN3(n1997), .IN4(n19284), .Q(
        n8021) );
  NAND4X0 U27021 ( .IN1(n8007), .IN2(n8008), .IN3(n8009), .IN4(n8010), .QN(
        s12_data_o[3]) );
  OA22X1 U27022 ( .IN1(n1738), .IN2(n19245), .IN3(n1633), .IN4(n19220), .Q(
        n8007) );
  OA22X1 U27023 ( .IN1(n1910), .IN2(n19278), .IN3(n1824), .IN4(n19253), .Q(
        n8008) );
  OA22X1 U27024 ( .IN1(n2082), .IN2(n19311), .IN3(n1996), .IN4(n19286), .Q(
        n8009) );
  NAND4X0 U27025 ( .IN1(n8003), .IN2(n8004), .IN3(n8005), .IN4(n8006), .QN(
        s12_data_o[4]) );
  OA22X1 U27026 ( .IN1(n1737), .IN2(n19246), .IN3(n1632), .IN4(n19235), .Q(
        n8003) );
  OA22X1 U27027 ( .IN1(n1909), .IN2(n19279), .IN3(n1823), .IN4(n19268), .Q(
        n8004) );
  OA22X1 U27028 ( .IN1(n2081), .IN2(n19312), .IN3(n1995), .IN4(n19301), .Q(
        n8005) );
  NAND4X0 U27029 ( .IN1(n7999), .IN2(n8000), .IN3(n8001), .IN4(n8002), .QN(
        s12_data_o[5]) );
  OA22X1 U27030 ( .IN1(n1736), .IN2(n19247), .IN3(n1631), .IN4(n19233), .Q(
        n7999) );
  OA22X1 U27031 ( .IN1(n1908), .IN2(n19280), .IN3(n1822), .IN4(n19266), .Q(
        n8000) );
  OA22X1 U27032 ( .IN1(n2080), .IN2(n19313), .IN3(n1994), .IN4(n19299), .Q(
        n8001) );
  NAND4X0 U27033 ( .IN1(n7995), .IN2(n7996), .IN3(n7997), .IN4(n7998), .QN(
        s12_data_o[6]) );
  OA22X1 U27034 ( .IN1(n1735), .IN2(n19243), .IN3(n1630), .IN4(n19233), .Q(
        n7995) );
  OA22X1 U27035 ( .IN1(n1907), .IN2(n19276), .IN3(n1821), .IN4(n19266), .Q(
        n7996) );
  OA22X1 U27036 ( .IN1(n2079), .IN2(n19309), .IN3(n1993), .IN4(n19299), .Q(
        n7997) );
  NAND4X0 U27037 ( .IN1(n7991), .IN2(n7992), .IN3(n7993), .IN4(n7994), .QN(
        s12_data_o[7]) );
  OA22X1 U27038 ( .IN1(n1734), .IN2(n19241), .IN3(n1629), .IN4(n19233), .Q(
        n7991) );
  OA22X1 U27039 ( .IN1(n1906), .IN2(n19274), .IN3(n1820), .IN4(n19266), .Q(
        n7992) );
  OA22X1 U27040 ( .IN1(n2078), .IN2(n19307), .IN3(n1992), .IN4(n19299), .Q(
        n7993) );
  NAND4X0 U27041 ( .IN1(n7987), .IN2(n7988), .IN3(n7989), .IN4(n7990), .QN(
        s12_data_o[8]) );
  OA22X1 U27042 ( .IN1(n1733), .IN2(n19248), .IN3(n1628), .IN4(n19233), .Q(
        n7987) );
  OA22X1 U27043 ( .IN1(n1905), .IN2(n19281), .IN3(n1819), .IN4(n19266), .Q(
        n7988) );
  OA22X1 U27044 ( .IN1(n2077), .IN2(n19314), .IN3(n1991), .IN4(n19299), .Q(
        n7989) );
  NAND4X0 U27045 ( .IN1(n7983), .IN2(n7984), .IN3(n7985), .IN4(n7986), .QN(
        s12_data_o[9]) );
  OA22X1 U27046 ( .IN1(n1732), .IN2(n19241), .IN3(n1627), .IN4(n19234), .Q(
        n7983) );
  OA22X1 U27047 ( .IN1(n1904), .IN2(n19274), .IN3(n1818), .IN4(n19267), .Q(
        n7984) );
  OA22X1 U27048 ( .IN1(n2076), .IN2(n19307), .IN3(n1990), .IN4(n19300), .Q(
        n7985) );
  NAND4X0 U27049 ( .IN1(n8103), .IN2(n8104), .IN3(n8105), .IN4(n8106), .QN(
        s12_data_o[10]) );
  OA22X1 U27050 ( .IN1(n1731), .IN2(n19243), .IN3(n1626), .IN4(n19228), .Q(
        n8103) );
  OA22X1 U27051 ( .IN1(n1903), .IN2(n19276), .IN3(n1817), .IN4(n19261), .Q(
        n8104) );
  OA22X1 U27052 ( .IN1(n2075), .IN2(n19309), .IN3(n1989), .IN4(n19294), .Q(
        n8105) );
  NAND4X0 U27053 ( .IN1(n8099), .IN2(n8100), .IN3(n8101), .IN4(n8102), .QN(
        s12_data_o[11]) );
  OA22X1 U27054 ( .IN1(n1730), .IN2(n19248), .IN3(n1625), .IN4(n19228), .Q(
        n8099) );
  OA22X1 U27055 ( .IN1(n1902), .IN2(n19281), .IN3(n1816), .IN4(n19261), .Q(
        n8100) );
  OA22X1 U27056 ( .IN1(n2074), .IN2(n19314), .IN3(n1988), .IN4(n19294), .Q(
        n8101) );
  NAND4X0 U27057 ( .IN1(n8095), .IN2(n8096), .IN3(n8097), .IN4(n8098), .QN(
        s12_data_o[12]) );
  OA22X1 U27058 ( .IN1(n1729), .IN2(n19244), .IN3(n1624), .IN4(n19228), .Q(
        n8095) );
  OA22X1 U27059 ( .IN1(n1901), .IN2(n19277), .IN3(n1815), .IN4(n19261), .Q(
        n8096) );
  OA22X1 U27060 ( .IN1(n2073), .IN2(n19310), .IN3(n1987), .IN4(n19294), .Q(
        n8097) );
  NAND4X0 U27061 ( .IN1(n8091), .IN2(n8092), .IN3(n8093), .IN4(n8094), .QN(
        s12_data_o[13]) );
  OA22X1 U27062 ( .IN1(n1728), .IN2(n19245), .IN3(n1623), .IN4(n19222), .Q(
        n8091) );
  OA22X1 U27063 ( .IN1(n1900), .IN2(n19278), .IN3(n1814), .IN4(n19255), .Q(
        n8092) );
  OA22X1 U27064 ( .IN1(n2072), .IN2(n19311), .IN3(n1986), .IN4(n19288), .Q(
        n8093) );
  NAND4X0 U27065 ( .IN1(n8087), .IN2(n8088), .IN3(n8089), .IN4(n8090), .QN(
        s12_data_o[14]) );
  OA22X1 U27066 ( .IN1(n1727), .IN2(n19245), .IN3(n1622), .IN4(n19227), .Q(
        n8087) );
  OA22X1 U27067 ( .IN1(n1899), .IN2(n19278), .IN3(n1813), .IN4(n19260), .Q(
        n8088) );
  OA22X1 U27068 ( .IN1(n2071), .IN2(n19311), .IN3(n1985), .IN4(n19293), .Q(
        n8089) );
  NAND4X0 U27069 ( .IN1(n8083), .IN2(n8084), .IN3(n8085), .IN4(n8086), .QN(
        s12_data_o[15]) );
  OA22X1 U27070 ( .IN1(n1726), .IN2(n19245), .IN3(n1621), .IN4(n19228), .Q(
        n8083) );
  OA22X1 U27071 ( .IN1(n1898), .IN2(n19278), .IN3(n1812), .IN4(n19261), .Q(
        n8084) );
  OA22X1 U27072 ( .IN1(n2070), .IN2(n19311), .IN3(n1984), .IN4(n19294), .Q(
        n8085) );
  NAND4X0 U27073 ( .IN1(n8079), .IN2(n8080), .IN3(n8081), .IN4(n8082), .QN(
        s12_data_o[16]) );
  OA22X1 U27074 ( .IN1(n1725), .IN2(n19245), .IN3(n1620), .IN4(n19229), .Q(
        n8079) );
  OA22X1 U27075 ( .IN1(n1897), .IN2(n19278), .IN3(n1811), .IN4(n19262), .Q(
        n8080) );
  OA22X1 U27076 ( .IN1(n2069), .IN2(n19311), .IN3(n1983), .IN4(n19295), .Q(
        n8081) );
  NAND4X0 U27077 ( .IN1(n8075), .IN2(n8076), .IN3(n8077), .IN4(n8078), .QN(
        s12_data_o[17]) );
  OA22X1 U27078 ( .IN1(n1724), .IN2(n19246), .IN3(n1619), .IN4(n19229), .Q(
        n8075) );
  OA22X1 U27079 ( .IN1(n1896), .IN2(n19279), .IN3(n1810), .IN4(n19262), .Q(
        n8076) );
  OA22X1 U27080 ( .IN1(n2068), .IN2(n19312), .IN3(n1982), .IN4(n19295), .Q(
        n8077) );
  NAND4X0 U27081 ( .IN1(n8071), .IN2(n8072), .IN3(n8073), .IN4(n8074), .QN(
        s12_data_o[18]) );
  OA22X1 U27082 ( .IN1(n1723), .IN2(n19246), .IN3(n1618), .IN4(n19229), .Q(
        n8071) );
  OA22X1 U27083 ( .IN1(n1895), .IN2(n19279), .IN3(n1809), .IN4(n19262), .Q(
        n8072) );
  OA22X1 U27084 ( .IN1(n2067), .IN2(n19312), .IN3(n1981), .IN4(n19295), .Q(
        n8073) );
  NAND4X0 U27085 ( .IN1(n8067), .IN2(n8068), .IN3(n8069), .IN4(n8070), .QN(
        s12_data_o[19]) );
  OA22X1 U27086 ( .IN1(n1722), .IN2(n19246), .IN3(n1617), .IN4(n19229), .Q(
        n8067) );
  OA22X1 U27087 ( .IN1(n1894), .IN2(n19279), .IN3(n1808), .IN4(n19262), .Q(
        n8068) );
  OA22X1 U27088 ( .IN1(n2066), .IN2(n19312), .IN3(n1980), .IN4(n19295), .Q(
        n8069) );
  NAND4X0 U27089 ( .IN1(n8059), .IN2(n8060), .IN3(n8061), .IN4(n8062), .QN(
        s12_data_o[20]) );
  OA22X1 U27090 ( .IN1(n1721), .IN2(n19247), .IN3(n1616), .IN4(n19226), .Q(
        n8059) );
  OA22X1 U27091 ( .IN1(n1893), .IN2(n19280), .IN3(n1807), .IN4(n19259), .Q(
        n8060) );
  OA22X1 U27092 ( .IN1(n2065), .IN2(n19313), .IN3(n1979), .IN4(n19292), .Q(
        n8061) );
  NAND4X0 U27093 ( .IN1(n8055), .IN2(n8056), .IN3(n8057), .IN4(n8058), .QN(
        s12_data_o[21]) );
  OA22X1 U27094 ( .IN1(n1720), .IN2(n19247), .IN3(n1615), .IN4(n19230), .Q(
        n8055) );
  OA22X1 U27095 ( .IN1(n1892), .IN2(n19280), .IN3(n1806), .IN4(n19263), .Q(
        n8056) );
  OA22X1 U27096 ( .IN1(n2064), .IN2(n19313), .IN3(n1978), .IN4(n19296), .Q(
        n8057) );
  NAND4X0 U27097 ( .IN1(n8051), .IN2(n8052), .IN3(n8053), .IN4(n8054), .QN(
        s12_data_o[22]) );
  OA22X1 U27098 ( .IN1(n1719), .IN2(n19245), .IN3(n1614), .IN4(n19230), .Q(
        n8051) );
  OA22X1 U27099 ( .IN1(n1891), .IN2(n19278), .IN3(n1805), .IN4(n19263), .Q(
        n8052) );
  OA22X1 U27100 ( .IN1(n2063), .IN2(n19311), .IN3(n1977), .IN4(n19296), .Q(
        n8053) );
  NAND4X0 U27101 ( .IN1(n8047), .IN2(n8048), .IN3(n8049), .IN4(n8050), .QN(
        s12_data_o[23]) );
  OA22X1 U27102 ( .IN1(n1718), .IN2(n19246), .IN3(n1613), .IN4(n19230), .Q(
        n8047) );
  OA22X1 U27103 ( .IN1(n1890), .IN2(n19279), .IN3(n1804), .IN4(n19263), .Q(
        n8048) );
  OA22X1 U27104 ( .IN1(n2062), .IN2(n19312), .IN3(n1976), .IN4(n19296), .Q(
        n8049) );
  NAND4X0 U27105 ( .IN1(n8043), .IN2(n8044), .IN3(n8045), .IN4(n8046), .QN(
        s12_data_o[24]) );
  OA22X1 U27106 ( .IN1(n1717), .IN2(n19244), .IN3(n1612), .IN4(n19231), .Q(
        n8043) );
  OA22X1 U27107 ( .IN1(n1889), .IN2(n19277), .IN3(n1803), .IN4(n19264), .Q(
        n8044) );
  OA22X1 U27108 ( .IN1(n2061), .IN2(n19310), .IN3(n1975), .IN4(n19297), .Q(
        n8045) );
  NAND4X0 U27109 ( .IN1(n8039), .IN2(n8040), .IN3(n8041), .IN4(n8042), .QN(
        s12_data_o[25]) );
  OA22X1 U27110 ( .IN1(n1716), .IN2(n19244), .IN3(n1611), .IN4(n19231), .Q(
        n8039) );
  OA22X1 U27111 ( .IN1(n1888), .IN2(n19277), .IN3(n1802), .IN4(n19264), .Q(
        n8040) );
  OA22X1 U27112 ( .IN1(n2060), .IN2(n19310), .IN3(n1974), .IN4(n19297), .Q(
        n8041) );
  NAND4X0 U27113 ( .IN1(n8035), .IN2(n8036), .IN3(n8037), .IN4(n8038), .QN(
        s12_data_o[26]) );
  OA22X1 U27114 ( .IN1(n1715), .IN2(n19243), .IN3(n1610), .IN4(n19231), .Q(
        n8035) );
  OA22X1 U27115 ( .IN1(n1887), .IN2(n19276), .IN3(n1801), .IN4(n19264), .Q(
        n8036) );
  OA22X1 U27116 ( .IN1(n2059), .IN2(n19309), .IN3(n1973), .IN4(n19297), .Q(
        n8037) );
  NAND4X0 U27117 ( .IN1(n8031), .IN2(n8032), .IN3(n8033), .IN4(n8034), .QN(
        s12_data_o[27]) );
  OA22X1 U27118 ( .IN1(n1714), .IN2(n19246), .IN3(n1609), .IN4(n19232), .Q(
        n8031) );
  OA22X1 U27119 ( .IN1(n1886), .IN2(n19279), .IN3(n1800), .IN4(n19265), .Q(
        n8032) );
  OA22X1 U27120 ( .IN1(n2058), .IN2(n19312), .IN3(n1972), .IN4(n19298), .Q(
        n8033) );
  NAND4X0 U27121 ( .IN1(n8027), .IN2(n8028), .IN3(n8029), .IN4(n8030), .QN(
        s12_data_o[28]) );
  OA22X1 U27122 ( .IN1(n1713), .IN2(n19247), .IN3(n1608), .IN4(n19232), .Q(
        n8027) );
  OA22X1 U27123 ( .IN1(n1885), .IN2(n19280), .IN3(n1799), .IN4(n19265), .Q(
        n8028) );
  OA22X1 U27124 ( .IN1(n2057), .IN2(n19313), .IN3(n1971), .IN4(n19298), .Q(
        n8029) );
  NAND4X0 U27125 ( .IN1(n8023), .IN2(n8024), .IN3(n8025), .IN4(n8026), .QN(
        s12_data_o[29]) );
  OA22X1 U27126 ( .IN1(n1712), .IN2(n19247), .IN3(n1607), .IN4(n19232), .Q(
        n8023) );
  OA22X1 U27127 ( .IN1(n1884), .IN2(n19280), .IN3(n1798), .IN4(n19265), .Q(
        n8024) );
  OA22X1 U27128 ( .IN1(n2056), .IN2(n19313), .IN3(n1970), .IN4(n19298), .Q(
        n8025) );
  NAND4X0 U27129 ( .IN1(n8015), .IN2(n8016), .IN3(n8017), .IN4(n8018), .QN(
        s12_data_o[30]) );
  OA22X1 U27130 ( .IN1(n1711), .IN2(n19247), .IN3(n1606), .IN4(n19234), .Q(
        n8015) );
  OA22X1 U27131 ( .IN1(n1883), .IN2(n19280), .IN3(n1797), .IN4(n19267), .Q(
        n8016) );
  OA22X1 U27132 ( .IN1(n2055), .IN2(n19313), .IN3(n1969), .IN4(n19300), .Q(
        n8017) );
  NAND4X0 U27133 ( .IN1(n8011), .IN2(n8012), .IN3(n8013), .IN4(n8014), .QN(
        s12_data_o[31]) );
  OA22X1 U27134 ( .IN1(n1710), .IN2(n19245), .IN3(n1605), .IN4(n19219), .Q(
        n8011) );
  OA22X1 U27135 ( .IN1(n1882), .IN2(n19278), .IN3(n1796), .IN4(n19252), .Q(
        n8012) );
  OA22X1 U27136 ( .IN1(n2054), .IN2(n19311), .IN3(n1968), .IN4(n19285), .Q(
        n8013) );
  NAND4X0 U27137 ( .IN1(n8251), .IN2(n8252), .IN3(n8253), .IN4(n8254), .QN(
        s11_stb_o) );
  OA22X1 U27138 ( .IN1(n1795), .IN2(n8261), .IN3(n1709), .IN4(n8262), .Q(n8251) );
  OA22X1 U27139 ( .IN1(n1967), .IN2(n8259), .IN3(n1881), .IN4(n8260), .Q(n8252) );
  OA22X1 U27140 ( .IN1(n2139), .IN2(n8257), .IN3(n2053), .IN4(n8258), .Q(n8253) );
  NAND4X0 U27141 ( .IN1(n8239), .IN2(n8240), .IN3(n8241), .IN4(n8242), .QN(
        s11_we_o) );
  OA22X1 U27142 ( .IN1(n1794), .IN2(n19109), .IN3(n1708), .IN4(n19103), .Q(
        n8239) );
  OA22X1 U27143 ( .IN1(n1966), .IN2(n19142), .IN3(n1880), .IN4(n19136), .Q(
        n8240) );
  OA22X1 U27144 ( .IN1(n2138), .IN2(n19182), .IN3(n2052), .IN4(n19169), .Q(
        n8241) );
  NAND4X0 U27145 ( .IN1(n8275), .IN2(n8276), .IN3(n8277), .IN4(n8278), .QN(
        s11_sel_o[0]) );
  OA22X1 U27146 ( .IN1(n1793), .IN2(n19116), .IN3(n1707), .IN4(n19102), .Q(
        n8275) );
  OA22X1 U27147 ( .IN1(n1965), .IN2(n19149), .IN3(n1879), .IN4(n19135), .Q(
        n8276) );
  OA22X1 U27148 ( .IN1(n2137), .IN2(n19182), .IN3(n2051), .IN4(n19167), .Q(
        n8277) );
  NAND4X0 U27149 ( .IN1(n8271), .IN2(n8272), .IN3(n8273), .IN4(n8274), .QN(
        s11_sel_o[1]) );
  OA22X1 U27150 ( .IN1(n1792), .IN2(n19116), .IN3(n1706), .IN4(n19102), .Q(
        n8271) );
  OA22X1 U27151 ( .IN1(n1964), .IN2(n19149), .IN3(n1878), .IN4(n19135), .Q(
        n8272) );
  OA22X1 U27152 ( .IN1(n2136), .IN2(n19182), .IN3(n2050), .IN4(n19167), .Q(
        n8273) );
  NAND4X0 U27153 ( .IN1(n8267), .IN2(n8268), .IN3(n8269), .IN4(n8270), .QN(
        s11_sel_o[2]) );
  OA22X1 U27154 ( .IN1(n1791), .IN2(n19116), .IN3(n1705), .IN4(n19103), .Q(
        n8267) );
  OA22X1 U27155 ( .IN1(n1963), .IN2(n19149), .IN3(n1877), .IN4(n19136), .Q(
        n8268) );
  OA22X1 U27156 ( .IN1(n2135), .IN2(n19182), .IN3(n2049), .IN4(n19169), .Q(
        n8269) );
  NAND4X0 U27157 ( .IN1(n8263), .IN2(n8264), .IN3(n8265), .IN4(n8266), .QN(
        s11_sel_o[3]) );
  OA22X1 U27158 ( .IN1(n1790), .IN2(n19116), .IN3(n1704), .IN4(n19103), .Q(
        n8263) );
  OA22X1 U27159 ( .IN1(n1962), .IN2(n19149), .IN3(n1876), .IN4(n19136), .Q(
        n8264) );
  OA22X1 U27160 ( .IN1(n2134), .IN2(n19182), .IN3(n2048), .IN4(n19169), .Q(
        n8265) );
  NAND4X0 U27161 ( .IN1(n8531), .IN2(n8532), .IN3(n8533), .IN4(n8534), .QN(
        s11_addr_o[0]) );
  OA22X1 U27162 ( .IN1(n1789), .IN2(n19109), .IN3(n1703), .IN4(n19086), .Q(
        n8531) );
  OA22X1 U27163 ( .IN1(n1961), .IN2(n19142), .IN3(n1875), .IN4(n19119), .Q(
        n8532) );
  OA22X1 U27164 ( .IN1(n2133), .IN2(n19177), .IN3(n2047), .IN4(n19152), .Q(
        n8533) );
  NAND4X0 U27165 ( .IN1(n8487), .IN2(n8488), .IN3(n8489), .IN4(n8490), .QN(
        s11_addr_o[1]) );
  OA22X1 U27166 ( .IN1(n1788), .IN2(n19111), .IN3(n1702), .IN4(n19089), .Q(
        n8487) );
  OA22X1 U27167 ( .IN1(n1960), .IN2(n19144), .IN3(n1874), .IN4(n19122), .Q(
        n8488) );
  OA22X1 U27168 ( .IN1(n2132), .IN2(n19176), .IN3(n2046), .IN4(n19155), .Q(
        n8489) );
  NAND4X0 U27169 ( .IN1(n8443), .IN2(n8444), .IN3(n8445), .IN4(n8446), .QN(
        s11_addr_o[2]) );
  OA22X1 U27170 ( .IN1(n1787), .IN2(n19111), .IN3(n1701), .IN4(n19093), .Q(
        n8443) );
  OA22X1 U27171 ( .IN1(n1959), .IN2(n19144), .IN3(n1873), .IN4(n19126), .Q(
        n8444) );
  OA22X1 U27172 ( .IN1(n2131), .IN2(n19176), .IN3(n2045), .IN4(n19159), .Q(
        n8445) );
  NAND4X0 U27173 ( .IN1(n8431), .IN2(n8432), .IN3(n8433), .IN4(n8434), .QN(
        s11_addr_o[3]) );
  OA22X1 U27174 ( .IN1(n1786), .IN2(n19116), .IN3(n1699), .IN4(n19094), .Q(
        n8431) );
  OA22X1 U27175 ( .IN1(n1958), .IN2(n19149), .IN3(n1872), .IN4(n19127), .Q(
        n8432) );
  OA22X1 U27176 ( .IN1(n2130), .IN2(n19182), .IN3(n2044), .IN4(n19160), .Q(
        n8433) );
  NAND4X0 U27177 ( .IN1(n8427), .IN2(n8428), .IN3(n8429), .IN4(n8430), .QN(
        s11_addr_o[4]) );
  OA22X1 U27178 ( .IN1(n1785), .IN2(n19109), .IN3(n1697), .IN4(n19094), .Q(
        n8427) );
  OA22X1 U27179 ( .IN1(n1957), .IN2(n19142), .IN3(n1871), .IN4(n19127), .Q(
        n8428) );
  OA22X1 U27180 ( .IN1(n2129), .IN2(n19177), .IN3(n2043), .IN4(n19160), .Q(
        n8429) );
  NAND4X0 U27181 ( .IN1(n8423), .IN2(n8424), .IN3(n8425), .IN4(n8426), .QN(
        s11_addr_o[5]) );
  OA22X1 U27182 ( .IN1(n1784), .IN2(n19116), .IN3(n1696), .IN4(n19093), .Q(
        n8423) );
  OA22X1 U27183 ( .IN1(n1956), .IN2(n19149), .IN3(n1870), .IN4(n19126), .Q(
        n8424) );
  OA22X1 U27184 ( .IN1(n2128), .IN2(n19182), .IN3(n2042), .IN4(n19161), .Q(
        n8425) );
  NAND4X0 U27185 ( .IN1(n8419), .IN2(n8420), .IN3(n8421), .IN4(n8422), .QN(
        s11_addr_o[6]) );
  OA22X1 U27186 ( .IN1(n1783), .IN2(n19112), .IN3(n1679), .IN4(n19094), .Q(
        n8419) );
  OA22X1 U27187 ( .IN1(n1955), .IN2(n19145), .IN3(n1869), .IN4(n19127), .Q(
        n8420) );
  OA22X1 U27188 ( .IN1(n2127), .IN2(n19178), .IN3(n2041), .IN4(n19161), .Q(
        n8421) );
  NAND4X0 U27189 ( .IN1(n8415), .IN2(n8416), .IN3(n8417), .IN4(n8418), .QN(
        s11_addr_o[7]) );
  OA22X1 U27190 ( .IN1(n1782), .IN2(n19112), .IN3(n1678), .IN4(n19086), .Q(
        n8415) );
  OA22X1 U27191 ( .IN1(n1954), .IN2(n19145), .IN3(n1868), .IN4(n19119), .Q(
        n8416) );
  OA22X1 U27192 ( .IN1(n2126), .IN2(n19178), .IN3(n2040), .IN4(n19161), .Q(
        n8417) );
  NAND4X0 U27193 ( .IN1(n8411), .IN2(n8412), .IN3(n8413), .IN4(n8414), .QN(
        s11_addr_o[8]) );
  OA22X1 U27194 ( .IN1(n1781), .IN2(n19112), .IN3(n1677), .IN4(n19095), .Q(
        n8411) );
  OA22X1 U27195 ( .IN1(n1953), .IN2(n19145), .IN3(n1867), .IN4(n19128), .Q(
        n8412) );
  OA22X1 U27196 ( .IN1(n2125), .IN2(n19178), .IN3(n2039), .IN4(n19162), .Q(
        n8413) );
  NAND4X0 U27197 ( .IN1(n8407), .IN2(n8408), .IN3(n8409), .IN4(n8410), .QN(
        s11_addr_o[9]) );
  OA22X1 U27198 ( .IN1(n1780), .IN2(n19112), .IN3(n1676), .IN4(n19095), .Q(
        n8407) );
  OA22X1 U27199 ( .IN1(n1952), .IN2(n19145), .IN3(n1866), .IN4(n19128), .Q(
        n8408) );
  OA22X1 U27200 ( .IN1(n2124), .IN2(n19178), .IN3(n2038), .IN4(n19162), .Q(
        n8409) );
  NAND4X0 U27201 ( .IN1(n8527), .IN2(n8528), .IN3(n8529), .IN4(n8530), .QN(
        s11_addr_o[10]) );
  OA22X1 U27202 ( .IN1(n1779), .IN2(n19109), .IN3(n1675), .IN4(n19086), .Q(
        n8527) );
  OA22X1 U27203 ( .IN1(n1951), .IN2(n19142), .IN3(n1865), .IN4(n19119), .Q(
        n8528) );
  OA22X1 U27204 ( .IN1(n2123), .IN2(n8245), .IN3(n2037), .IN4(n19152), .Q(
        n8529) );
  NAND4X0 U27205 ( .IN1(n8523), .IN2(n8524), .IN3(n8525), .IN4(n8526), .QN(
        s11_addr_o[11]) );
  OA22X1 U27206 ( .IN1(n1778), .IN2(n19109), .IN3(n1674), .IN4(n19086), .Q(
        n8523) );
  OA22X1 U27207 ( .IN1(n1950), .IN2(n19142), .IN3(n1864), .IN4(n19119), .Q(
        n8524) );
  OA22X1 U27208 ( .IN1(n2122), .IN2(n8245), .IN3(n2036), .IN4(n19152), .Q(
        n8525) );
  NAND4X0 U27209 ( .IN1(n8519), .IN2(n8520), .IN3(n8521), .IN4(n8522), .QN(
        s11_addr_o[12]) );
  OA22X1 U27210 ( .IN1(n1777), .IN2(n19109), .IN3(n1673), .IN4(n19087), .Q(
        n8519) );
  OA22X1 U27211 ( .IN1(n1949), .IN2(n19142), .IN3(n1863), .IN4(n19120), .Q(
        n8520) );
  OA22X1 U27212 ( .IN1(n2121), .IN2(n8245), .IN3(n2035), .IN4(n19153), .Q(
        n8521) );
  NAND4X0 U27213 ( .IN1(n8515), .IN2(n8516), .IN3(n8517), .IN4(n8518), .QN(
        s11_addr_o[13]) );
  OA22X1 U27214 ( .IN1(n1776), .IN2(n19110), .IN3(n1672), .IN4(n19087), .Q(
        n8515) );
  OA22X1 U27215 ( .IN1(n1948), .IN2(n19143), .IN3(n1862), .IN4(n19120), .Q(
        n8516) );
  OA22X1 U27216 ( .IN1(n2120), .IN2(n19175), .IN3(n2034), .IN4(n19153), .Q(
        n8517) );
  NAND4X0 U27217 ( .IN1(n8511), .IN2(n8512), .IN3(n8513), .IN4(n8514), .QN(
        s11_addr_o[14]) );
  OA22X1 U27218 ( .IN1(n1775), .IN2(n19110), .IN3(n1671), .IN4(n19087), .Q(
        n8511) );
  OA22X1 U27219 ( .IN1(n1947), .IN2(n19143), .IN3(n1861), .IN4(n19120), .Q(
        n8512) );
  OA22X1 U27220 ( .IN1(n2119), .IN2(n19175), .IN3(n2033), .IN4(n19153), .Q(
        n8513) );
  NAND4X0 U27221 ( .IN1(n8507), .IN2(n8508), .IN3(n8509), .IN4(n8510), .QN(
        s11_addr_o[15]) );
  OA22X1 U27222 ( .IN1(n1774), .IN2(n19110), .IN3(n1670), .IN4(n19088), .Q(
        n8507) );
  OA22X1 U27223 ( .IN1(n1946), .IN2(n19143), .IN3(n1860), .IN4(n19121), .Q(
        n8508) );
  OA22X1 U27224 ( .IN1(n2118), .IN2(n19175), .IN3(n2032), .IN4(n19154), .Q(
        n8509) );
  NAND4X0 U27225 ( .IN1(n8503), .IN2(n8504), .IN3(n8505), .IN4(n8506), .QN(
        s11_addr_o[16]) );
  OA22X1 U27226 ( .IN1(n1773), .IN2(n19110), .IN3(n1669), .IN4(n19088), .Q(
        n8503) );
  OA22X1 U27227 ( .IN1(n1945), .IN2(n19143), .IN3(n1859), .IN4(n19121), .Q(
        n8504) );
  OA22X1 U27228 ( .IN1(n2117), .IN2(n19175), .IN3(n2031), .IN4(n19154), .Q(
        n8505) );
  NAND4X0 U27229 ( .IN1(n8499), .IN2(n8500), .IN3(n8501), .IN4(n8502), .QN(
        s11_addr_o[17]) );
  OA22X1 U27230 ( .IN1(n1772), .IN2(n19111), .IN3(n1668), .IN4(n19088), .Q(
        n8499) );
  OA22X1 U27231 ( .IN1(n1944), .IN2(n19144), .IN3(n1858), .IN4(n19121), .Q(
        n8500) );
  OA22X1 U27232 ( .IN1(n2116), .IN2(n19176), .IN3(n2030), .IN4(n19154), .Q(
        n8501) );
  NAND4X0 U27233 ( .IN1(n8495), .IN2(n8496), .IN3(n8497), .IN4(n8498), .QN(
        s11_addr_o[18]) );
  OA22X1 U27234 ( .IN1(n1771), .IN2(n19111), .IN3(n1667), .IN4(n19089), .Q(
        n8495) );
  OA22X1 U27235 ( .IN1(n1943), .IN2(n19144), .IN3(n1857), .IN4(n19122), .Q(
        n8496) );
  OA22X1 U27236 ( .IN1(n2115), .IN2(n19176), .IN3(n2029), .IN4(n19155), .Q(
        n8497) );
  NAND4X0 U27237 ( .IN1(n8491), .IN2(n8492), .IN3(n8493), .IN4(n8494), .QN(
        s11_addr_o[19]) );
  OA22X1 U27238 ( .IN1(n1770), .IN2(n19111), .IN3(n1666), .IN4(n19089), .Q(
        n8491) );
  OA22X1 U27239 ( .IN1(n1942), .IN2(n19144), .IN3(n1856), .IN4(n19122), .Q(
        n8492) );
  OA22X1 U27240 ( .IN1(n2114), .IN2(n19176), .IN3(n2028), .IN4(n19155), .Q(
        n8493) );
  NAND4X0 U27241 ( .IN1(n8483), .IN2(n8484), .IN3(n8485), .IN4(n8486), .QN(
        s11_addr_o[20]) );
  OA22X1 U27242 ( .IN1(n1769), .IN2(n19110), .IN3(n1665), .IN4(n19090), .Q(
        n8483) );
  OA22X1 U27243 ( .IN1(n1941), .IN2(n19143), .IN3(n1855), .IN4(n19123), .Q(
        n8484) );
  OA22X1 U27244 ( .IN1(n2113), .IN2(n19175), .IN3(n2027), .IN4(n19156), .Q(
        n8485) );
  NAND4X0 U27245 ( .IN1(n8479), .IN2(n8480), .IN3(n8481), .IN4(n8482), .QN(
        s11_addr_o[21]) );
  OA22X1 U27246 ( .IN1(n1768), .IN2(n19110), .IN3(n1664), .IN4(n19090), .Q(
        n8479) );
  OA22X1 U27247 ( .IN1(n1940), .IN2(n19143), .IN3(n1854), .IN4(n19123), .Q(
        n8480) );
  OA22X1 U27248 ( .IN1(n2112), .IN2(n19175), .IN3(n2026), .IN4(n19156), .Q(
        n8481) );
  NAND4X0 U27249 ( .IN1(n8475), .IN2(n8476), .IN3(n8477), .IN4(n8478), .QN(
        s11_addr_o[22]) );
  OA22X1 U27250 ( .IN1(n1767), .IN2(n19109), .IN3(n1663), .IN4(n19090), .Q(
        n8475) );
  OA22X1 U27251 ( .IN1(n1939), .IN2(n19142), .IN3(n1853), .IN4(n19123), .Q(
        n8476) );
  OA22X1 U27252 ( .IN1(n2111), .IN2(n19177), .IN3(n2025), .IN4(n19156), .Q(
        n8477) );
  NAND4X0 U27253 ( .IN1(n8471), .IN2(n8472), .IN3(n8473), .IN4(n8474), .QN(
        s11_addr_o[23]) );
  OA22X1 U27254 ( .IN1(n1766), .IN2(n19110), .IN3(n1662), .IN4(n19091), .Q(
        n8471) );
  OA22X1 U27255 ( .IN1(n1938), .IN2(n19143), .IN3(n1852), .IN4(n19124), .Q(
        n8472) );
  OA22X1 U27256 ( .IN1(n2110), .IN2(n19175), .IN3(n2024), .IN4(n19157), .Q(
        n8473) );
  NAND4X0 U27257 ( .IN1(n8467), .IN2(n8468), .IN3(n8469), .IN4(n8470), .QN(
        s11_addr_o[24]) );
  OA22X1 U27258 ( .IN1(n1765), .IN2(n19116), .IN3(n1661), .IN4(n19091), .Q(
        n8467) );
  OA22X1 U27259 ( .IN1(n1937), .IN2(n19149), .IN3(n1851), .IN4(n19124), .Q(
        n8468) );
  OA22X1 U27260 ( .IN1(n2109), .IN2(n19177), .IN3(n2023), .IN4(n19157), .Q(
        n8469) );
  NAND4X0 U27261 ( .IN1(n8463), .IN2(n8464), .IN3(n8465), .IN4(n8466), .QN(
        s11_addr_o[25]) );
  OA22X1 U27262 ( .IN1(n1764), .IN2(n19112), .IN3(n1660), .IN4(n19091), .Q(
        n8463) );
  OA22X1 U27263 ( .IN1(n1936), .IN2(n19145), .IN3(n1850), .IN4(n19124), .Q(
        n8464) );
  OA22X1 U27264 ( .IN1(n2108), .IN2(n19177), .IN3(n2022), .IN4(n19157), .Q(
        n8465) );
  NAND4X0 U27265 ( .IN1(n8459), .IN2(n8460), .IN3(n8461), .IN4(n8462), .QN(
        s11_addr_o[26]) );
  OA22X1 U27266 ( .IN1(n1763), .IN2(n19111), .IN3(n1659), .IN4(n19092), .Q(
        n8459) );
  OA22X1 U27267 ( .IN1(n1935), .IN2(n19144), .IN3(n1849), .IN4(n19125), .Q(
        n8460) );
  OA22X1 U27268 ( .IN1(n2107), .IN2(n19177), .IN3(n2021), .IN4(n19158), .Q(
        n8461) );
  NAND4X0 U27269 ( .IN1(n8455), .IN2(n8456), .IN3(n8457), .IN4(n8458), .QN(
        s11_addr_o[27]) );
  OA22X1 U27270 ( .IN1(n1762), .IN2(n19110), .IN3(n1658), .IN4(n19092), .Q(
        n8455) );
  OA22X1 U27271 ( .IN1(n1934), .IN2(n19143), .IN3(n1848), .IN4(n19125), .Q(
        n8456) );
  OA22X1 U27272 ( .IN1(n2106), .IN2(n19177), .IN3(n2020), .IN4(n19158), .Q(
        n8457) );
  NAND4X0 U27273 ( .IN1(n8451), .IN2(n8452), .IN3(n8453), .IN4(n8454), .QN(
        s11_addr_o[28]) );
  OA22X1 U27274 ( .IN1(n1761), .IN2(n19110), .IN3(n1657), .IN4(n19092), .Q(
        n8451) );
  OA22X1 U27275 ( .IN1(n1933), .IN2(n19143), .IN3(n1847), .IN4(n19125), .Q(
        n8452) );
  OA22X1 U27276 ( .IN1(n2105), .IN2(n19175), .IN3(n2019), .IN4(n19158), .Q(
        n8453) );
  NAND4X0 U27277 ( .IN1(n8447), .IN2(n8448), .IN3(n8449), .IN4(n8450), .QN(
        s11_addr_o[29]) );
  OA22X1 U27278 ( .IN1(n1760), .IN2(n19114), .IN3(n1656), .IN4(n19093), .Q(
        n8447) );
  OA22X1 U27279 ( .IN1(n1932), .IN2(n19147), .IN3(n1846), .IN4(n19126), .Q(
        n8448) );
  OA22X1 U27280 ( .IN1(n2104), .IN2(n19180), .IN3(n2018), .IN4(n19159), .Q(
        n8449) );
  NAND4X0 U27281 ( .IN1(n8439), .IN2(n8440), .IN3(n8441), .IN4(n8442), .QN(
        s11_addr_o[30]) );
  OA22X1 U27282 ( .IN1(n1759), .IN2(n19115), .IN3(n1655), .IN4(n19093), .Q(
        n8439) );
  OA22X1 U27283 ( .IN1(n1931), .IN2(n19148), .IN3(n1845), .IN4(n19126), .Q(
        n8440) );
  OA22X1 U27284 ( .IN1(n2103), .IN2(n19181), .IN3(n2017), .IN4(n19159), .Q(
        n8441) );
  NAND4X0 U27285 ( .IN1(n8435), .IN2(n8436), .IN3(n8437), .IN4(n8438), .QN(
        s11_addr_o[31]) );
  OA22X1 U27286 ( .IN1(n1758), .IN2(n19113), .IN3(n1650), .IN4(n19094), .Q(
        n8435) );
  OA22X1 U27287 ( .IN1(n1930), .IN2(n19146), .IN3(n1844), .IN4(n19127), .Q(
        n8436) );
  OA22X1 U27288 ( .IN1(n2102), .IN2(n19179), .IN3(n2016), .IN4(n19160), .Q(
        n8437) );
  NAND4X0 U27289 ( .IN1(n8403), .IN2(n8404), .IN3(n8405), .IN4(n8406), .QN(
        s11_data_o[0]) );
  OA22X1 U27290 ( .IN1(n1741), .IN2(n19112), .IN3(n1636), .IN4(n19095), .Q(
        n8403) );
  OA22X1 U27291 ( .IN1(n1913), .IN2(n19145), .IN3(n1827), .IN4(n19128), .Q(
        n8404) );
  OA22X1 U27292 ( .IN1(n2085), .IN2(n19178), .IN3(n1999), .IN4(n19162), .Q(
        n8405) );
  NAND4X0 U27293 ( .IN1(n8359), .IN2(n8360), .IN3(n8361), .IN4(n8362), .QN(
        s11_data_o[1]) );
  OA22X1 U27294 ( .IN1(n1740), .IN2(n19114), .IN3(n1635), .IN4(n19093), .Q(
        n8359) );
  OA22X1 U27295 ( .IN1(n1912), .IN2(n19147), .IN3(n1826), .IN4(n19126), .Q(
        n8360) );
  OA22X1 U27296 ( .IN1(n2084), .IN2(n19180), .IN3(n1998), .IN4(n19163), .Q(
        n8361) );
  NAND4X0 U27297 ( .IN1(n8315), .IN2(n8316), .IN3(n8317), .IN4(n8318), .QN(
        s11_data_o[2]) );
  OA22X1 U27298 ( .IN1(n1739), .IN2(n19115), .IN3(n1634), .IN4(n19086), .Q(
        n8315) );
  OA22X1 U27299 ( .IN1(n1911), .IN2(n19148), .IN3(n1825), .IN4(n19119), .Q(
        n8316) );
  OA22X1 U27300 ( .IN1(n2083), .IN2(n19181), .IN3(n1997), .IN4(n19167), .Q(
        n8317) );
  NAND4X0 U27301 ( .IN1(n8303), .IN2(n8304), .IN3(n8305), .IN4(n8306), .QN(
        s11_data_o[3]) );
  OA22X1 U27302 ( .IN1(n1738), .IN2(n19113), .IN3(n1633), .IN4(n19088), .Q(
        n8303) );
  OA22X1 U27303 ( .IN1(n1910), .IN2(n19146), .IN3(n1824), .IN4(n19121), .Q(
        n8304) );
  OA22X1 U27304 ( .IN1(n2082), .IN2(n19179), .IN3(n1996), .IN4(n19167), .Q(
        n8305) );
  NAND4X0 U27305 ( .IN1(n8299), .IN2(n8300), .IN3(n8301), .IN4(n8302), .QN(
        s11_data_o[4]) );
  OA22X1 U27306 ( .IN1(n1737), .IN2(n19114), .IN3(n1632), .IN4(n19103), .Q(
        n8299) );
  OA22X1 U27307 ( .IN1(n1909), .IN2(n19147), .IN3(n1823), .IN4(n19136), .Q(
        n8300) );
  OA22X1 U27308 ( .IN1(n2081), .IN2(n19180), .IN3(n1995), .IN4(n19167), .Q(
        n8301) );
  NAND4X0 U27309 ( .IN1(n8295), .IN2(n8296), .IN3(n8297), .IN4(n8298), .QN(
        s11_data_o[5]) );
  OA22X1 U27310 ( .IN1(n1736), .IN2(n19115), .IN3(n1631), .IN4(n19101), .Q(
        n8295) );
  OA22X1 U27311 ( .IN1(n1908), .IN2(n19148), .IN3(n1822), .IN4(n19134), .Q(
        n8296) );
  OA22X1 U27312 ( .IN1(n2080), .IN2(n19181), .IN3(n1994), .IN4(n19167), .Q(
        n8297) );
  NAND4X0 U27313 ( .IN1(n8291), .IN2(n8292), .IN3(n8293), .IN4(n8294), .QN(
        s11_data_o[6]) );
  OA22X1 U27314 ( .IN1(n1735), .IN2(n19111), .IN3(n1630), .IN4(n19101), .Q(
        n8291) );
  OA22X1 U27315 ( .IN1(n1907), .IN2(n19144), .IN3(n1821), .IN4(n19134), .Q(
        n8292) );
  OA22X1 U27316 ( .IN1(n2079), .IN2(n19176), .IN3(n1993), .IN4(n19168), .Q(
        n8293) );
  NAND4X0 U27317 ( .IN1(n8287), .IN2(n8288), .IN3(n8289), .IN4(n8290), .QN(
        s11_data_o[7]) );
  OA22X1 U27318 ( .IN1(n1734), .IN2(n19109), .IN3(n1629), .IN4(n19101), .Q(
        n8287) );
  OA22X1 U27319 ( .IN1(n1906), .IN2(n19142), .IN3(n1820), .IN4(n19134), .Q(
        n8288) );
  OA22X1 U27320 ( .IN1(n2078), .IN2(n19182), .IN3(n1992), .IN4(n19168), .Q(
        n8289) );
  NAND4X0 U27321 ( .IN1(n8283), .IN2(n8284), .IN3(n8285), .IN4(n8286), .QN(
        s11_data_o[8]) );
  OA22X1 U27322 ( .IN1(n1733), .IN2(n19116), .IN3(n1628), .IN4(n19101), .Q(
        n8283) );
  OA22X1 U27323 ( .IN1(n1905), .IN2(n19149), .IN3(n1819), .IN4(n19134), .Q(
        n8284) );
  OA22X1 U27324 ( .IN1(n2077), .IN2(n19182), .IN3(n1991), .IN4(n19168), .Q(
        n8285) );
  NAND4X0 U27325 ( .IN1(n8279), .IN2(n8280), .IN3(n8281), .IN4(n8282), .QN(
        s11_data_o[9]) );
  OA22X1 U27326 ( .IN1(n1732), .IN2(n19109), .IN3(n1627), .IN4(n19102), .Q(
        n8279) );
  OA22X1 U27327 ( .IN1(n1904), .IN2(n19142), .IN3(n1818), .IN4(n19135), .Q(
        n8280) );
  OA22X1 U27328 ( .IN1(n2076), .IN2(n19177), .IN3(n1990), .IN4(n19167), .Q(
        n8281) );
  NAND4X0 U27329 ( .IN1(n8399), .IN2(n8400), .IN3(n8401), .IN4(n8402), .QN(
        s11_data_o[10]) );
  OA22X1 U27330 ( .IN1(n1731), .IN2(n19111), .IN3(n1626), .IN4(n19096), .Q(
        n8399) );
  OA22X1 U27331 ( .IN1(n1903), .IN2(n19144), .IN3(n1817), .IN4(n19129), .Q(
        n8400) );
  OA22X1 U27332 ( .IN1(n2075), .IN2(n19176), .IN3(n1989), .IN4(n19156), .Q(
        n8401) );
  NAND4X0 U27333 ( .IN1(n8395), .IN2(n8396), .IN3(n8397), .IN4(n8398), .QN(
        s11_data_o[11]) );
  OA22X1 U27334 ( .IN1(n1730), .IN2(n19116), .IN3(n1625), .IN4(n19096), .Q(
        n8395) );
  OA22X1 U27335 ( .IN1(n1902), .IN2(n19149), .IN3(n1816), .IN4(n19129), .Q(
        n8396) );
  OA22X1 U27336 ( .IN1(n2074), .IN2(n19177), .IN3(n1988), .IN4(n19162), .Q(
        n8397) );
  NAND4X0 U27337 ( .IN1(n8391), .IN2(n8392), .IN3(n8393), .IN4(n8394), .QN(
        s11_data_o[12]) );
  OA22X1 U27338 ( .IN1(n1729), .IN2(n19112), .IN3(n1624), .IN4(n19096), .Q(
        n8391) );
  OA22X1 U27339 ( .IN1(n1901), .IN2(n19145), .IN3(n1815), .IN4(n19129), .Q(
        n8392) );
  OA22X1 U27340 ( .IN1(n2073), .IN2(n19178), .IN3(n1987), .IN4(n19156), .Q(
        n8393) );
  NAND4X0 U27341 ( .IN1(n8387), .IN2(n8388), .IN3(n8389), .IN4(n8390), .QN(
        s11_data_o[13]) );
  OA22X1 U27342 ( .IN1(n1728), .IN2(n19113), .IN3(n1623), .IN4(n19090), .Q(
        n8387) );
  OA22X1 U27343 ( .IN1(n1900), .IN2(n19146), .IN3(n1814), .IN4(n19123), .Q(
        n8388) );
  OA22X1 U27344 ( .IN1(n2072), .IN2(n19179), .IN3(n1986), .IN4(n19163), .Q(
        n8389) );
  NAND4X0 U27345 ( .IN1(n8383), .IN2(n8384), .IN3(n8385), .IN4(n8386), .QN(
        s11_data_o[14]) );
  OA22X1 U27346 ( .IN1(n1727), .IN2(n19113), .IN3(n1622), .IN4(n19095), .Q(
        n8383) );
  OA22X1 U27347 ( .IN1(n1899), .IN2(n19146), .IN3(n1813), .IN4(n19128), .Q(
        n8384) );
  OA22X1 U27348 ( .IN1(n2071), .IN2(n19179), .IN3(n1985), .IN4(n19163), .Q(
        n8385) );
  NAND4X0 U27349 ( .IN1(n8379), .IN2(n8380), .IN3(n8381), .IN4(n8382), .QN(
        s11_data_o[15]) );
  OA22X1 U27350 ( .IN1(n1726), .IN2(n19113), .IN3(n1621), .IN4(n19096), .Q(
        n8379) );
  OA22X1 U27351 ( .IN1(n1898), .IN2(n19146), .IN3(n1812), .IN4(n19129), .Q(
        n8380) );
  OA22X1 U27352 ( .IN1(n2070), .IN2(n19179), .IN3(n1984), .IN4(n19163), .Q(
        n8381) );
  NAND4X0 U27353 ( .IN1(n8375), .IN2(n8376), .IN3(n8377), .IN4(n8378), .QN(
        s11_data_o[16]) );
  OA22X1 U27354 ( .IN1(n1725), .IN2(n19113), .IN3(n1620), .IN4(n19097), .Q(
        n8375) );
  OA22X1 U27355 ( .IN1(n1897), .IN2(n19146), .IN3(n1811), .IN4(n19130), .Q(
        n8376) );
  OA22X1 U27356 ( .IN1(n2069), .IN2(n19179), .IN3(n1983), .IN4(n19164), .Q(
        n8377) );
  NAND4X0 U27357 ( .IN1(n8371), .IN2(n8372), .IN3(n8373), .IN4(n8374), .QN(
        s11_data_o[17]) );
  OA22X1 U27358 ( .IN1(n1724), .IN2(n19114), .IN3(n1619), .IN4(n19097), .Q(
        n8371) );
  OA22X1 U27359 ( .IN1(n1896), .IN2(n19147), .IN3(n1810), .IN4(n19130), .Q(
        n8372) );
  OA22X1 U27360 ( .IN1(n2068), .IN2(n19180), .IN3(n1982), .IN4(n19164), .Q(
        n8373) );
  NAND4X0 U27361 ( .IN1(n8367), .IN2(n8368), .IN3(n8369), .IN4(n8370), .QN(
        s11_data_o[18]) );
  OA22X1 U27362 ( .IN1(n1723), .IN2(n19114), .IN3(n1618), .IN4(n19097), .Q(
        n8367) );
  OA22X1 U27363 ( .IN1(n1895), .IN2(n19147), .IN3(n1809), .IN4(n19130), .Q(
        n8368) );
  OA22X1 U27364 ( .IN1(n2067), .IN2(n19180), .IN3(n1981), .IN4(n19164), .Q(
        n8369) );
  NAND4X0 U27365 ( .IN1(n8363), .IN2(n8364), .IN3(n8365), .IN4(n8366), .QN(
        s11_data_o[19]) );
  OA22X1 U27366 ( .IN1(n1722), .IN2(n19114), .IN3(n1617), .IN4(n19097), .Q(
        n8363) );
  OA22X1 U27367 ( .IN1(n1894), .IN2(n19147), .IN3(n1808), .IN4(n19130), .Q(
        n8364) );
  OA22X1 U27368 ( .IN1(n2066), .IN2(n19180), .IN3(n1980), .IN4(n19164), .Q(
        n8365) );
  NAND4X0 U27369 ( .IN1(n8355), .IN2(n8356), .IN3(n8357), .IN4(n8358), .QN(
        s11_data_o[20]) );
  OA22X1 U27370 ( .IN1(n1721), .IN2(n19115), .IN3(n1616), .IN4(n19094), .Q(
        n8355) );
  OA22X1 U27371 ( .IN1(n1893), .IN2(n19148), .IN3(n1807), .IN4(n19127), .Q(
        n8356) );
  OA22X1 U27372 ( .IN1(n2065), .IN2(n19181), .IN3(n1979), .IN4(n19167), .Q(
        n8357) );
  NAND4X0 U27373 ( .IN1(n8351), .IN2(n8352), .IN3(n8353), .IN4(n8354), .QN(
        s11_data_o[21]) );
  OA22X1 U27374 ( .IN1(n1720), .IN2(n19115), .IN3(n1615), .IN4(n19098), .Q(
        n8351) );
  OA22X1 U27375 ( .IN1(n1892), .IN2(n19148), .IN3(n1806), .IN4(n19131), .Q(
        n8352) );
  OA22X1 U27376 ( .IN1(n2064), .IN2(n19181), .IN3(n1978), .IN4(n19165), .Q(
        n8353) );
  NAND4X0 U27377 ( .IN1(n8347), .IN2(n8348), .IN3(n8349), .IN4(n8350), .QN(
        s11_data_o[22]) );
  OA22X1 U27378 ( .IN1(n1719), .IN2(n19113), .IN3(n1614), .IN4(n19098), .Q(
        n8347) );
  OA22X1 U27379 ( .IN1(n1891), .IN2(n19146), .IN3(n1805), .IN4(n19131), .Q(
        n8348) );
  OA22X1 U27380 ( .IN1(n2063), .IN2(n19179), .IN3(n1977), .IN4(n19165), .Q(
        n8349) );
  NAND4X0 U27381 ( .IN1(n8343), .IN2(n8344), .IN3(n8345), .IN4(n8346), .QN(
        s11_data_o[23]) );
  OA22X1 U27382 ( .IN1(n1718), .IN2(n19114), .IN3(n1613), .IN4(n19098), .Q(
        n8343) );
  OA22X1 U27383 ( .IN1(n1890), .IN2(n19147), .IN3(n1804), .IN4(n19131), .Q(
        n8344) );
  OA22X1 U27384 ( .IN1(n2062), .IN2(n19180), .IN3(n1976), .IN4(n19165), .Q(
        n8345) );
  NAND4X0 U27385 ( .IN1(n8339), .IN2(n8340), .IN3(n8341), .IN4(n8342), .QN(
        s11_data_o[24]) );
  OA22X1 U27386 ( .IN1(n1717), .IN2(n19112), .IN3(n1612), .IN4(n19099), .Q(
        n8339) );
  OA22X1 U27387 ( .IN1(n1889), .IN2(n19145), .IN3(n1803), .IN4(n19132), .Q(
        n8340) );
  OA22X1 U27388 ( .IN1(n2061), .IN2(n19178), .IN3(n1975), .IN4(n19166), .Q(
        n8341) );
  NAND4X0 U27389 ( .IN1(n8335), .IN2(n8336), .IN3(n8337), .IN4(n8338), .QN(
        s11_data_o[25]) );
  OA22X1 U27390 ( .IN1(n1716), .IN2(n19112), .IN3(n1611), .IN4(n19099), .Q(
        n8335) );
  OA22X1 U27391 ( .IN1(n1888), .IN2(n19145), .IN3(n1802), .IN4(n19132), .Q(
        n8336) );
  OA22X1 U27392 ( .IN1(n2060), .IN2(n19178), .IN3(n1974), .IN4(n19166), .Q(
        n8337) );
  NAND4X0 U27393 ( .IN1(n8331), .IN2(n8332), .IN3(n8333), .IN4(n8334), .QN(
        s11_data_o[26]) );
  OA22X1 U27394 ( .IN1(n1715), .IN2(n19111), .IN3(n1610), .IN4(n19099), .Q(
        n8331) );
  OA22X1 U27395 ( .IN1(n1887), .IN2(n19144), .IN3(n1801), .IN4(n19132), .Q(
        n8332) );
  OA22X1 U27396 ( .IN1(n2059), .IN2(n19176), .IN3(n1973), .IN4(n19166), .Q(
        n8333) );
  NAND4X0 U27397 ( .IN1(n8327), .IN2(n8328), .IN3(n8329), .IN4(n8330), .QN(
        s11_data_o[27]) );
  OA22X1 U27398 ( .IN1(n1714), .IN2(n19114), .IN3(n1609), .IN4(n19100), .Q(
        n8327) );
  OA22X1 U27399 ( .IN1(n1886), .IN2(n19147), .IN3(n1800), .IN4(n19133), .Q(
        n8328) );
  OA22X1 U27400 ( .IN1(n2058), .IN2(n19180), .IN3(n1972), .IN4(n19165), .Q(
        n8329) );
  NAND4X0 U27401 ( .IN1(n8323), .IN2(n8324), .IN3(n8325), .IN4(n8326), .QN(
        s11_data_o[28]) );
  OA22X1 U27402 ( .IN1(n1713), .IN2(n19115), .IN3(n1608), .IN4(n19100), .Q(
        n8323) );
  OA22X1 U27403 ( .IN1(n1885), .IN2(n19148), .IN3(n1799), .IN4(n19133), .Q(
        n8324) );
  OA22X1 U27404 ( .IN1(n2057), .IN2(n19181), .IN3(n1971), .IN4(n19166), .Q(
        n8325) );
  NAND4X0 U27405 ( .IN1(n8319), .IN2(n8320), .IN3(n8321), .IN4(n8322), .QN(
        s11_data_o[29]) );
  OA22X1 U27406 ( .IN1(n1712), .IN2(n19115), .IN3(n1607), .IN4(n19100), .Q(
        n8319) );
  OA22X1 U27407 ( .IN1(n1884), .IN2(n19148), .IN3(n1798), .IN4(n19133), .Q(
        n8320) );
  OA22X1 U27408 ( .IN1(n2056), .IN2(n19181), .IN3(n1970), .IN4(n19165), .Q(
        n8321) );
  NAND4X0 U27409 ( .IN1(n8311), .IN2(n8312), .IN3(n8313), .IN4(n8314), .QN(
        s11_data_o[30]) );
  OA22X1 U27410 ( .IN1(n1711), .IN2(n19115), .IN3(n1606), .IN4(n19102), .Q(
        n8311) );
  OA22X1 U27411 ( .IN1(n1883), .IN2(n19148), .IN3(n1797), .IN4(n19135), .Q(
        n8312) );
  OA22X1 U27412 ( .IN1(n2055), .IN2(n19181), .IN3(n1969), .IN4(n19167), .Q(
        n8313) );
  NAND4X0 U27413 ( .IN1(n8307), .IN2(n8308), .IN3(n8309), .IN4(n8310), .QN(
        s11_data_o[31]) );
  OA22X1 U27414 ( .IN1(n1710), .IN2(n19113), .IN3(n1605), .IN4(n19087), .Q(
        n8307) );
  OA22X1 U27415 ( .IN1(n1882), .IN2(n19146), .IN3(n1796), .IN4(n19120), .Q(
        n8308) );
  OA22X1 U27416 ( .IN1(n2054), .IN2(n19179), .IN3(n1968), .IN4(n19167), .Q(
        n8309) );
  NAND4X0 U27417 ( .IN1(n8547), .IN2(n8548), .IN3(n8549), .IN4(n8550), .QN(
        s10_stb_o) );
  OA22X1 U27418 ( .IN1(n1795), .IN2(n8557), .IN3(n1709), .IN4(n8558), .Q(n8547) );
  OA22X1 U27419 ( .IN1(n1967), .IN2(n8555), .IN3(n1881), .IN4(n8556), .Q(n8548) );
  OA22X1 U27420 ( .IN1(n2139), .IN2(n8553), .IN3(n2053), .IN4(n8554), .Q(n8549) );
  NAND4X0 U27421 ( .IN1(n8535), .IN2(n8536), .IN3(n8537), .IN4(n8538), .QN(
        s10_we_o) );
  OA22X1 U27422 ( .IN1(n1794), .IN2(n18977), .IN3(n1708), .IN4(n18971), .Q(
        n8535) );
  OA22X1 U27423 ( .IN1(n1966), .IN2(n19010), .IN3(n1880), .IN4(n18987), .Q(
        n8536) );
  OA22X1 U27424 ( .IN1(n2138), .IN2(n19043), .IN3(n2052), .IN4(n19036), .Q(
        n8537) );
  NAND4X0 U27425 ( .IN1(n8571), .IN2(n8572), .IN3(n8573), .IN4(n8574), .QN(
        s10_sel_o[0]) );
  OA22X1 U27426 ( .IN1(n1793), .IN2(n8545), .IN3(n1707), .IN4(n18969), .Q(
        n8571) );
  OA22X1 U27427 ( .IN1(n1965), .IN2(n19017), .IN3(n1879), .IN4(n19004), .Q(
        n8572) );
  OA22X1 U27428 ( .IN1(n2137), .IN2(n8541), .IN3(n2051), .IN4(n19037), .Q(
        n8573) );
  NAND4X0 U27429 ( .IN1(n8567), .IN2(n8568), .IN3(n8569), .IN4(n8570), .QN(
        s10_sel_o[1]) );
  OA22X1 U27430 ( .IN1(n1792), .IN2(n8545), .IN3(n1706), .IN4(n18969), .Q(
        n8567) );
  OA22X1 U27431 ( .IN1(n1964), .IN2(n19017), .IN3(n1878), .IN4(n19004), .Q(
        n8568) );
  OA22X1 U27432 ( .IN1(n2136), .IN2(n8541), .IN3(n2050), .IN4(n19037), .Q(
        n8569) );
  NAND4X0 U27433 ( .IN1(n8563), .IN2(n8564), .IN3(n8565), .IN4(n8566), .QN(
        s10_sel_o[2]) );
  OA22X1 U27434 ( .IN1(n1791), .IN2(n8545), .IN3(n1705), .IN4(n18971), .Q(
        n8563) );
  OA22X1 U27435 ( .IN1(n1963), .IN2(n19017), .IN3(n1877), .IN4(n18988), .Q(
        n8564) );
  OA22X1 U27436 ( .IN1(n2135), .IN2(n8541), .IN3(n2049), .IN4(n19021), .Q(
        n8565) );
  NAND4X0 U27437 ( .IN1(n8559), .IN2(n8560), .IN3(n8561), .IN4(n8562), .QN(
        s10_sel_o[3]) );
  OA22X1 U27438 ( .IN1(n1790), .IN2(n8545), .IN3(n1704), .IN4(n18971), .Q(
        n8559) );
  OA22X1 U27439 ( .IN1(n1962), .IN2(n19017), .IN3(n1876), .IN4(n18989), .Q(
        n8560) );
  OA22X1 U27440 ( .IN1(n2134), .IN2(n8541), .IN3(n2048), .IN4(n19019), .Q(
        n8561) );
  NAND4X0 U27441 ( .IN1(n8827), .IN2(n8828), .IN3(n8829), .IN4(n8830), .QN(
        s10_addr_o[0]) );
  OA22X1 U27442 ( .IN1(n1789), .IN2(n18977), .IN3(n1703), .IN4(n18954), .Q(
        n8827) );
  OA22X1 U27443 ( .IN1(n1961), .IN2(n19010), .IN3(n1875), .IN4(n18987), .Q(
        n8828) );
  OA22X1 U27444 ( .IN1(n2133), .IN2(n19043), .IN3(n2047), .IN4(n19033), .Q(
        n8829) );
  NAND4X0 U27445 ( .IN1(n8783), .IN2(n8784), .IN3(n8785), .IN4(n8786), .QN(
        s10_addr_o[1]) );
  OA22X1 U27446 ( .IN1(n1788), .IN2(n18979), .IN3(n1702), .IN4(n18957), .Q(
        n8783) );
  OA22X1 U27447 ( .IN1(n1960), .IN2(n19012), .IN3(n1874), .IN4(n18990), .Q(
        n8784) );
  OA22X1 U27448 ( .IN1(n2132), .IN2(n19045), .IN3(n2046), .IN4(n19021), .Q(
        n8785) );
  NAND4X0 U27449 ( .IN1(n8739), .IN2(n8740), .IN3(n8741), .IN4(n8742), .QN(
        s10_addr_o[2]) );
  OA22X1 U27450 ( .IN1(n1787), .IN2(n18981), .IN3(n1701), .IN4(n18961), .Q(
        n8739) );
  OA22X1 U27451 ( .IN1(n1959), .IN2(n19014), .IN3(n1873), .IN4(n18994), .Q(
        n8740) );
  OA22X1 U27452 ( .IN1(n2131), .IN2(n19047), .IN3(n2045), .IN4(n19025), .Q(
        n8741) );
  NAND4X0 U27453 ( .IN1(n8727), .IN2(n8728), .IN3(n8729), .IN4(n8730), .QN(
        s10_addr_o[3]) );
  OA22X1 U27454 ( .IN1(n1786), .IN2(n8545), .IN3(n1699), .IN4(n18962), .Q(
        n8727) );
  OA22X1 U27455 ( .IN1(n1958), .IN2(n19017), .IN3(n1872), .IN4(n18995), .Q(
        n8728) );
  OA22X1 U27456 ( .IN1(n2130), .IN2(n8541), .IN3(n2044), .IN4(n19026), .Q(
        n8729) );
  NAND4X0 U27457 ( .IN1(n8723), .IN2(n8724), .IN3(n8725), .IN4(n8726), .QN(
        s10_addr_o[4]) );
  OA22X1 U27458 ( .IN1(n1785), .IN2(n18980), .IN3(n1697), .IN4(n18962), .Q(
        n8723) );
  OA22X1 U27459 ( .IN1(n1957), .IN2(n19013), .IN3(n1871), .IN4(n18995), .Q(
        n8724) );
  OA22X1 U27460 ( .IN1(n2129), .IN2(n19046), .IN3(n2043), .IN4(n19026), .Q(
        n8725) );
  NAND4X0 U27461 ( .IN1(n8719), .IN2(n8720), .IN3(n8721), .IN4(n8722), .QN(
        s10_addr_o[5]) );
  OA22X1 U27462 ( .IN1(n1784), .IN2(n8545), .IN3(n1696), .IN4(n18963), .Q(
        n8719) );
  OA22X1 U27463 ( .IN1(n1956), .IN2(n19017), .IN3(n1870), .IN4(n18996), .Q(
        n8720) );
  OA22X1 U27464 ( .IN1(n2128), .IN2(n8541), .IN3(n2042), .IN4(n19027), .Q(
        n8721) );
  NAND4X0 U27465 ( .IN1(n8715), .IN2(n8716), .IN3(n8717), .IN4(n8718), .QN(
        s10_addr_o[6]) );
  OA22X1 U27466 ( .IN1(n1783), .IN2(n18982), .IN3(n1679), .IN4(n18963), .Q(
        n8715) );
  OA22X1 U27467 ( .IN1(n1955), .IN2(n19015), .IN3(n1869), .IN4(n18996), .Q(
        n8716) );
  OA22X1 U27468 ( .IN1(n2127), .IN2(n19048), .IN3(n2041), .IN4(n19027), .Q(
        n8717) );
  NAND4X0 U27469 ( .IN1(n8711), .IN2(n8712), .IN3(n8713), .IN4(n8714), .QN(
        s10_addr_o[7]) );
  OA22X1 U27470 ( .IN1(n1782), .IN2(n18982), .IN3(n1678), .IN4(n18963), .Q(
        n8711) );
  OA22X1 U27471 ( .IN1(n1954), .IN2(n19015), .IN3(n1868), .IN4(n18996), .Q(
        n8712) );
  OA22X1 U27472 ( .IN1(n2126), .IN2(n19048), .IN3(n2040), .IN4(n19027), .Q(
        n8713) );
  NAND4X0 U27473 ( .IN1(n8707), .IN2(n8708), .IN3(n8709), .IN4(n8710), .QN(
        s10_addr_o[8]) );
  OA22X1 U27474 ( .IN1(n1781), .IN2(n18982), .IN3(n1677), .IN4(n18964), .Q(
        n8707) );
  OA22X1 U27475 ( .IN1(n1953), .IN2(n19015), .IN3(n1867), .IN4(n18997), .Q(
        n8708) );
  OA22X1 U27476 ( .IN1(n2125), .IN2(n19048), .IN3(n2039), .IN4(n19028), .Q(
        n8709) );
  NAND4X0 U27477 ( .IN1(n8703), .IN2(n8704), .IN3(n8705), .IN4(n8706), .QN(
        s10_addr_o[9]) );
  OA22X1 U27478 ( .IN1(n1780), .IN2(n18982), .IN3(n1676), .IN4(n18964), .Q(
        n8703) );
  OA22X1 U27479 ( .IN1(n1952), .IN2(n19015), .IN3(n1866), .IN4(n18997), .Q(
        n8704) );
  OA22X1 U27480 ( .IN1(n2124), .IN2(n19048), .IN3(n2038), .IN4(n19028), .Q(
        n8705) );
  NAND4X0 U27481 ( .IN1(n8823), .IN2(n8824), .IN3(n8825), .IN4(n8826), .QN(
        s10_addr_o[10]) );
  OA22X1 U27482 ( .IN1(n1779), .IN2(n18977), .IN3(n1675), .IN4(n18954), .Q(
        n8823) );
  OA22X1 U27483 ( .IN1(n1951), .IN2(n19010), .IN3(n1865), .IN4(n18987), .Q(
        n8824) );
  OA22X1 U27484 ( .IN1(n2123), .IN2(n19043), .IN3(n2037), .IN4(n19036), .Q(
        n8825) );
  NAND4X0 U27485 ( .IN1(n8819), .IN2(n8820), .IN3(n8821), .IN4(n8822), .QN(
        s10_addr_o[11]) );
  OA22X1 U27486 ( .IN1(n1778), .IN2(n18977), .IN3(n1674), .IN4(n18954), .Q(
        n8819) );
  OA22X1 U27487 ( .IN1(n1950), .IN2(n19010), .IN3(n1864), .IN4(n18987), .Q(
        n8820) );
  OA22X1 U27488 ( .IN1(n2122), .IN2(n19043), .IN3(n2036), .IN4(n19031), .Q(
        n8821) );
  NAND4X0 U27489 ( .IN1(n8815), .IN2(n8816), .IN3(n8817), .IN4(n8818), .QN(
        s10_addr_o[12]) );
  OA22X1 U27490 ( .IN1(n1777), .IN2(n18977), .IN3(n1673), .IN4(n18955), .Q(
        n8815) );
  OA22X1 U27491 ( .IN1(n1949), .IN2(n19010), .IN3(n1863), .IN4(n18988), .Q(
        n8816) );
  OA22X1 U27492 ( .IN1(n2121), .IN2(n19043), .IN3(n2035), .IN4(n19020), .Q(
        n8817) );
  NAND4X0 U27493 ( .IN1(n8811), .IN2(n8812), .IN3(n8813), .IN4(n8814), .QN(
        s10_addr_o[13]) );
  OA22X1 U27494 ( .IN1(n1776), .IN2(n18978), .IN3(n1672), .IN4(n18955), .Q(
        n8811) );
  OA22X1 U27495 ( .IN1(n1948), .IN2(n19011), .IN3(n1862), .IN4(n18988), .Q(
        n8812) );
  OA22X1 U27496 ( .IN1(n2120), .IN2(n19044), .IN3(n2034), .IN4(n19020), .Q(
        n8813) );
  NAND4X0 U27497 ( .IN1(n8807), .IN2(n8808), .IN3(n8809), .IN4(n8810), .QN(
        s10_addr_o[14]) );
  OA22X1 U27498 ( .IN1(n1775), .IN2(n18978), .IN3(n1671), .IN4(n18955), .Q(
        n8807) );
  OA22X1 U27499 ( .IN1(n1947), .IN2(n19011), .IN3(n1861), .IN4(n18988), .Q(
        n8808) );
  OA22X1 U27500 ( .IN1(n2119), .IN2(n19044), .IN3(n2033), .IN4(n19020), .Q(
        n8809) );
  NAND4X0 U27501 ( .IN1(n8803), .IN2(n8804), .IN3(n8805), .IN4(n8806), .QN(
        s10_addr_o[15]) );
  OA22X1 U27502 ( .IN1(n1774), .IN2(n18978), .IN3(n1670), .IN4(n18956), .Q(
        n8803) );
  OA22X1 U27503 ( .IN1(n1946), .IN2(n19011), .IN3(n1860), .IN4(n18989), .Q(
        n8804) );
  OA22X1 U27504 ( .IN1(n2118), .IN2(n19044), .IN3(n2032), .IN4(n19031), .Q(
        n8805) );
  NAND4X0 U27505 ( .IN1(n8799), .IN2(n8800), .IN3(n8801), .IN4(n8802), .QN(
        s10_addr_o[16]) );
  OA22X1 U27506 ( .IN1(n1773), .IN2(n18978), .IN3(n1669), .IN4(n18956), .Q(
        n8799) );
  OA22X1 U27507 ( .IN1(n1945), .IN2(n19011), .IN3(n1859), .IN4(n18989), .Q(
        n8800) );
  OA22X1 U27508 ( .IN1(n2117), .IN2(n19044), .IN3(n2031), .IN4(n19020), .Q(
        n8801) );
  NAND4X0 U27509 ( .IN1(n8795), .IN2(n8796), .IN3(n8797), .IN4(n8798), .QN(
        s10_addr_o[17]) );
  OA22X1 U27510 ( .IN1(n1772), .IN2(n18979), .IN3(n1668), .IN4(n18956), .Q(
        n8795) );
  OA22X1 U27511 ( .IN1(n1944), .IN2(n19012), .IN3(n1858), .IN4(n18989), .Q(
        n8796) );
  OA22X1 U27512 ( .IN1(n2116), .IN2(n19045), .IN3(n2030), .IN4(n19032), .Q(
        n8797) );
  NAND4X0 U27513 ( .IN1(n8791), .IN2(n8792), .IN3(n8793), .IN4(n8794), .QN(
        s10_addr_o[18]) );
  OA22X1 U27514 ( .IN1(n1771), .IN2(n18979), .IN3(n1667), .IN4(n18957), .Q(
        n8791) );
  OA22X1 U27515 ( .IN1(n1943), .IN2(n19012), .IN3(n1857), .IN4(n18990), .Q(
        n8792) );
  OA22X1 U27516 ( .IN1(n2115), .IN2(n19045), .IN3(n2029), .IN4(n19021), .Q(
        n8793) );
  NAND4X0 U27517 ( .IN1(n8787), .IN2(n8788), .IN3(n8789), .IN4(n8790), .QN(
        s10_addr_o[19]) );
  OA22X1 U27518 ( .IN1(n1770), .IN2(n18979), .IN3(n1666), .IN4(n18957), .Q(
        n8787) );
  OA22X1 U27519 ( .IN1(n1942), .IN2(n19012), .IN3(n1856), .IN4(n18990), .Q(
        n8788) );
  OA22X1 U27520 ( .IN1(n2114), .IN2(n19045), .IN3(n2028), .IN4(n19021), .Q(
        n8789) );
  NAND4X0 U27521 ( .IN1(n8779), .IN2(n8780), .IN3(n8781), .IN4(n8782), .QN(
        s10_addr_o[20]) );
  OA22X1 U27522 ( .IN1(n1769), .IN2(n18978), .IN3(n1665), .IN4(n18958), .Q(
        n8779) );
  OA22X1 U27523 ( .IN1(n1941), .IN2(n19011), .IN3(n1855), .IN4(n18991), .Q(
        n8780) );
  OA22X1 U27524 ( .IN1(n2113), .IN2(n19044), .IN3(n2027), .IN4(n19022), .Q(
        n8781) );
  NAND4X0 U27525 ( .IN1(n8775), .IN2(n8776), .IN3(n8777), .IN4(n8778), .QN(
        s10_addr_o[21]) );
  OA22X1 U27526 ( .IN1(n1768), .IN2(n18978), .IN3(n1664), .IN4(n18958), .Q(
        n8775) );
  OA22X1 U27527 ( .IN1(n1940), .IN2(n19011), .IN3(n1854), .IN4(n18991), .Q(
        n8776) );
  OA22X1 U27528 ( .IN1(n2112), .IN2(n19044), .IN3(n2026), .IN4(n19022), .Q(
        n8777) );
  NAND4X0 U27529 ( .IN1(n8771), .IN2(n8772), .IN3(n8773), .IN4(n8774), .QN(
        s10_addr_o[22]) );
  OA22X1 U27530 ( .IN1(n1767), .IN2(n18977), .IN3(n1663), .IN4(n18958), .Q(
        n8771) );
  OA22X1 U27531 ( .IN1(n1939), .IN2(n19010), .IN3(n1853), .IN4(n18991), .Q(
        n8772) );
  OA22X1 U27532 ( .IN1(n2111), .IN2(n19043), .IN3(n2025), .IN4(n19022), .Q(
        n8773) );
  NAND4X0 U27533 ( .IN1(n8767), .IN2(n8768), .IN3(n8769), .IN4(n8770), .QN(
        s10_addr_o[23]) );
  OA22X1 U27534 ( .IN1(n1766), .IN2(n18978), .IN3(n1662), .IN4(n18959), .Q(
        n8767) );
  OA22X1 U27535 ( .IN1(n1938), .IN2(n19011), .IN3(n1852), .IN4(n18992), .Q(
        n8768) );
  OA22X1 U27536 ( .IN1(n2110), .IN2(n19044), .IN3(n2024), .IN4(n19023), .Q(
        n8769) );
  NAND4X0 U27537 ( .IN1(n8763), .IN2(n8764), .IN3(n8765), .IN4(n8766), .QN(
        s10_addr_o[24]) );
  OA22X1 U27538 ( .IN1(n1765), .IN2(n18980), .IN3(n1661), .IN4(n18959), .Q(
        n8763) );
  OA22X1 U27539 ( .IN1(n1937), .IN2(n19013), .IN3(n1851), .IN4(n18992), .Q(
        n8764) );
  OA22X1 U27540 ( .IN1(n2109), .IN2(n19046), .IN3(n2023), .IN4(n19023), .Q(
        n8765) );
  NAND4X0 U27541 ( .IN1(n8759), .IN2(n8760), .IN3(n8761), .IN4(n8762), .QN(
        s10_addr_o[25]) );
  OA22X1 U27542 ( .IN1(n1764), .IN2(n18980), .IN3(n1660), .IN4(n18959), .Q(
        n8759) );
  OA22X1 U27543 ( .IN1(n1936), .IN2(n19013), .IN3(n1850), .IN4(n18992), .Q(
        n8760) );
  OA22X1 U27544 ( .IN1(n2108), .IN2(n19046), .IN3(n2022), .IN4(n19023), .Q(
        n8761) );
  NAND4X0 U27545 ( .IN1(n8755), .IN2(n8756), .IN3(n8757), .IN4(n8758), .QN(
        s10_addr_o[26]) );
  OA22X1 U27546 ( .IN1(n1763), .IN2(n18980), .IN3(n1659), .IN4(n18960), .Q(
        n8755) );
  OA22X1 U27547 ( .IN1(n1935), .IN2(n19013), .IN3(n1849), .IN4(n18993), .Q(
        n8756) );
  OA22X1 U27548 ( .IN1(n2107), .IN2(n19046), .IN3(n2021), .IN4(n19024), .Q(
        n8757) );
  NAND4X0 U27549 ( .IN1(n8751), .IN2(n8752), .IN3(n8753), .IN4(n8754), .QN(
        s10_addr_o[27]) );
  OA22X1 U27550 ( .IN1(n1762), .IN2(n18980), .IN3(n1658), .IN4(n18960), .Q(
        n8751) );
  OA22X1 U27551 ( .IN1(n1934), .IN2(n19013), .IN3(n1848), .IN4(n18993), .Q(
        n8752) );
  OA22X1 U27552 ( .IN1(n2106), .IN2(n19046), .IN3(n2020), .IN4(n19024), .Q(
        n8753) );
  NAND4X0 U27553 ( .IN1(n8747), .IN2(n8748), .IN3(n8749), .IN4(n8750), .QN(
        s10_addr_o[28]) );
  OA22X1 U27554 ( .IN1(n1761), .IN2(n18981), .IN3(n1657), .IN4(n18960), .Q(
        n8747) );
  OA22X1 U27555 ( .IN1(n1933), .IN2(n19014), .IN3(n1847), .IN4(n18993), .Q(
        n8748) );
  OA22X1 U27556 ( .IN1(n2105), .IN2(n19047), .IN3(n2019), .IN4(n19024), .Q(
        n8749) );
  NAND4X0 U27557 ( .IN1(n8743), .IN2(n8744), .IN3(n8745), .IN4(n8746), .QN(
        s10_addr_o[29]) );
  OA22X1 U27558 ( .IN1(n1760), .IN2(n18981), .IN3(n1656), .IN4(n18961), .Q(
        n8743) );
  OA22X1 U27559 ( .IN1(n1932), .IN2(n19014), .IN3(n1846), .IN4(n18994), .Q(
        n8744) );
  OA22X1 U27560 ( .IN1(n2104), .IN2(n19047), .IN3(n2018), .IN4(n19025), .Q(
        n8745) );
  NAND4X0 U27561 ( .IN1(n8735), .IN2(n8736), .IN3(n8737), .IN4(n8738), .QN(
        s10_addr_o[30]) );
  OA22X1 U27562 ( .IN1(n1759), .IN2(n18981), .IN3(n1655), .IN4(n18961), .Q(
        n8735) );
  OA22X1 U27563 ( .IN1(n1931), .IN2(n19014), .IN3(n1845), .IN4(n18994), .Q(
        n8736) );
  OA22X1 U27564 ( .IN1(n2103), .IN2(n19047), .IN3(n2017), .IN4(n19025), .Q(
        n8737) );
  NAND4X0 U27565 ( .IN1(n8731), .IN2(n8732), .IN3(n8733), .IN4(n8734), .QN(
        s10_addr_o[31]) );
  OA22X1 U27566 ( .IN1(n1758), .IN2(n18981), .IN3(n1650), .IN4(n18962), .Q(
        n8731) );
  OA22X1 U27567 ( .IN1(n1930), .IN2(n19014), .IN3(n1844), .IN4(n18995), .Q(
        n8732) );
  OA22X1 U27568 ( .IN1(n2102), .IN2(n19047), .IN3(n2016), .IN4(n19026), .Q(
        n8733) );
  NAND4X0 U27569 ( .IN1(n8699), .IN2(n8700), .IN3(n8701), .IN4(n8702), .QN(
        s10_data_o[0]) );
  OA22X1 U27570 ( .IN1(n1741), .IN2(n18983), .IN3(n1636), .IN4(n18964), .Q(
        n8699) );
  OA22X1 U27571 ( .IN1(n1913), .IN2(n19012), .IN3(n1827), .IN4(n18997), .Q(
        n8700) );
  OA22X1 U27572 ( .IN1(n2085), .IN2(n19049), .IN3(n1999), .IN4(n19028), .Q(
        n8701) );
  NAND4X0 U27573 ( .IN1(n8655), .IN2(n8656), .IN3(n8657), .IN4(n8658), .QN(
        s10_data_o[1]) );
  OA22X1 U27574 ( .IN1(n1740), .IN2(n18984), .IN3(n1635), .IN4(n18966), .Q(
        n8655) );
  OA22X1 U27575 ( .IN1(n1912), .IN2(n19016), .IN3(n1826), .IN4(n19001), .Q(
        n8656) );
  OA22X1 U27576 ( .IN1(n2084), .IN2(n19045), .IN3(n1998), .IN4(n19029), .Q(
        n8657) );
  NAND4X0 U27577 ( .IN1(n8611), .IN2(n8612), .IN3(n8613), .IN4(n8614), .QN(
        s10_data_o[2]) );
  OA22X1 U27578 ( .IN1(n1739), .IN2(n18979), .IN3(n1634), .IN4(n18969), .Q(
        n8611) );
  OA22X1 U27579 ( .IN1(n1911), .IN2(n8543), .IN3(n1825), .IN4(n19004), .Q(
        n8612) );
  OA22X1 U27580 ( .IN1(n2083), .IN2(n19050), .IN3(n1997), .IN4(n19034), .Q(
        n8613) );
  NAND4X0 U27581 ( .IN1(n8599), .IN2(n8600), .IN3(n8601), .IN4(n8602), .QN(
        s10_data_o[3]) );
  OA22X1 U27582 ( .IN1(n1738), .IN2(n18982), .IN3(n1633), .IN4(n18969), .Q(
        n8599) );
  OA22X1 U27583 ( .IN1(n1910), .IN2(n8543), .IN3(n1824), .IN4(n19004), .Q(
        n8600) );
  OA22X1 U27584 ( .IN1(n2082), .IN2(n19050), .IN3(n1996), .IN4(n19035), .Q(
        n8601) );
  NAND4X0 U27585 ( .IN1(n8595), .IN2(n8596), .IN3(n8597), .IN4(n8598), .QN(
        s10_data_o[4]) );
  OA22X1 U27586 ( .IN1(n1737), .IN2(n18980), .IN3(n1632), .IN4(n18969), .Q(
        n8595) );
  OA22X1 U27587 ( .IN1(n1909), .IN2(n19013), .IN3(n1823), .IN4(n19004), .Q(
        n8596) );
  OA22X1 U27588 ( .IN1(n2081), .IN2(n19046), .IN3(n1995), .IN4(n19035), .Q(
        n8597) );
  NAND4X0 U27589 ( .IN1(n8591), .IN2(n8592), .IN3(n8593), .IN4(n8594), .QN(
        s10_data_o[5]) );
  OA22X1 U27590 ( .IN1(n1736), .IN2(n18984), .IN3(n1631), .IN4(n18969), .Q(
        n8591) );
  OA22X1 U27591 ( .IN1(n1908), .IN2(n8543), .IN3(n1822), .IN4(n19004), .Q(
        n8592) );
  OA22X1 U27592 ( .IN1(n2080), .IN2(n19048), .IN3(n1994), .IN4(n19035), .Q(
        n8593) );
  NAND4X0 U27593 ( .IN1(n8587), .IN2(n8588), .IN3(n8589), .IN4(n8590), .QN(
        s10_data_o[6]) );
  OA22X1 U27594 ( .IN1(n1735), .IN2(n18984), .IN3(n1630), .IN4(n18970), .Q(
        n8587) );
  OA22X1 U27595 ( .IN1(n1907), .IN2(n19016), .IN3(n1821), .IN4(n19002), .Q(
        n8588) );
  OA22X1 U27596 ( .IN1(n2079), .IN2(n19050), .IN3(n1993), .IN4(n19036), .Q(
        n8589) );
  NAND4X0 U27597 ( .IN1(n8583), .IN2(n8584), .IN3(n8585), .IN4(n8586), .QN(
        s10_data_o[7]) );
  OA22X1 U27598 ( .IN1(n1734), .IN2(n18984), .IN3(n1629), .IN4(n18970), .Q(
        n8583) );
  OA22X1 U27599 ( .IN1(n1906), .IN2(n19016), .IN3(n1820), .IN4(n19002), .Q(
        n8584) );
  OA22X1 U27600 ( .IN1(n2078), .IN2(n19050), .IN3(n1992), .IN4(n19036), .Q(
        n8585) );
  NAND4X0 U27601 ( .IN1(n8579), .IN2(n8580), .IN3(n8581), .IN4(n8582), .QN(
        s10_data_o[8]) );
  OA22X1 U27602 ( .IN1(n1733), .IN2(n18984), .IN3(n1628), .IN4(n18970), .Q(
        n8579) );
  OA22X1 U27603 ( .IN1(n1905), .IN2(n19016), .IN3(n1819), .IN4(n19002), .Q(
        n8580) );
  OA22X1 U27604 ( .IN1(n2077), .IN2(n19050), .IN3(n1991), .IN4(n19036), .Q(
        n8581) );
  NAND4X0 U27605 ( .IN1(n8575), .IN2(n8576), .IN3(n8577), .IN4(n8578), .QN(
        s10_data_o[9]) );
  OA22X1 U27606 ( .IN1(n1732), .IN2(n18984), .IN3(n1627), .IN4(n18969), .Q(
        n8575) );
  OA22X1 U27607 ( .IN1(n1904), .IN2(n19016), .IN3(n1818), .IN4(n19002), .Q(
        n8576) );
  OA22X1 U27608 ( .IN1(n2076), .IN2(n19050), .IN3(n1990), .IN4(n19037), .Q(
        n8577) );
  NAND4X0 U27609 ( .IN1(n8695), .IN2(n8696), .IN3(n8697), .IN4(n8698), .QN(
        s10_data_o[10]) );
  OA22X1 U27610 ( .IN1(n1731), .IN2(n18983), .IN3(n1626), .IN4(n18965), .Q(
        n8695) );
  OA22X1 U27611 ( .IN1(n1903), .IN2(n19010), .IN3(n1817), .IN4(n18998), .Q(
        n8696) );
  OA22X1 U27612 ( .IN1(n2075), .IN2(n19049), .IN3(n1989), .IN4(n19022), .Q(
        n8697) );
  NAND4X0 U27613 ( .IN1(n8691), .IN2(n8692), .IN3(n8693), .IN4(n8694), .QN(
        s10_data_o[11]) );
  OA22X1 U27614 ( .IN1(n1730), .IN2(n18983), .IN3(n1625), .IN4(n18965), .Q(
        n8691) );
  OA22X1 U27615 ( .IN1(n1902), .IN2(n19017), .IN3(n1816), .IN4(n18998), .Q(
        n8692) );
  OA22X1 U27616 ( .IN1(n2074), .IN2(n19049), .IN3(n1988), .IN4(n19028), .Q(
        n8693) );
  NAND4X0 U27617 ( .IN1(n8687), .IN2(n8688), .IN3(n8689), .IN4(n8690), .QN(
        s10_data_o[12]) );
  OA22X1 U27618 ( .IN1(n1729), .IN2(n18983), .IN3(n1624), .IN4(n18965), .Q(
        n8687) );
  OA22X1 U27619 ( .IN1(n1901), .IN2(n19013), .IN3(n1815), .IN4(n18998), .Q(
        n8688) );
  OA22X1 U27620 ( .IN1(n2073), .IN2(n19049), .IN3(n1987), .IN4(n19022), .Q(
        n8689) );
  NAND4X0 U27621 ( .IN1(n8683), .IN2(n8684), .IN3(n8685), .IN4(n8686), .QN(
        s10_data_o[13]) );
  OA22X1 U27622 ( .IN1(n1728), .IN2(n18981), .IN3(n1623), .IN4(n18966), .Q(
        n8683) );
  OA22X1 U27623 ( .IN1(n1900), .IN2(n19014), .IN3(n1814), .IN4(n18999), .Q(
        n8684) );
  OA22X1 U27624 ( .IN1(n2072), .IN2(n19047), .IN3(n1986), .IN4(n19029), .Q(
        n8685) );
  NAND4X0 U27625 ( .IN1(n8679), .IN2(n8680), .IN3(n8681), .IN4(n8682), .QN(
        s10_data_o[14]) );
  OA22X1 U27626 ( .IN1(n1727), .IN2(n18980), .IN3(n1622), .IN4(n18966), .Q(
        n8679) );
  OA22X1 U27627 ( .IN1(n1899), .IN2(n19013), .IN3(n1813), .IN4(n18999), .Q(
        n8680) );
  OA22X1 U27628 ( .IN1(n2071), .IN2(n19046), .IN3(n1985), .IN4(n19029), .Q(
        n8681) );
  NAND4X0 U27629 ( .IN1(n8675), .IN2(n8676), .IN3(n8677), .IN4(n8678), .QN(
        s10_data_o[15]) );
  OA22X1 U27630 ( .IN1(n1726), .IN2(n18981), .IN3(n1621), .IN4(n18966), .Q(
        n8675) );
  OA22X1 U27631 ( .IN1(n1898), .IN2(n19014), .IN3(n1812), .IN4(n18999), .Q(
        n8676) );
  OA22X1 U27632 ( .IN1(n2070), .IN2(n19047), .IN3(n1984), .IN4(n19029), .Q(
        n8677) );
  NAND4X0 U27633 ( .IN1(n8671), .IN2(n8672), .IN3(n8673), .IN4(n8674), .QN(
        s10_data_o[16]) );
  OA22X1 U27634 ( .IN1(n1725), .IN2(n18977), .IN3(n1620), .IN4(n18967), .Q(
        n8671) );
  OA22X1 U27635 ( .IN1(n1897), .IN2(n19010), .IN3(n1811), .IN4(n19000), .Q(
        n8672) );
  OA22X1 U27636 ( .IN1(n2069), .IN2(n19043), .IN3(n1983), .IN4(n19030), .Q(
        n8673) );
  NAND4X0 U27637 ( .IN1(n8667), .IN2(n8668), .IN3(n8669), .IN4(n8670), .QN(
        s10_data_o[17]) );
  OA22X1 U27638 ( .IN1(n1724), .IN2(n18982), .IN3(n1619), .IN4(n18967), .Q(
        n8667) );
  OA22X1 U27639 ( .IN1(n1896), .IN2(n19015), .IN3(n1810), .IN4(n19000), .Q(
        n8668) );
  OA22X1 U27640 ( .IN1(n2068), .IN2(n19049), .IN3(n1982), .IN4(n19030), .Q(
        n8669) );
  NAND4X0 U27641 ( .IN1(n8663), .IN2(n8664), .IN3(n8665), .IN4(n8666), .QN(
        s10_data_o[18]) );
  OA22X1 U27642 ( .IN1(n1723), .IN2(n18979), .IN3(n1618), .IN4(n18967), .Q(
        n8663) );
  OA22X1 U27643 ( .IN1(n1895), .IN2(n19012), .IN3(n1809), .IN4(n19000), .Q(
        n8664) );
  OA22X1 U27644 ( .IN1(n2067), .IN2(n19043), .IN3(n1981), .IN4(n19030), .Q(
        n8665) );
  NAND4X0 U27645 ( .IN1(n8659), .IN2(n8660), .IN3(n8661), .IN4(n8662), .QN(
        s10_data_o[19]) );
  OA22X1 U27646 ( .IN1(n1722), .IN2(n18983), .IN3(n1617), .IN4(n18967), .Q(
        n8659) );
  OA22X1 U27647 ( .IN1(n1894), .IN2(n19016), .IN3(n1808), .IN4(n19001), .Q(
        n8660) );
  OA22X1 U27648 ( .IN1(n2066), .IN2(n19046), .IN3(n1980), .IN4(n19030), .Q(
        n8661) );
  NAND4X0 U27649 ( .IN1(n8651), .IN2(n8652), .IN3(n8653), .IN4(n8654), .QN(
        s10_data_o[20]) );
  OA22X1 U27650 ( .IN1(n1721), .IN2(n18984), .IN3(n1616), .IN4(n18966), .Q(
        n8651) );
  OA22X1 U27651 ( .IN1(n1893), .IN2(n19016), .IN3(n1807), .IN4(n19001), .Q(
        n8652) );
  OA22X1 U27652 ( .IN1(n2065), .IN2(n19050), .IN3(n1979), .IN4(n19029), .Q(
        n8653) );
  NAND4X0 U27653 ( .IN1(n8647), .IN2(n8648), .IN3(n8649), .IN4(n8650), .QN(
        s10_data_o[21]) );
  OA22X1 U27654 ( .IN1(n1720), .IN2(n18982), .IN3(n1615), .IN4(n18969), .Q(
        n8647) );
  OA22X1 U27655 ( .IN1(n1892), .IN2(n19015), .IN3(n1806), .IN4(n19002), .Q(
        n8648) );
  OA22X1 U27656 ( .IN1(n2064), .IN2(n19048), .IN3(n1978), .IN4(n19031), .Q(
        n8649) );
  NAND4X0 U27657 ( .IN1(n8643), .IN2(n8644), .IN3(n8645), .IN4(n8646), .QN(
        s10_data_o[22]) );
  OA22X1 U27658 ( .IN1(n1719), .IN2(n18979), .IN3(n1614), .IN4(n18953), .Q(
        n8643) );
  OA22X1 U27659 ( .IN1(n1891), .IN2(n19012), .IN3(n1805), .IN4(n19002), .Q(
        n8644) );
  OA22X1 U27660 ( .IN1(n2063), .IN2(n19045), .IN3(n1977), .IN4(n19031), .Q(
        n8645) );
  NAND4X0 U27661 ( .IN1(n8639), .IN2(n8640), .IN3(n8641), .IN4(n8642), .QN(
        s10_data_o[23]) );
  OA22X1 U27662 ( .IN1(n1718), .IN2(n18983), .IN3(n1613), .IN4(n18971), .Q(
        n8639) );
  OA22X1 U27663 ( .IN1(n1890), .IN2(n19011), .IN3(n1804), .IN4(n19002), .Q(
        n8640) );
  OA22X1 U27664 ( .IN1(n2062), .IN2(n19049), .IN3(n1976), .IN4(n19031), .Q(
        n8641) );
  NAND4X0 U27665 ( .IN1(n8635), .IN2(n8636), .IN3(n8637), .IN4(n8638), .QN(
        s10_data_o[24]) );
  OA22X1 U27666 ( .IN1(n1717), .IN2(n18984), .IN3(n1612), .IN4(n18968), .Q(
        n8635) );
  OA22X1 U27667 ( .IN1(n1889), .IN2(n19016), .IN3(n1803), .IN4(n19003), .Q(
        n8636) );
  OA22X1 U27668 ( .IN1(n2061), .IN2(n19050), .IN3(n1975), .IN4(n19032), .Q(
        n8637) );
  NAND4X0 U27669 ( .IN1(n8631), .IN2(n8632), .IN3(n8633), .IN4(n8634), .QN(
        s10_data_o[25]) );
  OA22X1 U27670 ( .IN1(n1716), .IN2(n18982), .IN3(n1611), .IN4(n18968), .Q(
        n8631) );
  OA22X1 U27671 ( .IN1(n1888), .IN2(n19015), .IN3(n1802), .IN4(n19003), .Q(
        n8632) );
  OA22X1 U27672 ( .IN1(n2060), .IN2(n19048), .IN3(n1974), .IN4(n19032), .Q(
        n8633) );
  NAND4X0 U27673 ( .IN1(n8627), .IN2(n8628), .IN3(n8629), .IN4(n8630), .QN(
        s10_data_o[26]) );
  OA22X1 U27674 ( .IN1(n1715), .IN2(n18979), .IN3(n1610), .IN4(n18968), .Q(
        n8627) );
  OA22X1 U27675 ( .IN1(n1887), .IN2(n19012), .IN3(n1801), .IN4(n19003), .Q(
        n8628) );
  OA22X1 U27676 ( .IN1(n2059), .IN2(n19045), .IN3(n1973), .IN4(n19032), .Q(
        n8629) );
  NAND4X0 U27677 ( .IN1(n8623), .IN2(n8624), .IN3(n8625), .IN4(n8626), .QN(
        s10_data_o[27]) );
  OA22X1 U27678 ( .IN1(n1714), .IN2(n18983), .IN3(n1609), .IN4(n18971), .Q(
        n8623) );
  OA22X1 U27679 ( .IN1(n1886), .IN2(n19015), .IN3(n1800), .IN4(n19002), .Q(
        n8624) );
  OA22X1 U27680 ( .IN1(n2058), .IN2(n19049), .IN3(n1972), .IN4(n19033), .Q(
        n8625) );
  NAND4X0 U27681 ( .IN1(n8619), .IN2(n8620), .IN3(n8621), .IN4(n8622), .QN(
        s10_data_o[28]) );
  OA22X1 U27682 ( .IN1(n1713), .IN2(n18983), .IN3(n1608), .IN4(n18968), .Q(
        n8619) );
  OA22X1 U27683 ( .IN1(n1885), .IN2(n8543), .IN3(n1799), .IN4(n19003), .Q(
        n8620) );
  OA22X1 U27684 ( .IN1(n2057), .IN2(n19048), .IN3(n1971), .IN4(n19033), .Q(
        n8621) );
  NAND4X0 U27685 ( .IN1(n8615), .IN2(n8616), .IN3(n8617), .IN4(n8618), .QN(
        s10_data_o[29]) );
  OA22X1 U27686 ( .IN1(n1712), .IN2(n18977), .IN3(n1607), .IN4(n18970), .Q(
        n8615) );
  OA22X1 U27687 ( .IN1(n1884), .IN2(n8543), .IN3(n1798), .IN4(n19002), .Q(
        n8616) );
  OA22X1 U27688 ( .IN1(n2056), .IN2(n19045), .IN3(n1970), .IN4(n19033), .Q(
        n8617) );
  NAND4X0 U27689 ( .IN1(n8607), .IN2(n8608), .IN3(n8609), .IN4(n8610), .QN(
        s10_data_o[30]) );
  OA22X1 U27690 ( .IN1(n1711), .IN2(n18980), .IN3(n1606), .IN4(n18969), .Q(
        n8607) );
  OA22X1 U27691 ( .IN1(n1883), .IN2(n8543), .IN3(n1797), .IN4(n19004), .Q(
        n8608) );
  OA22X1 U27692 ( .IN1(n2055), .IN2(n19049), .IN3(n1969), .IN4(n19034), .Q(
        n8609) );
  NAND4X0 U27693 ( .IN1(n8603), .IN2(n8604), .IN3(n8605), .IN4(n8606), .QN(
        s10_data_o[31]) );
  OA22X1 U27694 ( .IN1(n1710), .IN2(n18978), .IN3(n1605), .IN4(n18969), .Q(
        n8603) );
  OA22X1 U27695 ( .IN1(n1882), .IN2(n19017), .IN3(n1796), .IN4(n19004), .Q(
        n8604) );
  OA22X1 U27696 ( .IN1(n2054), .IN2(n19044), .IN3(n1968), .IN4(n19034), .Q(
        n8605) );
  NAND4X0 U27697 ( .IN1(n4515), .IN2(n4516), .IN3(n4517), .IN4(n4518), .QN(
        s9_stb_o) );
  OA22X1 U27698 ( .IN1(n4525), .IN2(n1795), .IN3(n4526), .IN4(n1709), .Q(n4515) );
  OA22X1 U27699 ( .IN1(n4523), .IN2(n1967), .IN3(n4524), .IN4(n1881), .Q(n4516) );
  OA22X1 U27700 ( .IN1(n4521), .IN2(n2139), .IN3(n4522), .IN4(n2053), .Q(n4517) );
  NAND4X0 U27701 ( .IN1(n4503), .IN2(n4504), .IN3(n4505), .IN4(n4506), .QN(
        s9_we_o) );
  OA22X1 U27702 ( .IN1(n20813), .IN2(n1794), .IN3(n20799), .IN4(n1708), .Q(
        n4503) );
  OA22X1 U27703 ( .IN1(n20831), .IN2(n1966), .IN3(n20817), .IN4(n1880), .Q(
        n4504) );
  OA22X1 U27704 ( .IN1(n20849), .IN2(n2138), .IN3(n20835), .IN4(n2052), .Q(
        n4505) );
  NAND4X0 U27705 ( .IN1(n4539), .IN2(n4540), .IN3(n4541), .IN4(n4542), .QN(
        s9_sel_o[0]) );
  OA22X1 U27706 ( .IN1(n20815), .IN2(n1793), .IN3(n4514), .IN4(n1707), .Q(
        n4539) );
  OA22X1 U27707 ( .IN1(n20833), .IN2(n1965), .IN3(n4512), .IN4(n1879), .Q(
        n4540) );
  OA22X1 U27708 ( .IN1(n20851), .IN2(n2137), .IN3(n4510), .IN4(n2051), .Q(
        n4541) );
  NAND4X0 U27709 ( .IN1(n4535), .IN2(n4536), .IN3(n4537), .IN4(n4538), .QN(
        s9_sel_o[1]) );
  OA22X1 U27710 ( .IN1(n20815), .IN2(n1792), .IN3(n4514), .IN4(n1706), .Q(
        n4535) );
  OA22X1 U27711 ( .IN1(n20833), .IN2(n1964), .IN3(n4512), .IN4(n1878), .Q(
        n4536) );
  OA22X1 U27712 ( .IN1(n20851), .IN2(n2136), .IN3(n4510), .IN4(n2050), .Q(
        n4537) );
  NAND4X0 U27713 ( .IN1(n4531), .IN2(n4532), .IN3(n4533), .IN4(n4534), .QN(
        s9_sel_o[2]) );
  OA22X1 U27714 ( .IN1(n20815), .IN2(n1791), .IN3(n4514), .IN4(n1705), .Q(
        n4531) );
  OA22X1 U27715 ( .IN1(n20833), .IN2(n1963), .IN3(n4512), .IN4(n1877), .Q(
        n4532) );
  OA22X1 U27716 ( .IN1(n20851), .IN2(n2135), .IN3(n4510), .IN4(n2049), .Q(
        n4533) );
  NAND4X0 U27717 ( .IN1(n4527), .IN2(n4528), .IN3(n4529), .IN4(n4530), .QN(
        s9_sel_o[3]) );
  OA22X1 U27718 ( .IN1(n20815), .IN2(n1790), .IN3(n4514), .IN4(n1704), .Q(
        n4527) );
  OA22X1 U27719 ( .IN1(n20833), .IN2(n1962), .IN3(n4512), .IN4(n1876), .Q(
        n4528) );
  OA22X1 U27720 ( .IN1(n20851), .IN2(n2134), .IN3(n4510), .IN4(n2048), .Q(
        n4529) );
  NAND4X0 U27721 ( .IN1(n4795), .IN2(n4796), .IN3(n4797), .IN4(n4798), .QN(
        s9_addr_o[0]) );
  OA22X1 U27722 ( .IN1(n20808), .IN2(n1789), .IN3(n20799), .IN4(n1703), .Q(
        n4795) );
  OA22X1 U27723 ( .IN1(n20826), .IN2(n1961), .IN3(n20817), .IN4(n1875), .Q(
        n4796) );
  OA22X1 U27724 ( .IN1(n20844), .IN2(n2133), .IN3(n20835), .IN4(n2047), .Q(
        n4797) );
  NAND4X0 U27725 ( .IN1(n4751), .IN2(n4752), .IN3(n4753), .IN4(n4754), .QN(
        s9_addr_o[1]) );
  OA22X1 U27726 ( .IN1(n20810), .IN2(n1788), .IN3(n20801), .IN4(n1702), .Q(
        n4751) );
  OA22X1 U27727 ( .IN1(n20828), .IN2(n1960), .IN3(n20819), .IN4(n1874), .Q(
        n4752) );
  OA22X1 U27728 ( .IN1(n20846), .IN2(n2132), .IN3(n20837), .IN4(n2046), .Q(
        n4753) );
  NAND4X0 U27729 ( .IN1(n4707), .IN2(n4708), .IN3(n4709), .IN4(n4710), .QN(
        s9_addr_o[2]) );
  OA22X1 U27730 ( .IN1(n20813), .IN2(n1787), .IN3(n20804), .IN4(n1701), .Q(
        n4707) );
  OA22X1 U27731 ( .IN1(n20831), .IN2(n1959), .IN3(n20822), .IN4(n1873), .Q(
        n4708) );
  OA22X1 U27732 ( .IN1(n20849), .IN2(n2131), .IN3(n20840), .IN4(n2045), .Q(
        n4709) );
  NAND4X0 U27733 ( .IN1(n4695), .IN2(n4696), .IN3(n4697), .IN4(n4698), .QN(
        s9_addr_o[3]) );
  OA22X1 U27734 ( .IN1(n20812), .IN2(n1786), .IN3(n4514), .IN4(n1699), .Q(
        n4695) );
  OA22X1 U27735 ( .IN1(n20830), .IN2(n1958), .IN3(n4512), .IN4(n1872), .Q(
        n4696) );
  OA22X1 U27736 ( .IN1(n20848), .IN2(n2130), .IN3(n4510), .IN4(n2044), .Q(
        n4697) );
  NAND4X0 U27737 ( .IN1(n4691), .IN2(n4692), .IN3(n4693), .IN4(n4694), .QN(
        s9_addr_o[4]) );
  OA22X1 U27738 ( .IN1(n20812), .IN2(n1785), .IN3(n20802), .IN4(n1697), .Q(
        n4691) );
  OA22X1 U27739 ( .IN1(n20830), .IN2(n1957), .IN3(n20820), .IN4(n1871), .Q(
        n4692) );
  OA22X1 U27740 ( .IN1(n20848), .IN2(n2129), .IN3(n20838), .IN4(n2043), .Q(
        n4693) );
  NAND4X0 U27741 ( .IN1(n4687), .IN2(n4688), .IN3(n4689), .IN4(n4690), .QN(
        s9_addr_o[5]) );
  OA22X1 U27742 ( .IN1(n20812), .IN2(n1784), .IN3(n4514), .IN4(n1696), .Q(
        n4687) );
  OA22X1 U27743 ( .IN1(n20830), .IN2(n1956), .IN3(n4512), .IN4(n1870), .Q(
        n4688) );
  OA22X1 U27744 ( .IN1(n20848), .IN2(n2128), .IN3(n4510), .IN4(n2042), .Q(
        n4689) );
  NAND4X0 U27745 ( .IN1(n4683), .IN2(n4684), .IN3(n4685), .IN4(n4686), .QN(
        s9_addr_o[6]) );
  OA22X1 U27746 ( .IN1(n20813), .IN2(n1783), .IN3(n20803), .IN4(n1679), .Q(
        n4683) );
  OA22X1 U27747 ( .IN1(n20831), .IN2(n1955), .IN3(n20821), .IN4(n1869), .Q(
        n4684) );
  OA22X1 U27748 ( .IN1(n20849), .IN2(n2127), .IN3(n20839), .IN4(n2041), .Q(
        n4685) );
  NAND4X0 U27749 ( .IN1(n4679), .IN2(n4680), .IN3(n4681), .IN4(n4682), .QN(
        s9_addr_o[7]) );
  OA22X1 U27750 ( .IN1(n20813), .IN2(n1782), .IN3(n20803), .IN4(n1678), .Q(
        n4679) );
  OA22X1 U27751 ( .IN1(n20831), .IN2(n1954), .IN3(n20821), .IN4(n1868), .Q(
        n4680) );
  OA22X1 U27752 ( .IN1(n20849), .IN2(n2126), .IN3(n20839), .IN4(n2040), .Q(
        n4681) );
  NAND4X0 U27753 ( .IN1(n4675), .IN2(n4676), .IN3(n4677), .IN4(n4678), .QN(
        s9_addr_o[8]) );
  OA22X1 U27754 ( .IN1(n20813), .IN2(n1781), .IN3(n20803), .IN4(n1677), .Q(
        n4675) );
  OA22X1 U27755 ( .IN1(n20831), .IN2(n1953), .IN3(n20821), .IN4(n1867), .Q(
        n4676) );
  OA22X1 U27756 ( .IN1(n20849), .IN2(n2125), .IN3(n20839), .IN4(n2039), .Q(
        n4677) );
  NAND4X0 U27757 ( .IN1(n4671), .IN2(n4672), .IN3(n4673), .IN4(n4674), .QN(
        s9_addr_o[9]) );
  OA22X1 U27758 ( .IN1(n20813), .IN2(n1780), .IN3(n20803), .IN4(n1676), .Q(
        n4671) );
  OA22X1 U27759 ( .IN1(n20831), .IN2(n1952), .IN3(n20821), .IN4(n1866), .Q(
        n4672) );
  OA22X1 U27760 ( .IN1(n20849), .IN2(n2124), .IN3(n20839), .IN4(n2038), .Q(
        n4673) );
  NAND4X0 U27761 ( .IN1(n4791), .IN2(n4792), .IN3(n4793), .IN4(n4794), .QN(
        s9_addr_o[10]) );
  OA22X1 U27762 ( .IN1(n20808), .IN2(n1779), .IN3(n20799), .IN4(n1675), .Q(
        n4791) );
  OA22X1 U27763 ( .IN1(n20826), .IN2(n1951), .IN3(n20817), .IN4(n1865), .Q(
        n4792) );
  OA22X1 U27764 ( .IN1(n20844), .IN2(n2123), .IN3(n20835), .IN4(n2037), .Q(
        n4793) );
  NAND4X0 U27765 ( .IN1(n4787), .IN2(n4788), .IN3(n4789), .IN4(n4790), .QN(
        s9_addr_o[11]) );
  OA22X1 U27766 ( .IN1(n20808), .IN2(n1778), .IN3(n20799), .IN4(n1674), .Q(
        n4787) );
  OA22X1 U27767 ( .IN1(n20826), .IN2(n1950), .IN3(n20817), .IN4(n1864), .Q(
        n4788) );
  OA22X1 U27768 ( .IN1(n20844), .IN2(n2122), .IN3(n20835), .IN4(n2036), .Q(
        n4789) );
  NAND4X0 U27769 ( .IN1(n4783), .IN2(n4784), .IN3(n4785), .IN4(n4786), .QN(
        s9_addr_o[12]) );
  OA22X1 U27770 ( .IN1(n20808), .IN2(n1777), .IN3(n20799), .IN4(n1673), .Q(
        n4783) );
  OA22X1 U27771 ( .IN1(n20826), .IN2(n1949), .IN3(n20817), .IN4(n1863), .Q(
        n4784) );
  OA22X1 U27772 ( .IN1(n20844), .IN2(n2121), .IN3(n20835), .IN4(n2035), .Q(
        n4785) );
  NAND4X0 U27773 ( .IN1(n4779), .IN2(n4780), .IN3(n4781), .IN4(n4782), .QN(
        s9_addr_o[13]) );
  OA22X1 U27774 ( .IN1(n20809), .IN2(n1776), .IN3(n20800), .IN4(n1672), .Q(
        n4779) );
  OA22X1 U27775 ( .IN1(n20827), .IN2(n1948), .IN3(n20818), .IN4(n1862), .Q(
        n4780) );
  OA22X1 U27776 ( .IN1(n20845), .IN2(n2120), .IN3(n20836), .IN4(n2034), .Q(
        n4781) );
  NAND4X0 U27777 ( .IN1(n4775), .IN2(n4776), .IN3(n4777), .IN4(n4778), .QN(
        s9_addr_o[14]) );
  OA22X1 U27778 ( .IN1(n20809), .IN2(n1775), .IN3(n20800), .IN4(n1671), .Q(
        n4775) );
  OA22X1 U27779 ( .IN1(n20827), .IN2(n1947), .IN3(n20818), .IN4(n1861), .Q(
        n4776) );
  OA22X1 U27780 ( .IN1(n20845), .IN2(n2119), .IN3(n20836), .IN4(n2033), .Q(
        n4777) );
  NAND4X0 U27781 ( .IN1(n4771), .IN2(n4772), .IN3(n4773), .IN4(n4774), .QN(
        s9_addr_o[15]) );
  OA22X1 U27782 ( .IN1(n20809), .IN2(n1774), .IN3(n20800), .IN4(n1670), .Q(
        n4771) );
  OA22X1 U27783 ( .IN1(n20827), .IN2(n1946), .IN3(n20818), .IN4(n1860), .Q(
        n4772) );
  OA22X1 U27784 ( .IN1(n20845), .IN2(n2118), .IN3(n20836), .IN4(n2032), .Q(
        n4773) );
  NAND4X0 U27785 ( .IN1(n4767), .IN2(n4768), .IN3(n4769), .IN4(n4770), .QN(
        s9_addr_o[16]) );
  OA22X1 U27786 ( .IN1(n20809), .IN2(n1773), .IN3(n20800), .IN4(n1669), .Q(
        n4767) );
  OA22X1 U27787 ( .IN1(n20827), .IN2(n1945), .IN3(n20818), .IN4(n1859), .Q(
        n4768) );
  OA22X1 U27788 ( .IN1(n20845), .IN2(n2117), .IN3(n20836), .IN4(n2031), .Q(
        n4769) );
  NAND4X0 U27789 ( .IN1(n4763), .IN2(n4764), .IN3(n4765), .IN4(n4766), .QN(
        s9_addr_o[17]) );
  OA22X1 U27790 ( .IN1(n20810), .IN2(n1772), .IN3(n20801), .IN4(n1668), .Q(
        n4763) );
  OA22X1 U27791 ( .IN1(n20828), .IN2(n1944), .IN3(n20819), .IN4(n1858), .Q(
        n4764) );
  OA22X1 U27792 ( .IN1(n20846), .IN2(n2116), .IN3(n20837), .IN4(n2030), .Q(
        n4765) );
  NAND4X0 U27793 ( .IN1(n4759), .IN2(n4760), .IN3(n4761), .IN4(n4762), .QN(
        s9_addr_o[18]) );
  OA22X1 U27794 ( .IN1(n20810), .IN2(n1771), .IN3(n20801), .IN4(n1667), .Q(
        n4759) );
  OA22X1 U27795 ( .IN1(n20828), .IN2(n1943), .IN3(n20819), .IN4(n1857), .Q(
        n4760) );
  OA22X1 U27796 ( .IN1(n20846), .IN2(n2115), .IN3(n20837), .IN4(n2029), .Q(
        n4761) );
  NAND4X0 U27797 ( .IN1(n4755), .IN2(n4756), .IN3(n4757), .IN4(n4758), .QN(
        s9_addr_o[19]) );
  OA22X1 U27798 ( .IN1(n20810), .IN2(n1770), .IN3(n20801), .IN4(n1666), .Q(
        n4755) );
  OA22X1 U27799 ( .IN1(n20828), .IN2(n1942), .IN3(n20819), .IN4(n1856), .Q(
        n4756) );
  OA22X1 U27800 ( .IN1(n20846), .IN2(n2114), .IN3(n20837), .IN4(n2028), .Q(
        n4757) );
  NAND4X0 U27801 ( .IN1(n4747), .IN2(n4748), .IN3(n4749), .IN4(n4750), .QN(
        s9_addr_o[20]) );
  OA22X1 U27802 ( .IN1(n20815), .IN2(n1769), .IN3(n20800), .IN4(n1665), .Q(
        n4747) );
  OA22X1 U27803 ( .IN1(n20833), .IN2(n1941), .IN3(n20818), .IN4(n1855), .Q(
        n4748) );
  OA22X1 U27804 ( .IN1(n20851), .IN2(n2113), .IN3(n20836), .IN4(n2027), .Q(
        n4749) );
  NAND4X0 U27805 ( .IN1(n4743), .IN2(n4744), .IN3(n4745), .IN4(n4746), .QN(
        s9_addr_o[21]) );
  OA22X1 U27806 ( .IN1(n20808), .IN2(n1768), .IN3(n20800), .IN4(n1664), .Q(
        n4743) );
  OA22X1 U27807 ( .IN1(n20826), .IN2(n1940), .IN3(n20818), .IN4(n1854), .Q(
        n4744) );
  OA22X1 U27808 ( .IN1(n20844), .IN2(n2112), .IN3(n20836), .IN4(n2026), .Q(
        n4745) );
  NAND4X0 U27809 ( .IN1(n4739), .IN2(n4740), .IN3(n4741), .IN4(n4742), .QN(
        s9_addr_o[22]) );
  OA22X1 U27810 ( .IN1(n20809), .IN2(n1767), .IN3(n20799), .IN4(n1663), .Q(
        n4739) );
  OA22X1 U27811 ( .IN1(n20827), .IN2(n1939), .IN3(n20817), .IN4(n1853), .Q(
        n4740) );
  OA22X1 U27812 ( .IN1(n20845), .IN2(n2111), .IN3(n20835), .IN4(n2025), .Q(
        n4741) );
  NAND4X0 U27813 ( .IN1(n4735), .IN2(n4736), .IN3(n4737), .IN4(n4738), .QN(
        s9_addr_o[23]) );
  OA22X1 U27814 ( .IN1(n20815), .IN2(n1766), .IN3(n20800), .IN4(n1662), .Q(
        n4735) );
  OA22X1 U27815 ( .IN1(n20833), .IN2(n1938), .IN3(n20818), .IN4(n1852), .Q(
        n4736) );
  OA22X1 U27816 ( .IN1(n20851), .IN2(n2110), .IN3(n20836), .IN4(n2024), .Q(
        n4737) );
  NAND4X0 U27817 ( .IN1(n4731), .IN2(n4732), .IN3(n4733), .IN4(n4734), .QN(
        s9_addr_o[24]) );
  OA22X1 U27818 ( .IN1(n20811), .IN2(n1765), .IN3(n20802), .IN4(n1661), .Q(
        n4731) );
  OA22X1 U27819 ( .IN1(n20829), .IN2(n1937), .IN3(n20820), .IN4(n1851), .Q(
        n4732) );
  OA22X1 U27820 ( .IN1(n20847), .IN2(n2109), .IN3(n20838), .IN4(n2023), .Q(
        n4733) );
  NAND4X0 U27821 ( .IN1(n4727), .IN2(n4728), .IN3(n4729), .IN4(n4730), .QN(
        s9_addr_o[25]) );
  OA22X1 U27822 ( .IN1(n20811), .IN2(n1764), .IN3(n20802), .IN4(n1660), .Q(
        n4727) );
  OA22X1 U27823 ( .IN1(n20829), .IN2(n1936), .IN3(n20820), .IN4(n1850), .Q(
        n4728) );
  OA22X1 U27824 ( .IN1(n20847), .IN2(n2108), .IN3(n20838), .IN4(n2022), .Q(
        n4729) );
  NAND4X0 U27825 ( .IN1(n4723), .IN2(n4724), .IN3(n4725), .IN4(n4726), .QN(
        s9_addr_o[26]) );
  OA22X1 U27826 ( .IN1(n20811), .IN2(n1763), .IN3(n20802), .IN4(n1659), .Q(
        n4723) );
  OA22X1 U27827 ( .IN1(n20829), .IN2(n1935), .IN3(n20820), .IN4(n1849), .Q(
        n4724) );
  OA22X1 U27828 ( .IN1(n20847), .IN2(n2107), .IN3(n20838), .IN4(n2021), .Q(
        n4725) );
  NAND4X0 U27829 ( .IN1(n4719), .IN2(n4720), .IN3(n4721), .IN4(n4722), .QN(
        s9_addr_o[27]) );
  OA22X1 U27830 ( .IN1(n20811), .IN2(n1762), .IN3(n20802), .IN4(n1658), .Q(
        n4719) );
  OA22X1 U27831 ( .IN1(n20829), .IN2(n1934), .IN3(n20820), .IN4(n1848), .Q(
        n4720) );
  OA22X1 U27832 ( .IN1(n20847), .IN2(n2106), .IN3(n20838), .IN4(n2020), .Q(
        n4721) );
  NAND4X0 U27833 ( .IN1(n4715), .IN2(n4716), .IN3(n4717), .IN4(n4718), .QN(
        s9_addr_o[28]) );
  OA22X1 U27834 ( .IN1(n20811), .IN2(n1761), .IN3(n4514), .IN4(n1657), .Q(
        n4715) );
  OA22X1 U27835 ( .IN1(n20829), .IN2(n1933), .IN3(n4512), .IN4(n1847), .Q(
        n4716) );
  OA22X1 U27836 ( .IN1(n20847), .IN2(n2105), .IN3(n4510), .IN4(n2019), .Q(
        n4717) );
  NAND4X0 U27837 ( .IN1(n4711), .IN2(n4712), .IN3(n4713), .IN4(n4714), .QN(
        s9_addr_o[29]) );
  OA22X1 U27838 ( .IN1(n4513), .IN2(n1760), .IN3(n20801), .IN4(n1656), .Q(
        n4711) );
  OA22X1 U27839 ( .IN1(n4511), .IN2(n1932), .IN3(n20819), .IN4(n1846), .Q(
        n4712) );
  OA22X1 U27840 ( .IN1(n4509), .IN2(n2104), .IN3(n20837), .IN4(n2018), .Q(
        n4713) );
  NAND4X0 U27841 ( .IN1(n4703), .IN2(n4704), .IN3(n4705), .IN4(n4706), .QN(
        s9_addr_o[30]) );
  OA22X1 U27842 ( .IN1(n20810), .IN2(n1759), .IN3(n20806), .IN4(n1655), .Q(
        n4703) );
  OA22X1 U27843 ( .IN1(n20828), .IN2(n1931), .IN3(n20824), .IN4(n1845), .Q(
        n4704) );
  OA22X1 U27844 ( .IN1(n20846), .IN2(n2103), .IN3(n20842), .IN4(n2017), .Q(
        n4705) );
  NAND4X0 U27845 ( .IN1(n4699), .IN2(n4700), .IN3(n4701), .IN4(n4702), .QN(
        s9_addr_o[31]) );
  OA22X1 U27846 ( .IN1(n20812), .IN2(n1758), .IN3(n20803), .IN4(n1650), .Q(
        n4699) );
  OA22X1 U27847 ( .IN1(n20830), .IN2(n1930), .IN3(n20821), .IN4(n1844), .Q(
        n4700) );
  OA22X1 U27848 ( .IN1(n20848), .IN2(n2102), .IN3(n20839), .IN4(n2016), .Q(
        n4701) );
  NAND4X0 U27849 ( .IN1(n4667), .IN2(n4668), .IN3(n4669), .IN4(n4670), .QN(
        s9_data_o[0]) );
  OA22X1 U27850 ( .IN1(n4513), .IN2(n1741), .IN3(n20804), .IN4(n1636), .Q(
        n4667) );
  OA22X1 U27851 ( .IN1(n4511), .IN2(n1913), .IN3(n20822), .IN4(n1827), .Q(
        n4668) );
  OA22X1 U27852 ( .IN1(n4509), .IN2(n2085), .IN3(n20840), .IN4(n1999), .Q(
        n4669) );
  NAND4X0 U27853 ( .IN1(n4623), .IN2(n4624), .IN3(n4625), .IN4(n4626), .QN(
        s9_data_o[1]) );
  OA22X1 U27854 ( .IN1(n20808), .IN2(n1740), .IN3(n4514), .IN4(n1635), .Q(
        n4623) );
  OA22X1 U27855 ( .IN1(n20826), .IN2(n1912), .IN3(n4512), .IN4(n1826), .Q(
        n4624) );
  OA22X1 U27856 ( .IN1(n20844), .IN2(n2084), .IN3(n4510), .IN4(n1998), .Q(
        n4625) );
  NAND4X0 U27857 ( .IN1(n4579), .IN2(n4580), .IN3(n4581), .IN4(n4582), .QN(
        s9_data_o[2]) );
  OA22X1 U27858 ( .IN1(n4513), .IN2(n1739), .IN3(n20806), .IN4(n1634), .Q(
        n4579) );
  OA22X1 U27859 ( .IN1(n4511), .IN2(n1911), .IN3(n20824), .IN4(n1825), .Q(
        n4580) );
  OA22X1 U27860 ( .IN1(n4509), .IN2(n2083), .IN3(n20842), .IN4(n1997), .Q(
        n4581) );
  NAND4X0 U27861 ( .IN1(n4567), .IN2(n4568), .IN3(n4569), .IN4(n4570), .QN(
        s9_data_o[3]) );
  OA22X1 U27862 ( .IN1(n20812), .IN2(n1738), .IN3(n4514), .IN4(n1633), .Q(
        n4567) );
  OA22X1 U27863 ( .IN1(n20830), .IN2(n1910), .IN3(n4512), .IN4(n1824), .Q(
        n4568) );
  OA22X1 U27864 ( .IN1(n20848), .IN2(n2082), .IN3(n4510), .IN4(n1996), .Q(
        n4569) );
  NAND4X0 U27865 ( .IN1(n4563), .IN2(n4564), .IN3(n4565), .IN4(n4566), .QN(
        s9_data_o[4]) );
  OA22X1 U27866 ( .IN1(n20814), .IN2(n1737), .IN3(n20805), .IN4(n1632), .Q(
        n4563) );
  OA22X1 U27867 ( .IN1(n20832), .IN2(n1909), .IN3(n20823), .IN4(n1823), .Q(
        n4564) );
  OA22X1 U27868 ( .IN1(n20850), .IN2(n2081), .IN3(n20841), .IN4(n1995), .Q(
        n4565) );
  NAND4X0 U27869 ( .IN1(n4559), .IN2(n4560), .IN3(n4561), .IN4(n4562), .QN(
        s9_data_o[5]) );
  OA22X1 U27870 ( .IN1(n20812), .IN2(n1736), .IN3(n4514), .IN4(n1631), .Q(
        n4559) );
  OA22X1 U27871 ( .IN1(n20830), .IN2(n1908), .IN3(n4512), .IN4(n1822), .Q(
        n4560) );
  OA22X1 U27872 ( .IN1(n20848), .IN2(n2080), .IN3(n4510), .IN4(n1994), .Q(
        n4561) );
  NAND4X0 U27873 ( .IN1(n4555), .IN2(n4556), .IN3(n4557), .IN4(n4558), .QN(
        s9_data_o[6]) );
  OA22X1 U27874 ( .IN1(n20814), .IN2(n1735), .IN3(n20806), .IN4(n1630), .Q(
        n4555) );
  OA22X1 U27875 ( .IN1(n20832), .IN2(n1907), .IN3(n20824), .IN4(n1821), .Q(
        n4556) );
  OA22X1 U27876 ( .IN1(n20850), .IN2(n2079), .IN3(n20842), .IN4(n1993), .Q(
        n4557) );
  NAND4X0 U27877 ( .IN1(n4551), .IN2(n4552), .IN3(n4553), .IN4(n4554), .QN(
        s9_data_o[7]) );
  OA22X1 U27878 ( .IN1(n20814), .IN2(n1734), .IN3(n20806), .IN4(n1629), .Q(
        n4551) );
  OA22X1 U27879 ( .IN1(n20832), .IN2(n1906), .IN3(n20824), .IN4(n1820), .Q(
        n4552) );
  OA22X1 U27880 ( .IN1(n20850), .IN2(n2078), .IN3(n20842), .IN4(n1992), .Q(
        n4553) );
  NAND4X0 U27881 ( .IN1(n4547), .IN2(n4548), .IN3(n4549), .IN4(n4550), .QN(
        s9_data_o[8]) );
  OA22X1 U27882 ( .IN1(n20814), .IN2(n1733), .IN3(n20806), .IN4(n1628), .Q(
        n4547) );
  OA22X1 U27883 ( .IN1(n20832), .IN2(n1905), .IN3(n20824), .IN4(n1819), .Q(
        n4548) );
  OA22X1 U27884 ( .IN1(n20850), .IN2(n2077), .IN3(n20842), .IN4(n1991), .Q(
        n4549) );
  NAND4X0 U27885 ( .IN1(n4543), .IN2(n4544), .IN3(n4545), .IN4(n4546), .QN(
        s9_data_o[9]) );
  OA22X1 U27886 ( .IN1(n20814), .IN2(n1732), .IN3(n20806), .IN4(n1627), .Q(
        n4543) );
  OA22X1 U27887 ( .IN1(n20832), .IN2(n1904), .IN3(n20824), .IN4(n1818), .Q(
        n4544) );
  OA22X1 U27888 ( .IN1(n20850), .IN2(n2076), .IN3(n20842), .IN4(n1990), .Q(
        n4545) );
  NAND4X0 U27889 ( .IN1(n4663), .IN2(n4664), .IN3(n4665), .IN4(n4666), .QN(
        s9_data_o[10]) );
  OA22X1 U27890 ( .IN1(n4513), .IN2(n1731), .IN3(n20804), .IN4(n1626), .Q(
        n4663) );
  OA22X1 U27891 ( .IN1(n4511), .IN2(n1903), .IN3(n20822), .IN4(n1817), .Q(
        n4664) );
  OA22X1 U27892 ( .IN1(n4509), .IN2(n2075), .IN3(n20840), .IN4(n1989), .Q(
        n4665) );
  NAND4X0 U27893 ( .IN1(n4659), .IN2(n4660), .IN3(n4661), .IN4(n4662), .QN(
        s9_data_o[11]) );
  OA22X1 U27894 ( .IN1(n4513), .IN2(n1730), .IN3(n20804), .IN4(n1625), .Q(
        n4659) );
  OA22X1 U27895 ( .IN1(n4511), .IN2(n1902), .IN3(n20822), .IN4(n1816), .Q(
        n4660) );
  OA22X1 U27896 ( .IN1(n4509), .IN2(n2074), .IN3(n20840), .IN4(n1988), .Q(
        n4661) );
  NAND4X0 U27897 ( .IN1(n4655), .IN2(n4656), .IN3(n4657), .IN4(n4658), .QN(
        s9_data_o[12]) );
  OA22X1 U27898 ( .IN1(n4513), .IN2(n1729), .IN3(n20804), .IN4(n1624), .Q(
        n4655) );
  OA22X1 U27899 ( .IN1(n4511), .IN2(n1901), .IN3(n20822), .IN4(n1815), .Q(
        n4656) );
  OA22X1 U27900 ( .IN1(n4509), .IN2(n2073), .IN3(n20840), .IN4(n1987), .Q(
        n4657) );
  NAND4X0 U27901 ( .IN1(n4651), .IN2(n4652), .IN3(n4653), .IN4(n4654), .QN(
        s9_data_o[13]) );
  OA22X1 U27902 ( .IN1(n4513), .IN2(n1728), .IN3(n20805), .IN4(n1623), .Q(
        n4651) );
  OA22X1 U27903 ( .IN1(n4511), .IN2(n1900), .IN3(n20823), .IN4(n1814), .Q(
        n4652) );
  OA22X1 U27904 ( .IN1(n4509), .IN2(n2072), .IN3(n20841), .IN4(n1986), .Q(
        n4653) );
  NAND4X0 U27905 ( .IN1(n4647), .IN2(n4648), .IN3(n4649), .IN4(n4650), .QN(
        s9_data_o[14]) );
  OA22X1 U27906 ( .IN1(n4513), .IN2(n1727), .IN3(n20805), .IN4(n1622), .Q(
        n4647) );
  OA22X1 U27907 ( .IN1(n4511), .IN2(n1899), .IN3(n20823), .IN4(n1813), .Q(
        n4648) );
  OA22X1 U27908 ( .IN1(n4509), .IN2(n2071), .IN3(n20841), .IN4(n1985), .Q(
        n4649) );
  NAND4X0 U27909 ( .IN1(n4643), .IN2(n4644), .IN3(n4645), .IN4(n4646), .QN(
        s9_data_o[15]) );
  OA22X1 U27910 ( .IN1(n4513), .IN2(n1726), .IN3(n20805), .IN4(n1621), .Q(
        n4643) );
  OA22X1 U27911 ( .IN1(n4511), .IN2(n1898), .IN3(n20823), .IN4(n1812), .Q(
        n4644) );
  OA22X1 U27912 ( .IN1(n4509), .IN2(n2070), .IN3(n20841), .IN4(n1984), .Q(
        n4645) );
  NAND4X0 U27913 ( .IN1(n4639), .IN2(n4640), .IN3(n4641), .IN4(n4642), .QN(
        s9_data_o[16]) );
  OA22X1 U27914 ( .IN1(n4513), .IN2(n1725), .IN3(n20805), .IN4(n1620), .Q(
        n4639) );
  OA22X1 U27915 ( .IN1(n4511), .IN2(n1897), .IN3(n20823), .IN4(n1811), .Q(
        n4640) );
  OA22X1 U27916 ( .IN1(n4509), .IN2(n2069), .IN3(n20841), .IN4(n1983), .Q(
        n4641) );
  NAND4X0 U27917 ( .IN1(n4635), .IN2(n4636), .IN3(n4637), .IN4(n4638), .QN(
        s9_data_o[17]) );
  OA22X1 U27918 ( .IN1(n20809), .IN2(n1724), .IN3(n4514), .IN4(n1619), .Q(
        n4635) );
  OA22X1 U27919 ( .IN1(n20827), .IN2(n1896), .IN3(n4512), .IN4(n1810), .Q(
        n4636) );
  OA22X1 U27920 ( .IN1(n20845), .IN2(n2068), .IN3(n4510), .IN4(n1982), .Q(
        n4637) );
  NAND4X0 U27921 ( .IN1(n4631), .IN2(n4632), .IN3(n4633), .IN4(n4634), .QN(
        s9_data_o[18]) );
  OA22X1 U27922 ( .IN1(n20811), .IN2(n1723), .IN3(n4514), .IN4(n1618), .Q(
        n4631) );
  OA22X1 U27923 ( .IN1(n20829), .IN2(n1895), .IN3(n4512), .IN4(n1809), .Q(
        n4632) );
  OA22X1 U27924 ( .IN1(n20847), .IN2(n2067), .IN3(n4510), .IN4(n1981), .Q(
        n4633) );
  NAND4X0 U27925 ( .IN1(n4627), .IN2(n4628), .IN3(n4629), .IN4(n4630), .QN(
        s9_data_o[19]) );
  OA22X1 U27926 ( .IN1(n20810), .IN2(n1722), .IN3(n4514), .IN4(n1617), .Q(
        n4627) );
  OA22X1 U27927 ( .IN1(n20828), .IN2(n1894), .IN3(n4512), .IN4(n1808), .Q(
        n4628) );
  OA22X1 U27928 ( .IN1(n20846), .IN2(n2066), .IN3(n4510), .IN4(n1980), .Q(
        n4629) );
  NAND4X0 U27929 ( .IN1(n4619), .IN2(n4620), .IN3(n4621), .IN4(n4622), .QN(
        s9_data_o[20]) );
  OA22X1 U27930 ( .IN1(n20813), .IN2(n1721), .IN3(n20802), .IN4(n1616), .Q(
        n4619) );
  OA22X1 U27931 ( .IN1(n20831), .IN2(n1893), .IN3(n20820), .IN4(n1807), .Q(
        n4620) );
  OA22X1 U27932 ( .IN1(n20849), .IN2(n2065), .IN3(n20838), .IN4(n1979), .Q(
        n4621) );
  NAND4X0 U27933 ( .IN1(n4615), .IN2(n4616), .IN3(n4617), .IN4(n4618), .QN(
        s9_data_o[21]) );
  OA22X1 U27934 ( .IN1(n20808), .IN2(n1720), .IN3(n20805), .IN4(n1615), .Q(
        n4615) );
  OA22X1 U27935 ( .IN1(n20826), .IN2(n1892), .IN3(n20823), .IN4(n1806), .Q(
        n4616) );
  OA22X1 U27936 ( .IN1(n20844), .IN2(n2064), .IN3(n20841), .IN4(n1978), .Q(
        n4617) );
  NAND4X0 U27937 ( .IN1(n4611), .IN2(n4612), .IN3(n4613), .IN4(n4614), .QN(
        s9_data_o[22]) );
  OA22X1 U27938 ( .IN1(n20809), .IN2(n1719), .IN3(n20802), .IN4(n1614), .Q(
        n4611) );
  OA22X1 U27939 ( .IN1(n20827), .IN2(n1891), .IN3(n20820), .IN4(n1805), .Q(
        n4612) );
  OA22X1 U27940 ( .IN1(n20845), .IN2(n2063), .IN3(n20838), .IN4(n1977), .Q(
        n4613) );
  NAND4X0 U27941 ( .IN1(n4607), .IN2(n4608), .IN3(n4609), .IN4(n4610), .QN(
        s9_data_o[23]) );
  OA22X1 U27942 ( .IN1(n4513), .IN2(n1718), .IN3(n20799), .IN4(n1613), .Q(
        n4607) );
  OA22X1 U27943 ( .IN1(n4511), .IN2(n1890), .IN3(n20817), .IN4(n1804), .Q(
        n4608) );
  OA22X1 U27944 ( .IN1(n4509), .IN2(n2062), .IN3(n20835), .IN4(n1976), .Q(
        n4609) );
  NAND4X0 U27945 ( .IN1(n4603), .IN2(n4604), .IN3(n4605), .IN4(n4606), .QN(
        s9_data_o[24]) );
  OA22X1 U27946 ( .IN1(n20811), .IN2(n1717), .IN3(n20806), .IN4(n1612), .Q(
        n4603) );
  OA22X1 U27947 ( .IN1(n20829), .IN2(n1889), .IN3(n20824), .IN4(n1803), .Q(
        n4604) );
  OA22X1 U27948 ( .IN1(n20847), .IN2(n2061), .IN3(n20842), .IN4(n1975), .Q(
        n4605) );
  NAND4X0 U27949 ( .IN1(n4599), .IN2(n4600), .IN3(n4601), .IN4(n4602), .QN(
        s9_data_o[25]) );
  OA22X1 U27950 ( .IN1(n20810), .IN2(n1716), .IN3(n20803), .IN4(n1611), .Q(
        n4599) );
  OA22X1 U27951 ( .IN1(n20828), .IN2(n1888), .IN3(n20821), .IN4(n1802), .Q(
        n4600) );
  OA22X1 U27952 ( .IN1(n20846), .IN2(n2060), .IN3(n20839), .IN4(n1974), .Q(
        n4601) );
  NAND4X0 U27953 ( .IN1(n4595), .IN2(n4596), .IN3(n4597), .IN4(n4598), .QN(
        s9_data_o[26]) );
  OA22X1 U27954 ( .IN1(n4513), .IN2(n1715), .IN3(n20801), .IN4(n1610), .Q(
        n4595) );
  OA22X1 U27955 ( .IN1(n4511), .IN2(n1887), .IN3(n20819), .IN4(n1801), .Q(
        n4596) );
  OA22X1 U27956 ( .IN1(n4509), .IN2(n2059), .IN3(n20837), .IN4(n1973), .Q(
        n4597) );
  NAND4X0 U27957 ( .IN1(n4591), .IN2(n4592), .IN3(n4593), .IN4(n4594), .QN(
        s9_data_o[27]) );
  OA22X1 U27958 ( .IN1(n20815), .IN2(n1714), .IN3(n20804), .IN4(n1609), .Q(
        n4591) );
  OA22X1 U27959 ( .IN1(n20833), .IN2(n1886), .IN3(n20822), .IN4(n1800), .Q(
        n4592) );
  OA22X1 U27960 ( .IN1(n20851), .IN2(n2058), .IN3(n20840), .IN4(n1972), .Q(
        n4593) );
  NAND4X0 U27961 ( .IN1(n4587), .IN2(n4588), .IN3(n4589), .IN4(n4590), .QN(
        s9_data_o[28]) );
  OA22X1 U27962 ( .IN1(n20814), .IN2(n1713), .IN3(n20803), .IN4(n1608), .Q(
        n4587) );
  OA22X1 U27963 ( .IN1(n20832), .IN2(n1885), .IN3(n20821), .IN4(n1799), .Q(
        n4588) );
  OA22X1 U27964 ( .IN1(n20850), .IN2(n2057), .IN3(n20839), .IN4(n1971), .Q(
        n4589) );
  NAND4X0 U27965 ( .IN1(n4583), .IN2(n4584), .IN3(n4585), .IN4(n4586), .QN(
        s9_data_o[29]) );
  OA22X1 U27966 ( .IN1(n20814), .IN2(n1712), .IN3(n20801), .IN4(n1607), .Q(
        n4583) );
  OA22X1 U27967 ( .IN1(n20832), .IN2(n1884), .IN3(n20819), .IN4(n1798), .Q(
        n4584) );
  OA22X1 U27968 ( .IN1(n20850), .IN2(n2056), .IN3(n20837), .IN4(n1970), .Q(
        n4585) );
  NAND4X0 U27969 ( .IN1(n4575), .IN2(n4576), .IN3(n4577), .IN4(n4578), .QN(
        s9_data_o[30]) );
  OA22X1 U27970 ( .IN1(n20812), .IN2(n1711), .IN3(n20804), .IN4(n1606), .Q(
        n4575) );
  OA22X1 U27971 ( .IN1(n20830), .IN2(n1883), .IN3(n20822), .IN4(n1797), .Q(
        n4576) );
  OA22X1 U27972 ( .IN1(n20848), .IN2(n2055), .IN3(n20840), .IN4(n1969), .Q(
        n4577) );
  NAND4X0 U27973 ( .IN1(n4571), .IN2(n4572), .IN3(n4573), .IN4(n4574), .QN(
        s9_data_o[31]) );
  OA22X1 U27974 ( .IN1(n4513), .IN2(n1710), .IN3(n20805), .IN4(n1605), .Q(
        n4571) );
  OA22X1 U27975 ( .IN1(n4511), .IN2(n1882), .IN3(n20823), .IN4(n1796), .Q(
        n4572) );
  OA22X1 U27976 ( .IN1(n4509), .IN2(n2054), .IN3(n20841), .IN4(n1968), .Q(
        n4573) );
  NAND4X0 U27977 ( .IN1(n4811), .IN2(n4812), .IN3(n4813), .IN4(n4814), .QN(
        s8_stb_o) );
  OA22X1 U27978 ( .IN1(n1795), .IN2(n4821), .IN3(n1709), .IN4(n4822), .Q(n4811) );
  OA22X1 U27979 ( .IN1(n1967), .IN2(n4819), .IN3(n1881), .IN4(n4820), .Q(n4812) );
  OA22X1 U27980 ( .IN1(n2139), .IN2(n4817), .IN3(n2053), .IN4(n4818), .Q(n4813) );
  NAND4X0 U27981 ( .IN1(n4799), .IN2(n4800), .IN3(n4801), .IN4(n4802), .QN(
        s8_we_o) );
  OA22X1 U27982 ( .IN1(n1794), .IN2(n20691), .IN3(n1708), .IN4(n20685), .Q(
        n4799) );
  OA22X1 U27983 ( .IN1(n1966), .IN2(n20724), .IN3(n1880), .IN4(n20701), .Q(
        n4800) );
  OA22X1 U27984 ( .IN1(n2138), .IN2(n20757), .IN3(n2052), .IN4(n20751), .Q(
        n4801) );
  NAND4X0 U27985 ( .IN1(n4835), .IN2(n4836), .IN3(n4837), .IN4(n4838), .QN(
        s8_sel_o[0]) );
  OA22X1 U27986 ( .IN1(n1793), .IN2(n4809), .IN3(n1707), .IN4(n20683), .Q(
        n4835) );
  OA22X1 U27987 ( .IN1(n1965), .IN2(n20731), .IN3(n1879), .IN4(n20718), .Q(
        n4836) );
  OA22X1 U27988 ( .IN1(n2137), .IN2(n4805), .IN3(n2051), .IN4(n20749), .Q(
        n4837) );
  NAND4X0 U27989 ( .IN1(n4831), .IN2(n4832), .IN3(n4833), .IN4(n4834), .QN(
        s8_sel_o[1]) );
  OA22X1 U27990 ( .IN1(n1792), .IN2(n4809), .IN3(n1706), .IN4(n20683), .Q(
        n4831) );
  OA22X1 U27991 ( .IN1(n1964), .IN2(n20731), .IN3(n1878), .IN4(n20718), .Q(
        n4832) );
  OA22X1 U27992 ( .IN1(n2136), .IN2(n4805), .IN3(n2050), .IN4(n20749), .Q(
        n4833) );
  NAND4X0 U27993 ( .IN1(n4827), .IN2(n4828), .IN3(n4829), .IN4(n4830), .QN(
        s8_sel_o[2]) );
  OA22X1 U27994 ( .IN1(n1791), .IN2(n4809), .IN3(n1705), .IN4(n20685), .Q(
        n4827) );
  OA22X1 U27995 ( .IN1(n1963), .IN2(n20731), .IN3(n1877), .IN4(n20702), .Q(
        n4828) );
  OA22X1 U27996 ( .IN1(n2135), .IN2(n4805), .IN3(n2049), .IN4(n20751), .Q(
        n4829) );
  NAND4X0 U27997 ( .IN1(n4823), .IN2(n4824), .IN3(n4825), .IN4(n4826), .QN(
        s8_sel_o[3]) );
  OA22X1 U27998 ( .IN1(n1790), .IN2(n4809), .IN3(n1704), .IN4(n20685), .Q(
        n4823) );
  OA22X1 U27999 ( .IN1(n1962), .IN2(n20731), .IN3(n1876), .IN4(n20703), .Q(
        n4824) );
  OA22X1 U28000 ( .IN1(n2134), .IN2(n4805), .IN3(n2048), .IN4(n20751), .Q(
        n4825) );
  NAND4X0 U28001 ( .IN1(n5091), .IN2(n5092), .IN3(n5093), .IN4(n5094), .QN(
        s8_addr_o[0]) );
  OA22X1 U28002 ( .IN1(n1789), .IN2(n20691), .IN3(n1703), .IN4(n20668), .Q(
        n5091) );
  OA22X1 U28003 ( .IN1(n1961), .IN2(n20724), .IN3(n1875), .IN4(n20701), .Q(
        n5092) );
  OA22X1 U28004 ( .IN1(n2133), .IN2(n20757), .IN3(n2047), .IN4(n20734), .Q(
        n5093) );
  NAND4X0 U28005 ( .IN1(n5047), .IN2(n5048), .IN3(n5049), .IN4(n5050), .QN(
        s8_addr_o[1]) );
  OA22X1 U28006 ( .IN1(n1788), .IN2(n20693), .IN3(n1702), .IN4(n20671), .Q(
        n5047) );
  OA22X1 U28007 ( .IN1(n1960), .IN2(n20726), .IN3(n1874), .IN4(n20704), .Q(
        n5048) );
  OA22X1 U28008 ( .IN1(n2132), .IN2(n20759), .IN3(n2046), .IN4(n20737), .Q(
        n5049) );
  NAND4X0 U28009 ( .IN1(n5003), .IN2(n5004), .IN3(n5005), .IN4(n5006), .QN(
        s8_addr_o[2]) );
  OA22X1 U28010 ( .IN1(n1787), .IN2(n20691), .IN3(n1701), .IN4(n20675), .Q(
        n5003) );
  OA22X1 U28011 ( .IN1(n1959), .IN2(n20724), .IN3(n1873), .IN4(n20708), .Q(
        n5004) );
  OA22X1 U28012 ( .IN1(n2131), .IN2(n20757), .IN3(n2045), .IN4(n20741), .Q(
        n5005) );
  NAND4X0 U28013 ( .IN1(n4991), .IN2(n4992), .IN3(n4993), .IN4(n4994), .QN(
        s8_addr_o[3]) );
  OA22X1 U28014 ( .IN1(n1786), .IN2(n4809), .IN3(n1699), .IN4(n20676), .Q(
        n4991) );
  OA22X1 U28015 ( .IN1(n1958), .IN2(n20731), .IN3(n1872), .IN4(n20709), .Q(
        n4992) );
  OA22X1 U28016 ( .IN1(n2130), .IN2(n4805), .IN3(n2044), .IN4(n20742), .Q(
        n4993) );
  NAND4X0 U28017 ( .IN1(n4987), .IN2(n4988), .IN3(n4989), .IN4(n4990), .QN(
        s8_addr_o[4]) );
  OA22X1 U28018 ( .IN1(n1785), .IN2(n20694), .IN3(n1697), .IN4(n20676), .Q(
        n4987) );
  OA22X1 U28019 ( .IN1(n1957), .IN2(n20727), .IN3(n1871), .IN4(n20709), .Q(
        n4988) );
  OA22X1 U28020 ( .IN1(n2129), .IN2(n20760), .IN3(n2043), .IN4(n20742), .Q(
        n4989) );
  NAND4X0 U28021 ( .IN1(n4983), .IN2(n4984), .IN3(n4985), .IN4(n4986), .QN(
        s8_addr_o[5]) );
  OA22X1 U28022 ( .IN1(n1784), .IN2(n4809), .IN3(n1696), .IN4(n20677), .Q(
        n4983) );
  OA22X1 U28023 ( .IN1(n1956), .IN2(n20731), .IN3(n1870), .IN4(n20710), .Q(
        n4984) );
  OA22X1 U28024 ( .IN1(n2128), .IN2(n4805), .IN3(n2042), .IN4(n20743), .Q(
        n4985) );
  NAND4X0 U28025 ( .IN1(n4979), .IN2(n4980), .IN3(n4981), .IN4(n4982), .QN(
        s8_addr_o[6]) );
  OA22X1 U28026 ( .IN1(n1783), .IN2(n20695), .IN3(n1679), .IN4(n20677), .Q(
        n4979) );
  OA22X1 U28027 ( .IN1(n1955), .IN2(n20728), .IN3(n1869), .IN4(n20710), .Q(
        n4980) );
  OA22X1 U28028 ( .IN1(n2127), .IN2(n20761), .IN3(n2041), .IN4(n20743), .Q(
        n4981) );
  NAND4X0 U28029 ( .IN1(n4975), .IN2(n4976), .IN3(n4977), .IN4(n4978), .QN(
        s8_addr_o[7]) );
  OA22X1 U28030 ( .IN1(n1782), .IN2(n20695), .IN3(n1678), .IN4(n20677), .Q(
        n4975) );
  OA22X1 U28031 ( .IN1(n1954), .IN2(n20728), .IN3(n1868), .IN4(n20710), .Q(
        n4976) );
  OA22X1 U28032 ( .IN1(n2126), .IN2(n20761), .IN3(n2040), .IN4(n20743), .Q(
        n4977) );
  NAND4X0 U28033 ( .IN1(n4971), .IN2(n4972), .IN3(n4973), .IN4(n4974), .QN(
        s8_addr_o[8]) );
  OA22X1 U28034 ( .IN1(n1781), .IN2(n20695), .IN3(n1677), .IN4(n20678), .Q(
        n4971) );
  OA22X1 U28035 ( .IN1(n1953), .IN2(n20728), .IN3(n1867), .IN4(n20711), .Q(
        n4972) );
  OA22X1 U28036 ( .IN1(n2125), .IN2(n20761), .IN3(n2039), .IN4(n20744), .Q(
        n4973) );
  NAND4X0 U28037 ( .IN1(n4967), .IN2(n4968), .IN3(n4969), .IN4(n4970), .QN(
        s8_addr_o[9]) );
  OA22X1 U28038 ( .IN1(n1780), .IN2(n20695), .IN3(n1676), .IN4(n20678), .Q(
        n4967) );
  OA22X1 U28039 ( .IN1(n1952), .IN2(n20728), .IN3(n1866), .IN4(n20711), .Q(
        n4968) );
  OA22X1 U28040 ( .IN1(n2124), .IN2(n20761), .IN3(n2038), .IN4(n20744), .Q(
        n4969) );
  NAND4X0 U28041 ( .IN1(n5087), .IN2(n5088), .IN3(n5089), .IN4(n5090), .QN(
        s8_addr_o[10]) );
  OA22X1 U28042 ( .IN1(n1779), .IN2(n20691), .IN3(n1675), .IN4(n20668), .Q(
        n5087) );
  OA22X1 U28043 ( .IN1(n1951), .IN2(n20724), .IN3(n1865), .IN4(n20701), .Q(
        n5088) );
  OA22X1 U28044 ( .IN1(n2123), .IN2(n20757), .IN3(n2037), .IN4(n20734), .Q(
        n5089) );
  NAND4X0 U28045 ( .IN1(n5083), .IN2(n5084), .IN3(n5085), .IN4(n5086), .QN(
        s8_addr_o[11]) );
  OA22X1 U28046 ( .IN1(n1778), .IN2(n20691), .IN3(n1674), .IN4(n20668), .Q(
        n5083) );
  OA22X1 U28047 ( .IN1(n1950), .IN2(n20724), .IN3(n1864), .IN4(n20701), .Q(
        n5084) );
  OA22X1 U28048 ( .IN1(n2122), .IN2(n20757), .IN3(n2036), .IN4(n20734), .Q(
        n5085) );
  NAND4X0 U28049 ( .IN1(n5079), .IN2(n5080), .IN3(n5081), .IN4(n5082), .QN(
        s8_addr_o[12]) );
  OA22X1 U28050 ( .IN1(n1777), .IN2(n20691), .IN3(n1673), .IN4(n20669), .Q(
        n5079) );
  OA22X1 U28051 ( .IN1(n1949), .IN2(n20724), .IN3(n1863), .IN4(n20702), .Q(
        n5080) );
  OA22X1 U28052 ( .IN1(n2121), .IN2(n20757), .IN3(n2035), .IN4(n20735), .Q(
        n5081) );
  NAND4X0 U28053 ( .IN1(n5075), .IN2(n5076), .IN3(n5077), .IN4(n5078), .QN(
        s8_addr_o[13]) );
  OA22X1 U28054 ( .IN1(n1776), .IN2(n20692), .IN3(n1672), .IN4(n20669), .Q(
        n5075) );
  OA22X1 U28055 ( .IN1(n1948), .IN2(n20725), .IN3(n1862), .IN4(n20702), .Q(
        n5076) );
  OA22X1 U28056 ( .IN1(n2120), .IN2(n20758), .IN3(n2034), .IN4(n20735), .Q(
        n5077) );
  NAND4X0 U28057 ( .IN1(n5071), .IN2(n5072), .IN3(n5073), .IN4(n5074), .QN(
        s8_addr_o[14]) );
  OA22X1 U28058 ( .IN1(n1775), .IN2(n20692), .IN3(n1671), .IN4(n20669), .Q(
        n5071) );
  OA22X1 U28059 ( .IN1(n1947), .IN2(n20725), .IN3(n1861), .IN4(n20702), .Q(
        n5072) );
  OA22X1 U28060 ( .IN1(n2119), .IN2(n20758), .IN3(n2033), .IN4(n20735), .Q(
        n5073) );
  NAND4X0 U28061 ( .IN1(n5067), .IN2(n5068), .IN3(n5069), .IN4(n5070), .QN(
        s8_addr_o[15]) );
  OA22X1 U28062 ( .IN1(n1774), .IN2(n20692), .IN3(n1670), .IN4(n20670), .Q(
        n5067) );
  OA22X1 U28063 ( .IN1(n1946), .IN2(n20725), .IN3(n1860), .IN4(n20703), .Q(
        n5068) );
  OA22X1 U28064 ( .IN1(n2118), .IN2(n20758), .IN3(n2032), .IN4(n20736), .Q(
        n5069) );
  NAND4X0 U28065 ( .IN1(n5063), .IN2(n5064), .IN3(n5065), .IN4(n5066), .QN(
        s8_addr_o[16]) );
  OA22X1 U28066 ( .IN1(n1773), .IN2(n20692), .IN3(n1669), .IN4(n20670), .Q(
        n5063) );
  OA22X1 U28067 ( .IN1(n1945), .IN2(n20725), .IN3(n1859), .IN4(n20703), .Q(
        n5064) );
  OA22X1 U28068 ( .IN1(n2117), .IN2(n20758), .IN3(n2031), .IN4(n20736), .Q(
        n5065) );
  NAND4X0 U28069 ( .IN1(n5059), .IN2(n5060), .IN3(n5061), .IN4(n5062), .QN(
        s8_addr_o[17]) );
  OA22X1 U28070 ( .IN1(n1772), .IN2(n20693), .IN3(n1668), .IN4(n20670), .Q(
        n5059) );
  OA22X1 U28071 ( .IN1(n1944), .IN2(n20726), .IN3(n1858), .IN4(n20703), .Q(
        n5060) );
  OA22X1 U28072 ( .IN1(n2116), .IN2(n20759), .IN3(n2030), .IN4(n20736), .Q(
        n5061) );
  NAND4X0 U28073 ( .IN1(n5055), .IN2(n5056), .IN3(n5057), .IN4(n5058), .QN(
        s8_addr_o[18]) );
  OA22X1 U28074 ( .IN1(n1771), .IN2(n20693), .IN3(n1667), .IN4(n20671), .Q(
        n5055) );
  OA22X1 U28075 ( .IN1(n1943), .IN2(n20726), .IN3(n1857), .IN4(n20704), .Q(
        n5056) );
  OA22X1 U28076 ( .IN1(n2115), .IN2(n20759), .IN3(n2029), .IN4(n20737), .Q(
        n5057) );
  NAND4X0 U28077 ( .IN1(n5051), .IN2(n5052), .IN3(n5053), .IN4(n5054), .QN(
        s8_addr_o[19]) );
  OA22X1 U28078 ( .IN1(n1770), .IN2(n20693), .IN3(n1666), .IN4(n20671), .Q(
        n5051) );
  OA22X1 U28079 ( .IN1(n1942), .IN2(n20726), .IN3(n1856), .IN4(n20704), .Q(
        n5052) );
  OA22X1 U28080 ( .IN1(n2114), .IN2(n20759), .IN3(n2028), .IN4(n20737), .Q(
        n5053) );
  NAND4X0 U28081 ( .IN1(n5043), .IN2(n5044), .IN3(n5045), .IN4(n5046), .QN(
        s8_addr_o[20]) );
  OA22X1 U28082 ( .IN1(n1769), .IN2(n20692), .IN3(n1665), .IN4(n20672), .Q(
        n5043) );
  OA22X1 U28083 ( .IN1(n1941), .IN2(n20725), .IN3(n1855), .IN4(n20705), .Q(
        n5044) );
  OA22X1 U28084 ( .IN1(n2113), .IN2(n20758), .IN3(n2027), .IN4(n20738), .Q(
        n5045) );
  NAND4X0 U28085 ( .IN1(n5039), .IN2(n5040), .IN3(n5041), .IN4(n5042), .QN(
        s8_addr_o[21]) );
  OA22X1 U28086 ( .IN1(n1768), .IN2(n20692), .IN3(n1664), .IN4(n20672), .Q(
        n5039) );
  OA22X1 U28087 ( .IN1(n1940), .IN2(n20725), .IN3(n1854), .IN4(n20705), .Q(
        n5040) );
  OA22X1 U28088 ( .IN1(n2112), .IN2(n20758), .IN3(n2026), .IN4(n20738), .Q(
        n5041) );
  NAND4X0 U28089 ( .IN1(n5035), .IN2(n5036), .IN3(n5037), .IN4(n5038), .QN(
        s8_addr_o[22]) );
  OA22X1 U28090 ( .IN1(n1767), .IN2(n20691), .IN3(n1663), .IN4(n20672), .Q(
        n5035) );
  OA22X1 U28091 ( .IN1(n1939), .IN2(n20724), .IN3(n1853), .IN4(n20705), .Q(
        n5036) );
  OA22X1 U28092 ( .IN1(n2111), .IN2(n20757), .IN3(n2025), .IN4(n20738), .Q(
        n5037) );
  NAND4X0 U28093 ( .IN1(n5031), .IN2(n5032), .IN3(n5033), .IN4(n5034), .QN(
        s8_addr_o[23]) );
  OA22X1 U28094 ( .IN1(n1766), .IN2(n20692), .IN3(n1662), .IN4(n20673), .Q(
        n5031) );
  OA22X1 U28095 ( .IN1(n1938), .IN2(n20725), .IN3(n1852), .IN4(n20706), .Q(
        n5032) );
  OA22X1 U28096 ( .IN1(n2110), .IN2(n20758), .IN3(n2024), .IN4(n20739), .Q(
        n5033) );
  NAND4X0 U28097 ( .IN1(n5027), .IN2(n5028), .IN3(n5029), .IN4(n5030), .QN(
        s8_addr_o[24]) );
  OA22X1 U28098 ( .IN1(n1765), .IN2(n20694), .IN3(n1661), .IN4(n20673), .Q(
        n5027) );
  OA22X1 U28099 ( .IN1(n1937), .IN2(n20727), .IN3(n1851), .IN4(n20706), .Q(
        n5028) );
  OA22X1 U28100 ( .IN1(n2109), .IN2(n20760), .IN3(n2023), .IN4(n20739), .Q(
        n5029) );
  NAND4X0 U28101 ( .IN1(n5023), .IN2(n5024), .IN3(n5025), .IN4(n5026), .QN(
        s8_addr_o[25]) );
  OA22X1 U28102 ( .IN1(n1764), .IN2(n20694), .IN3(n1660), .IN4(n20673), .Q(
        n5023) );
  OA22X1 U28103 ( .IN1(n1936), .IN2(n20727), .IN3(n1850), .IN4(n20706), .Q(
        n5024) );
  OA22X1 U28104 ( .IN1(n2108), .IN2(n20760), .IN3(n2022), .IN4(n20739), .Q(
        n5025) );
  NAND4X0 U28105 ( .IN1(n5019), .IN2(n5020), .IN3(n5021), .IN4(n5022), .QN(
        s8_addr_o[26]) );
  OA22X1 U28106 ( .IN1(n1763), .IN2(n20694), .IN3(n1659), .IN4(n20674), .Q(
        n5019) );
  OA22X1 U28107 ( .IN1(n1935), .IN2(n20727), .IN3(n1849), .IN4(n20707), .Q(
        n5020) );
  OA22X1 U28108 ( .IN1(n2107), .IN2(n20760), .IN3(n2021), .IN4(n20740), .Q(
        n5021) );
  NAND4X0 U28109 ( .IN1(n5015), .IN2(n5016), .IN3(n5017), .IN4(n5018), .QN(
        s8_addr_o[27]) );
  OA22X1 U28110 ( .IN1(n1762), .IN2(n20694), .IN3(n1658), .IN4(n20674), .Q(
        n5015) );
  OA22X1 U28111 ( .IN1(n1934), .IN2(n20727), .IN3(n1848), .IN4(n20707), .Q(
        n5016) );
  OA22X1 U28112 ( .IN1(n2106), .IN2(n20760), .IN3(n2020), .IN4(n20740), .Q(
        n5017) );
  NAND4X0 U28113 ( .IN1(n5011), .IN2(n5012), .IN3(n5013), .IN4(n5014), .QN(
        s8_addr_o[28]) );
  OA22X1 U28114 ( .IN1(n1761), .IN2(n20694), .IN3(n1657), .IN4(n20674), .Q(
        n5011) );
  OA22X1 U28115 ( .IN1(n1933), .IN2(n20727), .IN3(n1847), .IN4(n20707), .Q(
        n5012) );
  OA22X1 U28116 ( .IN1(n2105), .IN2(n20760), .IN3(n2019), .IN4(n20740), .Q(
        n5013) );
  NAND4X0 U28117 ( .IN1(n5007), .IN2(n5008), .IN3(n5009), .IN4(n5010), .QN(
        s8_addr_o[29]) );
  OA22X1 U28118 ( .IN1(n1760), .IN2(n20693), .IN3(n1656), .IN4(n20675), .Q(
        n5007) );
  OA22X1 U28119 ( .IN1(n1932), .IN2(n20726), .IN3(n1846), .IN4(n20708), .Q(
        n5008) );
  OA22X1 U28120 ( .IN1(n2104), .IN2(n20761), .IN3(n2018), .IN4(n20741), .Q(
        n5009) );
  NAND4X0 U28121 ( .IN1(n4999), .IN2(n5000), .IN3(n5001), .IN4(n5002), .QN(
        s8_addr_o[30]) );
  OA22X1 U28122 ( .IN1(n1759), .IN2(n20694), .IN3(n1655), .IN4(n20675), .Q(
        n4999) );
  OA22X1 U28123 ( .IN1(n1931), .IN2(n20727), .IN3(n1845), .IN4(n20708), .Q(
        n5000) );
  OA22X1 U28124 ( .IN1(n2103), .IN2(n20760), .IN3(n2017), .IN4(n20741), .Q(
        n5001) );
  NAND4X0 U28125 ( .IN1(n4995), .IN2(n4996), .IN3(n4997), .IN4(n4998), .QN(
        s8_addr_o[31]) );
  OA22X1 U28126 ( .IN1(n1758), .IN2(n20695), .IN3(n1650), .IN4(n20676), .Q(
        n4995) );
  OA22X1 U28127 ( .IN1(n1930), .IN2(n20728), .IN3(n1844), .IN4(n20709), .Q(
        n4996) );
  OA22X1 U28128 ( .IN1(n2102), .IN2(n20764), .IN3(n2016), .IN4(n20742), .Q(
        n4997) );
  NAND4X0 U28129 ( .IN1(n4963), .IN2(n4964), .IN3(n4965), .IN4(n4966), .QN(
        s8_data_o[0]) );
  OA22X1 U28130 ( .IN1(n1741), .IN2(n20696), .IN3(n1636), .IN4(n20678), .Q(
        n4963) );
  OA22X1 U28131 ( .IN1(n1913), .IN2(n20729), .IN3(n1827), .IN4(n20711), .Q(
        n4964) );
  OA22X1 U28132 ( .IN1(n2085), .IN2(n20762), .IN3(n1999), .IN4(n20744), .Q(
        n4965) );
  NAND4X0 U28133 ( .IN1(n4919), .IN2(n4920), .IN3(n4921), .IN4(n4922), .QN(
        s8_data_o[1]) );
  OA22X1 U28134 ( .IN1(n1740), .IN2(n20698), .IN3(n1635), .IN4(n20680), .Q(
        n4919) );
  OA22X1 U28135 ( .IN1(n1912), .IN2(n20724), .IN3(n1826), .IN4(n20715), .Q(
        n4920) );
  OA22X1 U28136 ( .IN1(n2084), .IN2(n20763), .IN3(n1998), .IN4(n20745), .Q(
        n4921) );
  NAND4X0 U28137 ( .IN1(n4875), .IN2(n4876), .IN3(n4877), .IN4(n4878), .QN(
        s8_data_o[2]) );
  OA22X1 U28138 ( .IN1(n1739), .IN2(n20698), .IN3(n1634), .IN4(n20683), .Q(
        n4875) );
  OA22X1 U28139 ( .IN1(n1911), .IN2(n4807), .IN3(n1825), .IN4(n20718), .Q(
        n4876) );
  OA22X1 U28140 ( .IN1(n2083), .IN2(n20763), .IN3(n1997), .IN4(n20749), .Q(
        n4877) );
  NAND4X0 U28141 ( .IN1(n4863), .IN2(n4864), .IN3(n4865), .IN4(n4866), .QN(
        s8_data_o[3]) );
  OA22X1 U28142 ( .IN1(n1738), .IN2(n20692), .IN3(n1633), .IN4(n20683), .Q(
        n4863) );
  OA22X1 U28143 ( .IN1(n1910), .IN2(n4807), .IN3(n1824), .IN4(n20718), .Q(
        n4864) );
  OA22X1 U28144 ( .IN1(n2082), .IN2(n20758), .IN3(n1996), .IN4(n20749), .Q(
        n4865) );
  NAND4X0 U28145 ( .IN1(n4859), .IN2(n4860), .IN3(n4861), .IN4(n4862), .QN(
        s8_data_o[4]) );
  OA22X1 U28146 ( .IN1(n1737), .IN2(n20697), .IN3(n1632), .IN4(n20683), .Q(
        n4859) );
  OA22X1 U28147 ( .IN1(n1909), .IN2(n20730), .IN3(n1823), .IN4(n20718), .Q(
        n4860) );
  OA22X1 U28148 ( .IN1(n2081), .IN2(n20762), .IN3(n1995), .IN4(n20749), .Q(
        n4861) );
  NAND4X0 U28149 ( .IN1(n4855), .IN2(n4856), .IN3(n4857), .IN4(n4858), .QN(
        s8_data_o[5]) );
  OA22X1 U28150 ( .IN1(n1736), .IN2(n20698), .IN3(n1631), .IN4(n20683), .Q(
        n4855) );
  OA22X1 U28151 ( .IN1(n1908), .IN2(n20725), .IN3(n1822), .IN4(n20718), .Q(
        n4856) );
  OA22X1 U28152 ( .IN1(n2080), .IN2(n20763), .IN3(n1994), .IN4(n20749), .Q(
        n4857) );
  NAND4X0 U28153 ( .IN1(n4851), .IN2(n4852), .IN3(n4853), .IN4(n4854), .QN(
        s8_data_o[6]) );
  OA22X1 U28154 ( .IN1(n1735), .IN2(n20697), .IN3(n1630), .IN4(n20684), .Q(
        n4851) );
  OA22X1 U28155 ( .IN1(n1907), .IN2(n20730), .IN3(n1821), .IN4(n20716), .Q(
        n4852) );
  OA22X1 U28156 ( .IN1(n2079), .IN2(n20764), .IN3(n1993), .IN4(n20750), .Q(
        n4853) );
  NAND4X0 U28157 ( .IN1(n4847), .IN2(n4848), .IN3(n4849), .IN4(n4850), .QN(
        s8_data_o[7]) );
  OA22X1 U28158 ( .IN1(n1734), .IN2(n20698), .IN3(n1629), .IN4(n20684), .Q(
        n4847) );
  OA22X1 U28159 ( .IN1(n1906), .IN2(n20729), .IN3(n1820), .IN4(n20716), .Q(
        n4848) );
  OA22X1 U28160 ( .IN1(n2078), .IN2(n20764), .IN3(n1992), .IN4(n20750), .Q(
        n4849) );
  NAND4X0 U28161 ( .IN1(n4843), .IN2(n4844), .IN3(n4845), .IN4(n4846), .QN(
        s8_data_o[8]) );
  OA22X1 U28162 ( .IN1(n1733), .IN2(n20695), .IN3(n1628), .IN4(n20684), .Q(
        n4843) );
  OA22X1 U28163 ( .IN1(n1905), .IN2(n20728), .IN3(n1819), .IN4(n20716), .Q(
        n4844) );
  OA22X1 U28164 ( .IN1(n2077), .IN2(n20764), .IN3(n1991), .IN4(n20750), .Q(
        n4845) );
  NAND4X0 U28165 ( .IN1(n4839), .IN2(n4840), .IN3(n4841), .IN4(n4842), .QN(
        s8_data_o[9]) );
  OA22X1 U28166 ( .IN1(n1732), .IN2(n20693), .IN3(n1627), .IN4(n20683), .Q(
        n4839) );
  OA22X1 U28167 ( .IN1(n1904), .IN2(n20726), .IN3(n1818), .IN4(n20716), .Q(
        n4840) );
  OA22X1 U28168 ( .IN1(n2076), .IN2(n20764), .IN3(n1990), .IN4(n20749), .Q(
        n4841) );
  NAND4X0 U28169 ( .IN1(n4959), .IN2(n4960), .IN3(n4961), .IN4(n4962), .QN(
        s8_data_o[10]) );
  OA22X1 U28170 ( .IN1(n1731), .IN2(n20696), .IN3(n1626), .IN4(n20679), .Q(
        n4959) );
  OA22X1 U28171 ( .IN1(n1903), .IN2(n20729), .IN3(n1817), .IN4(n20712), .Q(
        n4960) );
  OA22X1 U28172 ( .IN1(n2075), .IN2(n20763), .IN3(n1989), .IN4(n20738), .Q(
        n4961) );
  NAND4X0 U28173 ( .IN1(n4955), .IN2(n4956), .IN3(n4957), .IN4(n4958), .QN(
        s8_data_o[11]) );
  OA22X1 U28174 ( .IN1(n1730), .IN2(n20696), .IN3(n1625), .IN4(n20679), .Q(
        n4955) );
  OA22X1 U28175 ( .IN1(n1902), .IN2(n20729), .IN3(n1816), .IN4(n20712), .Q(
        n4956) );
  OA22X1 U28176 ( .IN1(n2074), .IN2(n20764), .IN3(n1988), .IN4(n20744), .Q(
        n4957) );
  NAND4X0 U28177 ( .IN1(n4951), .IN2(n4952), .IN3(n4953), .IN4(n4954), .QN(
        s8_data_o[12]) );
  OA22X1 U28178 ( .IN1(n1729), .IN2(n20696), .IN3(n1624), .IN4(n20679), .Q(
        n4951) );
  OA22X1 U28179 ( .IN1(n1901), .IN2(n20729), .IN3(n1815), .IN4(n20712), .Q(
        n4952) );
  OA22X1 U28180 ( .IN1(n2073), .IN2(n20761), .IN3(n1987), .IN4(n20738), .Q(
        n4953) );
  NAND4X0 U28181 ( .IN1(n4947), .IN2(n4948), .IN3(n4949), .IN4(n4950), .QN(
        s8_data_o[13]) );
  OA22X1 U28182 ( .IN1(n1728), .IN2(n20697), .IN3(n1623), .IN4(n20680), .Q(
        n4947) );
  OA22X1 U28183 ( .IN1(n1900), .IN2(n20730), .IN3(n1814), .IN4(n20713), .Q(
        n4948) );
  OA22X1 U28184 ( .IN1(n2072), .IN2(n20762), .IN3(n1986), .IN4(n20745), .Q(
        n4949) );
  NAND4X0 U28185 ( .IN1(n4943), .IN2(n4944), .IN3(n4945), .IN4(n4946), .QN(
        s8_data_o[14]) );
  OA22X1 U28186 ( .IN1(n1727), .IN2(n20697), .IN3(n1622), .IN4(n20680), .Q(
        n4943) );
  OA22X1 U28187 ( .IN1(n1899), .IN2(n20730), .IN3(n1813), .IN4(n20713), .Q(
        n4944) );
  OA22X1 U28188 ( .IN1(n2071), .IN2(n20762), .IN3(n1985), .IN4(n20745), .Q(
        n4945) );
  NAND4X0 U28189 ( .IN1(n4939), .IN2(n4940), .IN3(n4941), .IN4(n4942), .QN(
        s8_data_o[15]) );
  OA22X1 U28190 ( .IN1(n1726), .IN2(n20697), .IN3(n1621), .IN4(n20680), .Q(
        n4939) );
  OA22X1 U28191 ( .IN1(n1898), .IN2(n20730), .IN3(n1812), .IN4(n20713), .Q(
        n4940) );
  OA22X1 U28192 ( .IN1(n2070), .IN2(n20762), .IN3(n1984), .IN4(n20745), .Q(
        n4941) );
  NAND4X0 U28193 ( .IN1(n4935), .IN2(n4936), .IN3(n4937), .IN4(n4938), .QN(
        s8_data_o[16]) );
  OA22X1 U28194 ( .IN1(n1725), .IN2(n20697), .IN3(n1620), .IN4(n20681), .Q(
        n4935) );
  OA22X1 U28195 ( .IN1(n1897), .IN2(n20730), .IN3(n1811), .IN4(n20714), .Q(
        n4936) );
  OA22X1 U28196 ( .IN1(n2069), .IN2(n20762), .IN3(n1983), .IN4(n20746), .Q(
        n4937) );
  NAND4X0 U28197 ( .IN1(n4931), .IN2(n4932), .IN3(n4933), .IN4(n4934), .QN(
        s8_data_o[17]) );
  OA22X1 U28198 ( .IN1(n1724), .IN2(n20698), .IN3(n1619), .IN4(n20681), .Q(
        n4931) );
  OA22X1 U28199 ( .IN1(n1896), .IN2(n20731), .IN3(n1810), .IN4(n20714), .Q(
        n4932) );
  OA22X1 U28200 ( .IN1(n2068), .IN2(n20763), .IN3(n1982), .IN4(n20746), .Q(
        n4933) );
  NAND4X0 U28201 ( .IN1(n4927), .IN2(n4928), .IN3(n4929), .IN4(n4930), .QN(
        s8_data_o[18]) );
  OA22X1 U28202 ( .IN1(n1723), .IN2(n20698), .IN3(n1618), .IN4(n20681), .Q(
        n4927) );
  OA22X1 U28203 ( .IN1(n1895), .IN2(n4807), .IN3(n1809), .IN4(n20714), .Q(
        n4928) );
  OA22X1 U28204 ( .IN1(n2067), .IN2(n20763), .IN3(n1981), .IN4(n20746), .Q(
        n4929) );
  NAND4X0 U28205 ( .IN1(n4923), .IN2(n4924), .IN3(n4925), .IN4(n4926), .QN(
        s8_data_o[19]) );
  OA22X1 U28206 ( .IN1(n1722), .IN2(n20698), .IN3(n1617), .IN4(n20681), .Q(
        n4923) );
  OA22X1 U28207 ( .IN1(n1894), .IN2(n4807), .IN3(n1808), .IN4(n20715), .Q(
        n4924) );
  OA22X1 U28208 ( .IN1(n2066), .IN2(n20763), .IN3(n1980), .IN4(n20746), .Q(
        n4925) );
  NAND4X0 U28209 ( .IN1(n4915), .IN2(n4916), .IN3(n4917), .IN4(n4918), .QN(
        s8_data_o[20]) );
  OA22X1 U28210 ( .IN1(n1721), .IN2(n20696), .IN3(n1616), .IN4(n20680), .Q(
        n4915) );
  OA22X1 U28211 ( .IN1(n1893), .IN2(n20729), .IN3(n1807), .IN4(n20715), .Q(
        n4916) );
  OA22X1 U28212 ( .IN1(n2065), .IN2(n20759), .IN3(n1979), .IN4(n20749), .Q(
        n4917) );
  NAND4X0 U28213 ( .IN1(n4911), .IN2(n4912), .IN3(n4913), .IN4(n4914), .QN(
        s8_data_o[21]) );
  OA22X1 U28214 ( .IN1(n1720), .IN2(n20697), .IN3(n1615), .IN4(n20683), .Q(
        n4911) );
  OA22X1 U28215 ( .IN1(n1892), .IN2(n4807), .IN3(n1806), .IN4(n20716), .Q(
        n4912) );
  OA22X1 U28216 ( .IN1(n2064), .IN2(n20762), .IN3(n1978), .IN4(n20747), .Q(
        n4913) );
  NAND4X0 U28217 ( .IN1(n4907), .IN2(n4908), .IN3(n4909), .IN4(n4910), .QN(
        s8_data_o[22]) );
  OA22X1 U28218 ( .IN1(n1719), .IN2(n20697), .IN3(n1614), .IN4(n20667), .Q(
        n4907) );
  OA22X1 U28219 ( .IN1(n1891), .IN2(n20730), .IN3(n1805), .IN4(n20716), .Q(
        n4908) );
  OA22X1 U28220 ( .IN1(n2063), .IN2(n20762), .IN3(n1977), .IN4(n20747), .Q(
        n4909) );
  NAND4X0 U28221 ( .IN1(n4903), .IN2(n4904), .IN3(n4905), .IN4(n4906), .QN(
        s8_data_o[23]) );
  OA22X1 U28222 ( .IN1(n1718), .IN2(n20698), .IN3(n1613), .IN4(n20685), .Q(
        n4903) );
  OA22X1 U28223 ( .IN1(n1890), .IN2(n20730), .IN3(n1804), .IN4(n20716), .Q(
        n4904) );
  OA22X1 U28224 ( .IN1(n2062), .IN2(n20763), .IN3(n1976), .IN4(n20747), .Q(
        n4905) );
  NAND4X0 U28225 ( .IN1(n4899), .IN2(n4900), .IN3(n4901), .IN4(n4902), .QN(
        s8_data_o[24]) );
  OA22X1 U28226 ( .IN1(n1717), .IN2(n20696), .IN3(n1612), .IN4(n20682), .Q(
        n4899) );
  OA22X1 U28227 ( .IN1(n1889), .IN2(n20731), .IN3(n1803), .IN4(n20717), .Q(
        n4900) );
  OA22X1 U28228 ( .IN1(n2061), .IN2(n20764), .IN3(n1975), .IN4(n20748), .Q(
        n4901) );
  NAND4X0 U28229 ( .IN1(n4895), .IN2(n4896), .IN3(n4897), .IN4(n4898), .QN(
        s8_data_o[25]) );
  OA22X1 U28230 ( .IN1(n1716), .IN2(n20695), .IN3(n1611), .IN4(n20682), .Q(
        n4895) );
  OA22X1 U28231 ( .IN1(n1888), .IN2(n20728), .IN3(n1802), .IN4(n20717), .Q(
        n4896) );
  OA22X1 U28232 ( .IN1(n2060), .IN2(n20761), .IN3(n1974), .IN4(n20748), .Q(
        n4897) );
  NAND4X0 U28233 ( .IN1(n4891), .IN2(n4892), .IN3(n4893), .IN4(n4894), .QN(
        s8_data_o[26]) );
  OA22X1 U28234 ( .IN1(n1715), .IN2(n20693), .IN3(n1610), .IN4(n20682), .Q(
        n4891) );
  OA22X1 U28235 ( .IN1(n1887), .IN2(n20726), .IN3(n1801), .IN4(n20717), .Q(
        n4892) );
  OA22X1 U28236 ( .IN1(n2059), .IN2(n20759), .IN3(n1973), .IN4(n20748), .Q(
        n4893) );
  NAND4X0 U28237 ( .IN1(n4887), .IN2(n4888), .IN3(n4889), .IN4(n4890), .QN(
        s8_data_o[27]) );
  OA22X1 U28238 ( .IN1(n1714), .IN2(n20696), .IN3(n1609), .IN4(n20685), .Q(
        n4887) );
  OA22X1 U28239 ( .IN1(n1886), .IN2(n20729), .IN3(n1800), .IN4(n20716), .Q(
        n4888) );
  OA22X1 U28240 ( .IN1(n2058), .IN2(n20759), .IN3(n1972), .IN4(n20747), .Q(
        n4889) );
  NAND4X0 U28241 ( .IN1(n4883), .IN2(n4884), .IN3(n4885), .IN4(n4886), .QN(
        s8_data_o[28]) );
  OA22X1 U28242 ( .IN1(n1713), .IN2(n20691), .IN3(n1608), .IN4(n20682), .Q(
        n4883) );
  OA22X1 U28243 ( .IN1(n1885), .IN2(n4807), .IN3(n1799), .IN4(n20717), .Q(
        n4884) );
  OA22X1 U28244 ( .IN1(n2057), .IN2(n20757), .IN3(n1971), .IN4(n20748), .Q(
        n4885) );
  NAND4X0 U28245 ( .IN1(n4879), .IN2(n4880), .IN3(n4881), .IN4(n4882), .QN(
        s8_data_o[29]) );
  OA22X1 U28246 ( .IN1(n1712), .IN2(n20694), .IN3(n1607), .IN4(n20684), .Q(
        n4879) );
  OA22X1 U28247 ( .IN1(n1884), .IN2(n4807), .IN3(n1798), .IN4(n20716), .Q(
        n4880) );
  OA22X1 U28248 ( .IN1(n2056), .IN2(n4805), .IN3(n1970), .IN4(n20747), .Q(
        n4881) );
  NAND4X0 U28249 ( .IN1(n4871), .IN2(n4872), .IN3(n4873), .IN4(n4874), .QN(
        s8_data_o[30]) );
  OA22X1 U28250 ( .IN1(n1711), .IN2(n20695), .IN3(n1606), .IN4(n20683), .Q(
        n4871) );
  OA22X1 U28251 ( .IN1(n1883), .IN2(n4807), .IN3(n1797), .IN4(n20718), .Q(
        n4872) );
  OA22X1 U28252 ( .IN1(n2055), .IN2(n4805), .IN3(n1969), .IN4(n20749), .Q(
        n4873) );
  NAND4X0 U28253 ( .IN1(n4867), .IN2(n4868), .IN3(n4869), .IN4(n4870), .QN(
        s8_data_o[31]) );
  OA22X1 U28254 ( .IN1(n1710), .IN2(n20696), .IN3(n1605), .IN4(n20683), .Q(
        n4867) );
  OA22X1 U28255 ( .IN1(n1882), .IN2(n20729), .IN3(n1796), .IN4(n20718), .Q(
        n4868) );
  OA22X1 U28256 ( .IN1(n2054), .IN2(n20759), .IN3(n1968), .IN4(n20749), .Q(
        n4869) );
  NAND4X0 U28257 ( .IN1(n5107), .IN2(n5108), .IN3(n5109), .IN4(n5110), .QN(
        s7_stb_o) );
  OA22X1 U28258 ( .IN1(n1795), .IN2(n5117), .IN3(n1709), .IN4(n5118), .Q(n5107) );
  OA22X1 U28259 ( .IN1(n1967), .IN2(n5115), .IN3(n1881), .IN4(n5116), .Q(n5108) );
  OA22X1 U28260 ( .IN1(n2139), .IN2(n5113), .IN3(n2053), .IN4(n5114), .Q(n5109) );
  NAND4X0 U28261 ( .IN1(n5095), .IN2(n5096), .IN3(n5097), .IN4(n5098), .QN(
        s7_we_o) );
  OA22X1 U28262 ( .IN1(n1794), .IN2(n20566), .IN3(n1708), .IN4(n20553), .Q(
        n5095) );
  OA22X1 U28263 ( .IN1(n1966), .IN2(n20592), .IN3(n1880), .IN4(n20586), .Q(
        n5096) );
  OA22X1 U28264 ( .IN1(n2138), .IN2(n20625), .IN3(n2052), .IN4(n20620), .Q(
        n5097) );
  NAND4X0 U28265 ( .IN1(n5131), .IN2(n5132), .IN3(n5133), .IN4(n5134), .QN(
        s7_sel_o[0]) );
  OA22X1 U28266 ( .IN1(n1793), .IN2(n20566), .IN3(n1707), .IN4(n20552), .Q(
        n5131) );
  OA22X1 U28267 ( .IN1(n1965), .IN2(n20599), .IN3(n1879), .IN4(n20585), .Q(
        n5132) );
  OA22X1 U28268 ( .IN1(n2137), .IN2(n20629), .IN3(n2051), .IN4(n20619), .Q(
        n5133) );
  NAND4X0 U28269 ( .IN1(n5127), .IN2(n5128), .IN3(n5129), .IN4(n5130), .QN(
        s7_sel_o[1]) );
  OA22X1 U28270 ( .IN1(n1792), .IN2(n20566), .IN3(n1706), .IN4(n20552), .Q(
        n5127) );
  OA22X1 U28271 ( .IN1(n1964), .IN2(n20599), .IN3(n1878), .IN4(n20585), .Q(
        n5128) );
  OA22X1 U28272 ( .IN1(n2136), .IN2(n20630), .IN3(n2050), .IN4(n20619), .Q(
        n5129) );
  NAND4X0 U28273 ( .IN1(n5123), .IN2(n5124), .IN3(n5125), .IN4(n5126), .QN(
        s7_sel_o[2]) );
  OA22X1 U28274 ( .IN1(n1791), .IN2(n20566), .IN3(n1705), .IN4(n20553), .Q(
        n5123) );
  OA22X1 U28275 ( .IN1(n1963), .IN2(n20599), .IN3(n1877), .IN4(n20586), .Q(
        n5124) );
  OA22X1 U28276 ( .IN1(n2135), .IN2(n20631), .IN3(n2049), .IN4(n20620), .Q(
        n5125) );
  NAND4X0 U28277 ( .IN1(n5119), .IN2(n5120), .IN3(n5121), .IN4(n5122), .QN(
        s7_sel_o[3]) );
  OA22X1 U28278 ( .IN1(n1790), .IN2(n20566), .IN3(n1704), .IN4(n20553), .Q(
        n5119) );
  OA22X1 U28279 ( .IN1(n1962), .IN2(n20599), .IN3(n1876), .IN4(n20586), .Q(
        n5120) );
  OA22X1 U28280 ( .IN1(n2134), .IN2(n20625), .IN3(n2048), .IN4(n20620), .Q(
        n5121) );
  NAND4X0 U28281 ( .IN1(n5387), .IN2(n5388), .IN3(n5389), .IN4(n5390), .QN(
        s7_addr_o[0]) );
  OA22X1 U28282 ( .IN1(n1789), .IN2(n20561), .IN3(n1703), .IN4(n20536), .Q(
        n5387) );
  OA22X1 U28283 ( .IN1(n1961), .IN2(n20592), .IN3(n1875), .IN4(n20569), .Q(
        n5388) );
  OA22X1 U28284 ( .IN1(n2133), .IN2(n20625), .IN3(n2047), .IN4(n20602), .Q(
        n5389) );
  NAND4X0 U28285 ( .IN1(n5343), .IN2(n5344), .IN3(n5345), .IN4(n5346), .QN(
        s7_addr_o[1]) );
  OA22X1 U28286 ( .IN1(n1788), .IN2(n20560), .IN3(n1702), .IN4(n20539), .Q(
        n5343) );
  OA22X1 U28287 ( .IN1(n1960), .IN2(n20594), .IN3(n1874), .IN4(n20572), .Q(
        n5344) );
  OA22X1 U28288 ( .IN1(n2132), .IN2(n20627), .IN3(n2046), .IN4(n20605), .Q(
        n5345) );
  NAND4X0 U28289 ( .IN1(n5299), .IN2(n5300), .IN3(n5301), .IN4(n5302), .QN(
        s7_addr_o[2]) );
  OA22X1 U28290 ( .IN1(n1787), .IN2(n20560), .IN3(n1701), .IN4(n20543), .Q(
        n5299) );
  OA22X1 U28291 ( .IN1(n1959), .IN2(n20594), .IN3(n1873), .IN4(n20576), .Q(
        n5300) );
  OA22X1 U28292 ( .IN1(n2131), .IN2(n20625), .IN3(n2045), .IN4(n20609), .Q(
        n5301) );
  NAND4X0 U28293 ( .IN1(n5287), .IN2(n5288), .IN3(n5289), .IN4(n5290), .QN(
        s7_addr_o[3]) );
  OA22X1 U28294 ( .IN1(n1786), .IN2(n20566), .IN3(n1699), .IN4(n20544), .Q(
        n5287) );
  OA22X1 U28295 ( .IN1(n1958), .IN2(n20599), .IN3(n1872), .IN4(n20577), .Q(
        n5288) );
  OA22X1 U28296 ( .IN1(n2130), .IN2(n20626), .IN3(n2044), .IN4(n20610), .Q(
        n5289) );
  NAND4X0 U28297 ( .IN1(n5283), .IN2(n5284), .IN3(n5285), .IN4(n5286), .QN(
        s7_addr_o[4]) );
  OA22X1 U28298 ( .IN1(n1785), .IN2(n20561), .IN3(n1697), .IN4(n20544), .Q(
        n5283) );
  OA22X1 U28299 ( .IN1(n1957), .IN2(n20592), .IN3(n1871), .IN4(n20577), .Q(
        n5284) );
  OA22X1 U28300 ( .IN1(n2129), .IN2(n20628), .IN3(n2043), .IN4(n20610), .Q(
        n5285) );
  NAND4X0 U28301 ( .IN1(n5279), .IN2(n5280), .IN3(n5281), .IN4(n5282), .QN(
        s7_addr_o[5]) );
  OA22X1 U28302 ( .IN1(n1784), .IN2(n20566), .IN3(n1696), .IN4(n20544), .Q(
        n5279) );
  OA22X1 U28303 ( .IN1(n1956), .IN2(n20599), .IN3(n1870), .IN4(n20576), .Q(
        n5280) );
  OA22X1 U28304 ( .IN1(n2128), .IN2(n20632), .IN3(n2042), .IN4(n20611), .Q(
        n5281) );
  NAND4X0 U28305 ( .IN1(n5275), .IN2(n5276), .IN3(n5277), .IN4(n5278), .QN(
        s7_addr_o[6]) );
  OA22X1 U28306 ( .IN1(n1783), .IN2(n20562), .IN3(n1679), .IN4(n20544), .Q(
        n5275) );
  OA22X1 U28307 ( .IN1(n1955), .IN2(n20595), .IN3(n1869), .IN4(n20577), .Q(
        n5276) );
  OA22X1 U28308 ( .IN1(n2127), .IN2(n20628), .IN3(n2041), .IN4(n20611), .Q(
        n5277) );
  NAND4X0 U28309 ( .IN1(n5271), .IN2(n5272), .IN3(n5273), .IN4(n5274), .QN(
        s7_addr_o[7]) );
  OA22X1 U28310 ( .IN1(n1782), .IN2(n20562), .IN3(n1678), .IN4(n20544), .Q(
        n5271) );
  OA22X1 U28311 ( .IN1(n1954), .IN2(n20595), .IN3(n1868), .IN4(n20569), .Q(
        n5272) );
  OA22X1 U28312 ( .IN1(n2126), .IN2(n20628), .IN3(n2040), .IN4(n20611), .Q(
        n5273) );
  NAND4X0 U28313 ( .IN1(n5267), .IN2(n5268), .IN3(n5269), .IN4(n5270), .QN(
        s7_addr_o[8]) );
  OA22X1 U28314 ( .IN1(n1781), .IN2(n20562), .IN3(n1677), .IN4(n20545), .Q(
        n5267) );
  OA22X1 U28315 ( .IN1(n1953), .IN2(n20595), .IN3(n1867), .IN4(n20578), .Q(
        n5268) );
  OA22X1 U28316 ( .IN1(n2125), .IN2(n20628), .IN3(n2039), .IN4(n20612), .Q(
        n5269) );
  NAND4X0 U28317 ( .IN1(n5263), .IN2(n5264), .IN3(n5265), .IN4(n5266), .QN(
        s7_addr_o[9]) );
  OA22X1 U28318 ( .IN1(n1780), .IN2(n20562), .IN3(n1676), .IN4(n20545), .Q(
        n5263) );
  OA22X1 U28319 ( .IN1(n1952), .IN2(n20595), .IN3(n1866), .IN4(n20578), .Q(
        n5264) );
  OA22X1 U28320 ( .IN1(n2124), .IN2(n20628), .IN3(n2038), .IN4(n20612), .Q(
        n5265) );
  NAND4X0 U28321 ( .IN1(n5383), .IN2(n5384), .IN3(n5385), .IN4(n5386), .QN(
        s7_addr_o[10]) );
  OA22X1 U28322 ( .IN1(n1779), .IN2(n20562), .IN3(n1675), .IN4(n20536), .Q(
        n5383) );
  OA22X1 U28323 ( .IN1(n1951), .IN2(n20592), .IN3(n1865), .IN4(n20569), .Q(
        n5384) );
  OA22X1 U28324 ( .IN1(n2123), .IN2(n20625), .IN3(n2037), .IN4(n20602), .Q(
        n5385) );
  NAND4X0 U28325 ( .IN1(n5379), .IN2(n5380), .IN3(n5381), .IN4(n5382), .QN(
        s7_addr_o[11]) );
  OA22X1 U28326 ( .IN1(n1778), .IN2(n20560), .IN3(n1674), .IN4(n20536), .Q(
        n5379) );
  OA22X1 U28327 ( .IN1(n1950), .IN2(n20592), .IN3(n1864), .IN4(n20569), .Q(
        n5380) );
  OA22X1 U28328 ( .IN1(n2122), .IN2(n20625), .IN3(n2036), .IN4(n20602), .Q(
        n5381) );
  NAND4X0 U28329 ( .IN1(n5375), .IN2(n5376), .IN3(n5377), .IN4(n5378), .QN(
        s7_addr_o[12]) );
  OA22X1 U28330 ( .IN1(n1777), .IN2(n20559), .IN3(n1673), .IN4(n20537), .Q(
        n5375) );
  OA22X1 U28331 ( .IN1(n1949), .IN2(n20592), .IN3(n1863), .IN4(n20570), .Q(
        n5376) );
  OA22X1 U28332 ( .IN1(n2121), .IN2(n20625), .IN3(n2035), .IN4(n20603), .Q(
        n5377) );
  NAND4X0 U28333 ( .IN1(n5371), .IN2(n5372), .IN3(n5373), .IN4(n5374), .QN(
        s7_addr_o[13]) );
  OA22X1 U28334 ( .IN1(n1776), .IN2(n20559), .IN3(n1672), .IN4(n20537), .Q(
        n5371) );
  OA22X1 U28335 ( .IN1(n1948), .IN2(n20593), .IN3(n1862), .IN4(n20570), .Q(
        n5372) );
  OA22X1 U28336 ( .IN1(n2120), .IN2(n20626), .IN3(n2034), .IN4(n20603), .Q(
        n5373) );
  NAND4X0 U28337 ( .IN1(n5367), .IN2(n5368), .IN3(n5369), .IN4(n5370), .QN(
        s7_addr_o[14]) );
  OA22X1 U28338 ( .IN1(n1775), .IN2(n20559), .IN3(n1671), .IN4(n20537), .Q(
        n5367) );
  OA22X1 U28339 ( .IN1(n1947), .IN2(n20593), .IN3(n1861), .IN4(n20570), .Q(
        n5368) );
  OA22X1 U28340 ( .IN1(n2119), .IN2(n20626), .IN3(n2033), .IN4(n20603), .Q(
        n5369) );
  NAND4X0 U28341 ( .IN1(n5363), .IN2(n5364), .IN3(n5365), .IN4(n5366), .QN(
        s7_addr_o[15]) );
  OA22X1 U28342 ( .IN1(n1774), .IN2(n20559), .IN3(n1670), .IN4(n20538), .Q(
        n5363) );
  OA22X1 U28343 ( .IN1(n1946), .IN2(n20593), .IN3(n1860), .IN4(n20571), .Q(
        n5364) );
  OA22X1 U28344 ( .IN1(n2118), .IN2(n20626), .IN3(n2032), .IN4(n20604), .Q(
        n5365) );
  NAND4X0 U28345 ( .IN1(n5359), .IN2(n5360), .IN3(n5361), .IN4(n5362), .QN(
        s7_addr_o[16]) );
  OA22X1 U28346 ( .IN1(n1773), .IN2(n20559), .IN3(n1669), .IN4(n20538), .Q(
        n5359) );
  OA22X1 U28347 ( .IN1(n1945), .IN2(n20593), .IN3(n1859), .IN4(n20571), .Q(
        n5360) );
  OA22X1 U28348 ( .IN1(n2117), .IN2(n20626), .IN3(n2031), .IN4(n20604), .Q(
        n5361) );
  NAND4X0 U28349 ( .IN1(n5355), .IN2(n5356), .IN3(n5357), .IN4(n5358), .QN(
        s7_addr_o[17]) );
  OA22X1 U28350 ( .IN1(n1772), .IN2(n20560), .IN3(n1668), .IN4(n20538), .Q(
        n5355) );
  OA22X1 U28351 ( .IN1(n1944), .IN2(n20594), .IN3(n1858), .IN4(n20571), .Q(
        n5356) );
  OA22X1 U28352 ( .IN1(n2116), .IN2(n20627), .IN3(n2030), .IN4(n20604), .Q(
        n5357) );
  NAND4X0 U28353 ( .IN1(n5351), .IN2(n5352), .IN3(n5353), .IN4(n5354), .QN(
        s7_addr_o[18]) );
  OA22X1 U28354 ( .IN1(n1771), .IN2(n20560), .IN3(n1667), .IN4(n20539), .Q(
        n5351) );
  OA22X1 U28355 ( .IN1(n1943), .IN2(n20594), .IN3(n1857), .IN4(n20572), .Q(
        n5352) );
  OA22X1 U28356 ( .IN1(n2115), .IN2(n20627), .IN3(n2029), .IN4(n20605), .Q(
        n5353) );
  NAND4X0 U28357 ( .IN1(n5347), .IN2(n5348), .IN3(n5349), .IN4(n5350), .QN(
        s7_addr_o[19]) );
  OA22X1 U28358 ( .IN1(n1770), .IN2(n20560), .IN3(n1666), .IN4(n20539), .Q(
        n5347) );
  OA22X1 U28359 ( .IN1(n1942), .IN2(n20594), .IN3(n1856), .IN4(n20572), .Q(
        n5348) );
  OA22X1 U28360 ( .IN1(n2114), .IN2(n20627), .IN3(n2028), .IN4(n20605), .Q(
        n5349) );
  NAND4X0 U28361 ( .IN1(n5339), .IN2(n5340), .IN3(n5341), .IN4(n5342), .QN(
        s7_addr_o[20]) );
  OA22X1 U28362 ( .IN1(n1769), .IN2(n20559), .IN3(n1665), .IN4(n20540), .Q(
        n5339) );
  OA22X1 U28363 ( .IN1(n1941), .IN2(n20593), .IN3(n1855), .IN4(n20573), .Q(
        n5340) );
  OA22X1 U28364 ( .IN1(n2113), .IN2(n20626), .IN3(n2027), .IN4(n20606), .Q(
        n5341) );
  NAND4X0 U28365 ( .IN1(n5335), .IN2(n5336), .IN3(n5337), .IN4(n5338), .QN(
        s7_addr_o[21]) );
  OA22X1 U28366 ( .IN1(n1768), .IN2(n20559), .IN3(n1664), .IN4(n20540), .Q(
        n5335) );
  OA22X1 U28367 ( .IN1(n1940), .IN2(n20593), .IN3(n1854), .IN4(n20573), .Q(
        n5336) );
  OA22X1 U28368 ( .IN1(n2112), .IN2(n20626), .IN3(n2026), .IN4(n20606), .Q(
        n5337) );
  NAND4X0 U28369 ( .IN1(n5331), .IN2(n5332), .IN3(n5333), .IN4(n5334), .QN(
        s7_addr_o[22]) );
  OA22X1 U28370 ( .IN1(n1767), .IN2(n20561), .IN3(n1663), .IN4(n20540), .Q(
        n5331) );
  OA22X1 U28371 ( .IN1(n1939), .IN2(n20592), .IN3(n1853), .IN4(n20573), .Q(
        n5332) );
  OA22X1 U28372 ( .IN1(n2111), .IN2(n20625), .IN3(n2025), .IN4(n20606), .Q(
        n5333) );
  NAND4X0 U28373 ( .IN1(n5327), .IN2(n5328), .IN3(n5329), .IN4(n5330), .QN(
        s7_addr_o[23]) );
  OA22X1 U28374 ( .IN1(n1766), .IN2(n20559), .IN3(n1662), .IN4(n20541), .Q(
        n5327) );
  OA22X1 U28375 ( .IN1(n1938), .IN2(n20593), .IN3(n1852), .IN4(n20574), .Q(
        n5328) );
  OA22X1 U28376 ( .IN1(n2110), .IN2(n20626), .IN3(n2024), .IN4(n20607), .Q(
        n5329) );
  NAND4X0 U28377 ( .IN1(n5323), .IN2(n5324), .IN3(n5325), .IN4(n5326), .QN(
        s7_addr_o[24]) );
  OA22X1 U28378 ( .IN1(n1765), .IN2(n20561), .IN3(n1661), .IN4(n20541), .Q(
        n5323) );
  OA22X1 U28379 ( .IN1(n1937), .IN2(n20599), .IN3(n1851), .IN4(n20574), .Q(
        n5324) );
  OA22X1 U28380 ( .IN1(n2109), .IN2(n20627), .IN3(n2023), .IN4(n20607), .Q(
        n5325) );
  NAND4X0 U28381 ( .IN1(n5319), .IN2(n5320), .IN3(n5321), .IN4(n5322), .QN(
        s7_addr_o[25]) );
  OA22X1 U28382 ( .IN1(n1764), .IN2(n20561), .IN3(n1660), .IN4(n20541), .Q(
        n5319) );
  OA22X1 U28383 ( .IN1(n1936), .IN2(n20595), .IN3(n1850), .IN4(n20574), .Q(
        n5320) );
  OA22X1 U28384 ( .IN1(n2108), .IN2(n20626), .IN3(n2022), .IN4(n20607), .Q(
        n5321) );
  NAND4X0 U28385 ( .IN1(n5315), .IN2(n5316), .IN3(n5317), .IN4(n5318), .QN(
        s7_addr_o[26]) );
  OA22X1 U28386 ( .IN1(n1763), .IN2(n20561), .IN3(n1659), .IN4(n20542), .Q(
        n5315) );
  OA22X1 U28387 ( .IN1(n1935), .IN2(n20594), .IN3(n1849), .IN4(n20575), .Q(
        n5316) );
  OA22X1 U28388 ( .IN1(n2107), .IN2(n20632), .IN3(n2021), .IN4(n20608), .Q(
        n5317) );
  NAND4X0 U28389 ( .IN1(n5311), .IN2(n5312), .IN3(n5313), .IN4(n5314), .QN(
        s7_addr_o[27]) );
  OA22X1 U28390 ( .IN1(n1762), .IN2(n20561), .IN3(n1658), .IN4(n20542), .Q(
        n5311) );
  OA22X1 U28391 ( .IN1(n1934), .IN2(n20593), .IN3(n1848), .IN4(n20575), .Q(
        n5312) );
  OA22X1 U28392 ( .IN1(n2106), .IN2(n20629), .IN3(n2020), .IN4(n20608), .Q(
        n5313) );
  NAND4X0 U28393 ( .IN1(n5307), .IN2(n5308), .IN3(n5309), .IN4(n5310), .QN(
        s7_addr_o[28]) );
  OA22X1 U28394 ( .IN1(n1761), .IN2(n20559), .IN3(n1657), .IN4(n20542), .Q(
        n5307) );
  OA22X1 U28395 ( .IN1(n1933), .IN2(n20593), .IN3(n1847), .IN4(n20575), .Q(
        n5308) );
  OA22X1 U28396 ( .IN1(n2105), .IN2(n20628), .IN3(n2019), .IN4(n20608), .Q(
        n5309) );
  NAND4X0 U28397 ( .IN1(n5303), .IN2(n5304), .IN3(n5305), .IN4(n5306), .QN(
        s7_addr_o[29]) );
  OA22X1 U28398 ( .IN1(n1760), .IN2(n20565), .IN3(n1656), .IN4(n20543), .Q(
        n5303) );
  OA22X1 U28399 ( .IN1(n1932), .IN2(n20597), .IN3(n1846), .IN4(n20576), .Q(
        n5304) );
  OA22X1 U28400 ( .IN1(n2104), .IN2(n20627), .IN3(n2018), .IN4(n20609), .Q(
        n5305) );
  NAND4X0 U28401 ( .IN1(n5295), .IN2(n5296), .IN3(n5297), .IN4(n5298), .QN(
        s7_addr_o[30]) );
  OA22X1 U28402 ( .IN1(n1759), .IN2(n20564), .IN3(n1655), .IN4(n20543), .Q(
        n5295) );
  OA22X1 U28403 ( .IN1(n1931), .IN2(n20598), .IN3(n1845), .IN4(n20576), .Q(
        n5296) );
  OA22X1 U28404 ( .IN1(n2103), .IN2(n20627), .IN3(n2017), .IN4(n20609), .Q(
        n5297) );
  NAND4X0 U28405 ( .IN1(n5291), .IN2(n5292), .IN3(n5293), .IN4(n5294), .QN(
        s7_addr_o[31]) );
  OA22X1 U28406 ( .IN1(n1758), .IN2(n20563), .IN3(n1650), .IN4(n20543), .Q(
        n5291) );
  OA22X1 U28407 ( .IN1(n1930), .IN2(n20596), .IN3(n1844), .IN4(n20577), .Q(
        n5292) );
  OA22X1 U28408 ( .IN1(n2102), .IN2(n20628), .IN3(n2016), .IN4(n20610), .Q(
        n5293) );
  NAND4X0 U28409 ( .IN1(n5259), .IN2(n5260), .IN3(n5261), .IN4(n5262), .QN(
        s7_data_o[0]) );
  OA22X1 U28410 ( .IN1(n1741), .IN2(n20562), .IN3(n1636), .IN4(n20545), .Q(
        n5259) );
  OA22X1 U28411 ( .IN1(n1913), .IN2(n20595), .IN3(n1827), .IN4(n20578), .Q(
        n5260) );
  OA22X1 U28412 ( .IN1(n2085), .IN2(n20629), .IN3(n1999), .IN4(n20612), .Q(
        n5261) );
  NAND4X0 U28413 ( .IN1(n5215), .IN2(n5216), .IN3(n5217), .IN4(n5218), .QN(
        s7_data_o[1]) );
  OA22X1 U28414 ( .IN1(n1740), .IN2(n20560), .IN3(n1635), .IN4(n20547), .Q(
        n5215) );
  OA22X1 U28415 ( .IN1(n1912), .IN2(n20597), .IN3(n1826), .IN4(n20576), .Q(
        n5216) );
  OA22X1 U28416 ( .IN1(n2084), .IN2(n20630), .IN3(n1998), .IN4(n20613), .Q(
        n5217) );
  NAND4X0 U28417 ( .IN1(n5171), .IN2(n5172), .IN3(n5173), .IN4(n5174), .QN(
        s7_data_o[2]) );
  OA22X1 U28418 ( .IN1(n1739), .IN2(n20564), .IN3(n1634), .IN4(n20551), .Q(
        n5171) );
  OA22X1 U28419 ( .IN1(n1911), .IN2(n20598), .IN3(n1825), .IN4(n20569), .Q(
        n5172) );
  OA22X1 U28420 ( .IN1(n2083), .IN2(n20632), .IN3(n1997), .IN4(n20601), .Q(
        n5173) );
  NAND4X0 U28421 ( .IN1(n5159), .IN2(n5160), .IN3(n5161), .IN4(n5162), .QN(
        s7_data_o[3]) );
  OA22X1 U28422 ( .IN1(n1738), .IN2(n20563), .IN3(n1633), .IN4(n20551), .Q(
        n5159) );
  OA22X1 U28423 ( .IN1(n1910), .IN2(n20596), .IN3(n1824), .IN4(n20571), .Q(
        n5160) );
  OA22X1 U28424 ( .IN1(n2082), .IN2(n20632), .IN3(n1996), .IN4(n20615), .Q(
        n5161) );
  NAND4X0 U28425 ( .IN1(n5155), .IN2(n5156), .IN3(n5157), .IN4(n5158), .QN(
        s7_data_o[4]) );
  OA22X1 U28426 ( .IN1(n1737), .IN2(n20565), .IN3(n1632), .IN4(n20551), .Q(
        n5155) );
  OA22X1 U28427 ( .IN1(n1909), .IN2(n20597), .IN3(n1823), .IN4(n20586), .Q(
        n5156) );
  OA22X1 U28428 ( .IN1(n2081), .IN2(n20629), .IN3(n1995), .IN4(n20616), .Q(
        n5157) );
  NAND4X0 U28429 ( .IN1(n5151), .IN2(n5152), .IN3(n5153), .IN4(n5154), .QN(
        s7_data_o[5]) );
  OA22X1 U28430 ( .IN1(n1736), .IN2(n20564), .IN3(n1631), .IN4(n20551), .Q(
        n5151) );
  OA22X1 U28431 ( .IN1(n1908), .IN2(n20598), .IN3(n1822), .IN4(n20584), .Q(
        n5152) );
  OA22X1 U28432 ( .IN1(n2080), .IN2(n20630), .IN3(n1994), .IN4(n20617), .Q(
        n5153) );
  NAND4X0 U28433 ( .IN1(n5147), .IN2(n5148), .IN3(n5149), .IN4(n5150), .QN(
        s7_data_o[6]) );
  OA22X1 U28434 ( .IN1(n1735), .IN2(n20565), .IN3(n1630), .IN4(n20553), .Q(
        n5147) );
  OA22X1 U28435 ( .IN1(n1907), .IN2(n20594), .IN3(n1821), .IN4(n20584), .Q(
        n5148) );
  OA22X1 U28436 ( .IN1(n2079), .IN2(n20630), .IN3(n1993), .IN4(n20618), .Q(
        n5149) );
  NAND4X0 U28437 ( .IN1(n5143), .IN2(n5144), .IN3(n5145), .IN4(n5146), .QN(
        s7_data_o[7]) );
  OA22X1 U28438 ( .IN1(n1734), .IN2(n20565), .IN3(n1629), .IN4(n20553), .Q(
        n5143) );
  OA22X1 U28439 ( .IN1(n1906), .IN2(n20592), .IN3(n1820), .IN4(n20584), .Q(
        n5144) );
  OA22X1 U28440 ( .IN1(n2078), .IN2(n20631), .IN3(n1992), .IN4(n20618), .Q(
        n5145) );
  NAND4X0 U28441 ( .IN1(n5139), .IN2(n5140), .IN3(n5141), .IN4(n5142), .QN(
        s7_data_o[8]) );
  OA22X1 U28442 ( .IN1(n1733), .IN2(n20565), .IN3(n1628), .IN4(n20553), .Q(
        n5139) );
  OA22X1 U28443 ( .IN1(n1905), .IN2(n20599), .IN3(n1819), .IN4(n20584), .Q(
        n5140) );
  OA22X1 U28444 ( .IN1(n2077), .IN2(n20628), .IN3(n1991), .IN4(n20618), .Q(
        n5141) );
  NAND4X0 U28445 ( .IN1(n5135), .IN2(n5136), .IN3(n5137), .IN4(n5138), .QN(
        s7_data_o[9]) );
  OA22X1 U28446 ( .IN1(n1732), .IN2(n20565), .IN3(n1627), .IN4(n20552), .Q(
        n5135) );
  OA22X1 U28447 ( .IN1(n1904), .IN2(n20592), .IN3(n1818), .IN4(n20585), .Q(
        n5136) );
  OA22X1 U28448 ( .IN1(n2076), .IN2(n20627), .IN3(n1990), .IN4(n20619), .Q(
        n5137) );
  NAND4X0 U28449 ( .IN1(n5255), .IN2(n5256), .IN3(n5257), .IN4(n5258), .QN(
        s7_data_o[10]) );
  OA22X1 U28450 ( .IN1(n1731), .IN2(n20560), .IN3(n1626), .IN4(n20546), .Q(
        n5255) );
  OA22X1 U28451 ( .IN1(n1903), .IN2(n20594), .IN3(n1817), .IN4(n20579), .Q(
        n5256) );
  OA22X1 U28452 ( .IN1(n2075), .IN2(n20630), .IN3(n1989), .IN4(n20606), .Q(
        n5257) );
  NAND4X0 U28453 ( .IN1(n5251), .IN2(n5252), .IN3(n5253), .IN4(n5254), .QN(
        s7_data_o[11]) );
  OA22X1 U28454 ( .IN1(n1730), .IN2(n20561), .IN3(n1625), .IN4(n20546), .Q(
        n5251) );
  OA22X1 U28455 ( .IN1(n1902), .IN2(n20599), .IN3(n1816), .IN4(n20579), .Q(
        n5252) );
  OA22X1 U28456 ( .IN1(n2074), .IN2(n20631), .IN3(n1988), .IN4(n20612), .Q(
        n5253) );
  NAND4X0 U28457 ( .IN1(n5247), .IN2(n5248), .IN3(n5249), .IN4(n5250), .QN(
        s7_data_o[12]) );
  OA22X1 U28458 ( .IN1(n1729), .IN2(n20562), .IN3(n1624), .IN4(n20546), .Q(
        n5247) );
  OA22X1 U28459 ( .IN1(n1901), .IN2(n20595), .IN3(n1815), .IN4(n20579), .Q(
        n5248) );
  OA22X1 U28460 ( .IN1(n2073), .IN2(n20632), .IN3(n1987), .IN4(n20606), .Q(
        n5249) );
  NAND4X0 U28461 ( .IN1(n5243), .IN2(n5244), .IN3(n5245), .IN4(n5246), .QN(
        s7_data_o[13]) );
  OA22X1 U28462 ( .IN1(n1728), .IN2(n20563), .IN3(n1623), .IN4(n20547), .Q(
        n5243) );
  OA22X1 U28463 ( .IN1(n1900), .IN2(n20596), .IN3(n1814), .IN4(n20573), .Q(
        n5244) );
  OA22X1 U28464 ( .IN1(n2072), .IN2(n20629), .IN3(n1986), .IN4(n20613), .Q(
        n5245) );
  NAND4X0 U28465 ( .IN1(n5239), .IN2(n5240), .IN3(n5241), .IN4(n5242), .QN(
        s7_data_o[14]) );
  OA22X1 U28466 ( .IN1(n1727), .IN2(n20563), .IN3(n1622), .IN4(n20547), .Q(
        n5239) );
  OA22X1 U28467 ( .IN1(n1899), .IN2(n20596), .IN3(n1813), .IN4(n20578), .Q(
        n5240) );
  OA22X1 U28468 ( .IN1(n2071), .IN2(n20629), .IN3(n1985), .IN4(n20613), .Q(
        n5241) );
  NAND4X0 U28469 ( .IN1(n5235), .IN2(n5236), .IN3(n5237), .IN4(n5238), .QN(
        s7_data_o[15]) );
  OA22X1 U28470 ( .IN1(n1726), .IN2(n20563), .IN3(n1621), .IN4(n20547), .Q(
        n5235) );
  OA22X1 U28471 ( .IN1(n1898), .IN2(n20596), .IN3(n1812), .IN4(n20579), .Q(
        n5236) );
  OA22X1 U28472 ( .IN1(n2070), .IN2(n20629), .IN3(n1984), .IN4(n20613), .Q(
        n5237) );
  NAND4X0 U28473 ( .IN1(n5231), .IN2(n5232), .IN3(n5233), .IN4(n5234), .QN(
        s7_data_o[16]) );
  OA22X1 U28474 ( .IN1(n1725), .IN2(n20563), .IN3(n1620), .IN4(n20548), .Q(
        n5231) );
  OA22X1 U28475 ( .IN1(n1897), .IN2(n20596), .IN3(n1811), .IN4(n20580), .Q(
        n5232) );
  OA22X1 U28476 ( .IN1(n2069), .IN2(n20629), .IN3(n1983), .IN4(n20614), .Q(
        n5233) );
  NAND4X0 U28477 ( .IN1(n5227), .IN2(n5228), .IN3(n5229), .IN4(n5230), .QN(
        s7_data_o[17]) );
  OA22X1 U28478 ( .IN1(n1724), .IN2(n20566), .IN3(n1619), .IN4(n20548), .Q(
        n5227) );
  OA22X1 U28479 ( .IN1(n1896), .IN2(n20597), .IN3(n1810), .IN4(n20580), .Q(
        n5228) );
  OA22X1 U28480 ( .IN1(n2068), .IN2(n20630), .IN3(n1982), .IN4(n20614), .Q(
        n5229) );
  NAND4X0 U28481 ( .IN1(n5223), .IN2(n5224), .IN3(n5225), .IN4(n5226), .QN(
        s7_data_o[18]) );
  OA22X1 U28482 ( .IN1(n1723), .IN2(n20566), .IN3(n1618), .IN4(n20548), .Q(
        n5223) );
  OA22X1 U28483 ( .IN1(n1895), .IN2(n20597), .IN3(n1809), .IN4(n20580), .Q(
        n5224) );
  OA22X1 U28484 ( .IN1(n2067), .IN2(n20630), .IN3(n1981), .IN4(n20614), .Q(
        n5225) );
  NAND4X0 U28485 ( .IN1(n5219), .IN2(n5220), .IN3(n5221), .IN4(n5222), .QN(
        s7_data_o[19]) );
  OA22X1 U28486 ( .IN1(n1722), .IN2(n20561), .IN3(n1617), .IN4(n20548), .Q(
        n5219) );
  OA22X1 U28487 ( .IN1(n1894), .IN2(n20597), .IN3(n1808), .IN4(n20580), .Q(
        n5220) );
  OA22X1 U28488 ( .IN1(n2066), .IN2(n20630), .IN3(n1980), .IN4(n20614), .Q(
        n5221) );
  NAND4X0 U28489 ( .IN1(n5211), .IN2(n5212), .IN3(n5213), .IN4(n5214), .QN(
        s7_data_o[20]) );
  OA22X1 U28490 ( .IN1(n1721), .IN2(n20564), .IN3(n1616), .IN4(n20547), .Q(
        n5211) );
  OA22X1 U28491 ( .IN1(n1893), .IN2(n20598), .IN3(n1807), .IN4(n20577), .Q(
        n5212) );
  OA22X1 U28492 ( .IN1(n2065), .IN2(n20631), .IN3(n1979), .IN4(n20613), .Q(
        n5213) );
  NAND4X0 U28493 ( .IN1(n5207), .IN2(n5208), .IN3(n5209), .IN4(n5210), .QN(
        s7_data_o[21]) );
  OA22X1 U28494 ( .IN1(n1720), .IN2(n20564), .IN3(n1615), .IN4(n20549), .Q(
        n5207) );
  OA22X1 U28495 ( .IN1(n1892), .IN2(n20598), .IN3(n1806), .IN4(n20581), .Q(
        n5208) );
  OA22X1 U28496 ( .IN1(n2064), .IN2(n20631), .IN3(n1978), .IN4(n20615), .Q(
        n5209) );
  NAND4X0 U28497 ( .IN1(n5203), .IN2(n5204), .IN3(n5205), .IN4(n5206), .QN(
        s7_data_o[22]) );
  OA22X1 U28498 ( .IN1(n1719), .IN2(n20563), .IN3(n1614), .IN4(n20549), .Q(
        n5203) );
  OA22X1 U28499 ( .IN1(n1891), .IN2(n20596), .IN3(n1805), .IN4(n20581), .Q(
        n5204) );
  OA22X1 U28500 ( .IN1(n2063), .IN2(n20631), .IN3(n1977), .IN4(n20615), .Q(
        n5205) );
  NAND4X0 U28501 ( .IN1(n5199), .IN2(n5200), .IN3(n5201), .IN4(n5202), .QN(
        s7_data_o[23]) );
  OA22X1 U28502 ( .IN1(n1718), .IN2(n20562), .IN3(n1613), .IN4(n20549), .Q(
        n5199) );
  OA22X1 U28503 ( .IN1(n1890), .IN2(n20597), .IN3(n1804), .IN4(n20581), .Q(
        n5200) );
  OA22X1 U28504 ( .IN1(n2062), .IN2(n20631), .IN3(n1976), .IN4(n20615), .Q(
        n5201) );
  NAND4X0 U28505 ( .IN1(n5195), .IN2(n5196), .IN3(n5197), .IN4(n5198), .QN(
        s7_data_o[24]) );
  OA22X1 U28506 ( .IN1(n1717), .IN2(n20565), .IN3(n1612), .IN4(n20550), .Q(
        n5195) );
  OA22X1 U28507 ( .IN1(n1889), .IN2(n20595), .IN3(n1803), .IN4(n20582), .Q(
        n5196) );
  OA22X1 U28508 ( .IN1(n2061), .IN2(n20629), .IN3(n1975), .IN4(n20616), .Q(
        n5197) );
  NAND4X0 U28509 ( .IN1(n5191), .IN2(n5192), .IN3(n5193), .IN4(n5194), .QN(
        s7_data_o[25]) );
  OA22X1 U28510 ( .IN1(n1716), .IN2(n20562), .IN3(n1611), .IN4(n20550), .Q(
        n5191) );
  OA22X1 U28511 ( .IN1(n1888), .IN2(n20595), .IN3(n1802), .IN4(n20582), .Q(
        n5192) );
  OA22X1 U28512 ( .IN1(n2060), .IN2(n20628), .IN3(n1974), .IN4(n20616), .Q(
        n5193) );
  NAND4X0 U28513 ( .IN1(n5187), .IN2(n5188), .IN3(n5189), .IN4(n5190), .QN(
        s7_data_o[26]) );
  OA22X1 U28514 ( .IN1(n1715), .IN2(n20560), .IN3(n1610), .IN4(n20550), .Q(
        n5187) );
  OA22X1 U28515 ( .IN1(n1887), .IN2(n20594), .IN3(n1801), .IN4(n20582), .Q(
        n5188) );
  OA22X1 U28516 ( .IN1(n2059), .IN2(n20627), .IN3(n1973), .IN4(n20616), .Q(
        n5189) );
  NAND4X0 U28517 ( .IN1(n5183), .IN2(n5184), .IN3(n5185), .IN4(n5186), .QN(
        s7_data_o[27]) );
  OA22X1 U28518 ( .IN1(n1714), .IN2(n20565), .IN3(n1609), .IN4(n20549), .Q(
        n5183) );
  OA22X1 U28519 ( .IN1(n1886), .IN2(n20597), .IN3(n1800), .IN4(n20583), .Q(
        n5184) );
  OA22X1 U28520 ( .IN1(n2058), .IN2(n20632), .IN3(n1972), .IN4(n20617), .Q(
        n5185) );
  NAND4X0 U28521 ( .IN1(n5179), .IN2(n5180), .IN3(n5181), .IN4(n5182), .QN(
        s7_data_o[28]) );
  OA22X1 U28522 ( .IN1(n1713), .IN2(n20564), .IN3(n1608), .IN4(n20550), .Q(
        n5179) );
  OA22X1 U28523 ( .IN1(n1885), .IN2(n20598), .IN3(n1799), .IN4(n20583), .Q(
        n5180) );
  OA22X1 U28524 ( .IN1(n2057), .IN2(n20632), .IN3(n1971), .IN4(n20617), .Q(
        n5181) );
  NAND4X0 U28525 ( .IN1(n5175), .IN2(n5176), .IN3(n5177), .IN4(n5178), .QN(
        s7_data_o[29]) );
  OA22X1 U28526 ( .IN1(n1712), .IN2(n20564), .IN3(n1607), .IN4(n20549), .Q(
        n5175) );
  OA22X1 U28527 ( .IN1(n1884), .IN2(n20598), .IN3(n1798), .IN4(n20583), .Q(
        n5176) );
  OA22X1 U28528 ( .IN1(n2056), .IN2(n20632), .IN3(n1970), .IN4(n20617), .Q(
        n5177) );
  NAND4X0 U28529 ( .IN1(n5167), .IN2(n5168), .IN3(n5169), .IN4(n5170), .QN(
        s7_data_o[30]) );
  OA22X1 U28530 ( .IN1(n1711), .IN2(n20564), .IN3(n1606), .IN4(n20552), .Q(
        n5167) );
  OA22X1 U28531 ( .IN1(n1883), .IN2(n20598), .IN3(n1797), .IN4(n20585), .Q(
        n5168) );
  OA22X1 U28532 ( .IN1(n2055), .IN2(n20632), .IN3(n1969), .IN4(n20619), .Q(
        n5169) );
  NAND4X0 U28533 ( .IN1(n5163), .IN2(n5164), .IN3(n5165), .IN4(n5166), .QN(
        s7_data_o[31]) );
  OA22X1 U28534 ( .IN1(n1710), .IN2(n20563), .IN3(n1605), .IN4(n20551), .Q(
        n5163) );
  OA22X1 U28535 ( .IN1(n1882), .IN2(n20596), .IN3(n1796), .IN4(n20570), .Q(
        n5164) );
  OA22X1 U28536 ( .IN1(n2054), .IN2(n20631), .IN3(n1968), .IN4(n20618), .Q(
        n5165) );
  NAND4X0 U28537 ( .IN1(n5403), .IN2(n5404), .IN3(n5405), .IN4(n5406), .QN(
        s6_stb_o) );
  OA22X1 U28538 ( .IN1(n1795), .IN2(n5413), .IN3(n1709), .IN4(n5414), .Q(n5403) );
  OA22X1 U28539 ( .IN1(n1967), .IN2(n5411), .IN3(n1881), .IN4(n5412), .Q(n5404) );
  OA22X1 U28540 ( .IN1(n2139), .IN2(n5409), .IN3(n2053), .IN4(n5410), .Q(n5405) );
  NAND4X0 U28541 ( .IN1(n5391), .IN2(n5392), .IN3(n5393), .IN4(n5394), .QN(
        s6_we_o) );
  OA22X1 U28542 ( .IN1(n1794), .IN2(n20434), .IN3(n1708), .IN4(n20421), .Q(
        n5391) );
  OA22X1 U28543 ( .IN1(n1966), .IN2(n20460), .IN3(n1880), .IN4(n20454), .Q(
        n5392) );
  OA22X1 U28544 ( .IN1(n2138), .IN2(n20493), .IN3(n2052), .IN4(n20488), .Q(
        n5393) );
  NAND4X0 U28545 ( .IN1(n5427), .IN2(n5428), .IN3(n5429), .IN4(n5430), .QN(
        s6_sel_o[0]) );
  OA22X1 U28546 ( .IN1(n1793), .IN2(n20434), .IN3(n1707), .IN4(n20420), .Q(
        n5427) );
  OA22X1 U28547 ( .IN1(n1965), .IN2(n20467), .IN3(n1879), .IN4(n20453), .Q(
        n5428) );
  OA22X1 U28548 ( .IN1(n2137), .IN2(n20500), .IN3(n2051), .IN4(n20486), .Q(
        n5429) );
  NAND4X0 U28549 ( .IN1(n5423), .IN2(n5424), .IN3(n5425), .IN4(n5426), .QN(
        s6_sel_o[1]) );
  OA22X1 U28550 ( .IN1(n1792), .IN2(n20434), .IN3(n1706), .IN4(n20420), .Q(
        n5423) );
  OA22X1 U28551 ( .IN1(n1964), .IN2(n20467), .IN3(n1878), .IN4(n20453), .Q(
        n5424) );
  OA22X1 U28552 ( .IN1(n2136), .IN2(n20500), .IN3(n2050), .IN4(n20488), .Q(
        n5425) );
  NAND4X0 U28553 ( .IN1(n5419), .IN2(n5420), .IN3(n5421), .IN4(n5422), .QN(
        s6_sel_o[2]) );
  OA22X1 U28554 ( .IN1(n1791), .IN2(n20434), .IN3(n1705), .IN4(n20421), .Q(
        n5419) );
  OA22X1 U28555 ( .IN1(n1963), .IN2(n20467), .IN3(n1877), .IN4(n20454), .Q(
        n5420) );
  OA22X1 U28556 ( .IN1(n2135), .IN2(n20500), .IN3(n2049), .IN4(n20488), .Q(
        n5421) );
  NAND4X0 U28557 ( .IN1(n5415), .IN2(n5416), .IN3(n5417), .IN4(n5418), .QN(
        s6_sel_o[3]) );
  OA22X1 U28558 ( .IN1(n1790), .IN2(n20434), .IN3(n1704), .IN4(n20421), .Q(
        n5415) );
  OA22X1 U28559 ( .IN1(n1962), .IN2(n20467), .IN3(n1876), .IN4(n20454), .Q(
        n5416) );
  OA22X1 U28560 ( .IN1(n2134), .IN2(n20500), .IN3(n2048), .IN4(n20488), .Q(
        n5417) );
  NAND4X0 U28561 ( .IN1(n5683), .IN2(n5684), .IN3(n5685), .IN4(n5686), .QN(
        s6_addr_o[0]) );
  OA22X1 U28562 ( .IN1(n1789), .IN2(n20429), .IN3(n1703), .IN4(n20404), .Q(
        n5683) );
  OA22X1 U28563 ( .IN1(n1961), .IN2(n20460), .IN3(n1875), .IN4(n20437), .Q(
        n5684) );
  OA22X1 U28564 ( .IN1(n2133), .IN2(n20493), .IN3(n2047), .IN4(n20470), .Q(
        n5685) );
  NAND4X0 U28565 ( .IN1(n5639), .IN2(n5640), .IN3(n5641), .IN4(n5642), .QN(
        s6_addr_o[1]) );
  OA22X1 U28566 ( .IN1(n1788), .IN2(n20428), .IN3(n1702), .IN4(n20407), .Q(
        n5639) );
  OA22X1 U28567 ( .IN1(n1960), .IN2(n20462), .IN3(n1874), .IN4(n20440), .Q(
        n5640) );
  OA22X1 U28568 ( .IN1(n2132), .IN2(n20495), .IN3(n2046), .IN4(n20473), .Q(
        n5641) );
  NAND4X0 U28569 ( .IN1(n5595), .IN2(n5596), .IN3(n5597), .IN4(n5598), .QN(
        s6_addr_o[2]) );
  OA22X1 U28570 ( .IN1(n1787), .IN2(n20428), .IN3(n1701), .IN4(n20411), .Q(
        n5595) );
  OA22X1 U28571 ( .IN1(n1959), .IN2(n20462), .IN3(n1873), .IN4(n20444), .Q(
        n5596) );
  OA22X1 U28572 ( .IN1(n2131), .IN2(n20499), .IN3(n2045), .IN4(n20477), .Q(
        n5597) );
  NAND4X0 U28573 ( .IN1(n5583), .IN2(n5584), .IN3(n5585), .IN4(n5586), .QN(
        s6_addr_o[3]) );
  OA22X1 U28574 ( .IN1(n1786), .IN2(n20434), .IN3(n1699), .IN4(n20412), .Q(
        n5583) );
  OA22X1 U28575 ( .IN1(n1958), .IN2(n20467), .IN3(n1872), .IN4(n20445), .Q(
        n5584) );
  OA22X1 U28576 ( .IN1(n2130), .IN2(n20500), .IN3(n2044), .IN4(n20470), .Q(
        n5585) );
  NAND4X0 U28577 ( .IN1(n5579), .IN2(n5580), .IN3(n5581), .IN4(n5582), .QN(
        s6_addr_o[4]) );
  OA22X1 U28578 ( .IN1(n1785), .IN2(n20429), .IN3(n1697), .IN4(n20412), .Q(
        n5579) );
  OA22X1 U28579 ( .IN1(n1957), .IN2(n20460), .IN3(n1871), .IN4(n20445), .Q(
        n5580) );
  OA22X1 U28580 ( .IN1(n2129), .IN2(n20496), .IN3(n2043), .IN4(n20472), .Q(
        n5581) );
  NAND4X0 U28581 ( .IN1(n5575), .IN2(n5576), .IN3(n5577), .IN4(n5578), .QN(
        s6_addr_o[5]) );
  OA22X1 U28582 ( .IN1(n1784), .IN2(n20434), .IN3(n1696), .IN4(n20412), .Q(
        n5575) );
  OA22X1 U28583 ( .IN1(n1956), .IN2(n20467), .IN3(n1870), .IN4(n20444), .Q(
        n5576) );
  OA22X1 U28584 ( .IN1(n2128), .IN2(n20500), .IN3(n2042), .IN4(n20478), .Q(
        n5577) );
  NAND4X0 U28585 ( .IN1(n5571), .IN2(n5572), .IN3(n5573), .IN4(n5574), .QN(
        s6_addr_o[6]) );
  OA22X1 U28586 ( .IN1(n1783), .IN2(n20430), .IN3(n1679), .IN4(n20412), .Q(
        n5571) );
  OA22X1 U28587 ( .IN1(n1955), .IN2(n20463), .IN3(n1869), .IN4(n20445), .Q(
        n5572) );
  OA22X1 U28588 ( .IN1(n2127), .IN2(n20497), .IN3(n2041), .IN4(n20478), .Q(
        n5573) );
  NAND4X0 U28589 ( .IN1(n5567), .IN2(n5568), .IN3(n5569), .IN4(n5570), .QN(
        s6_addr_o[7]) );
  OA22X1 U28590 ( .IN1(n1782), .IN2(n20430), .IN3(n1678), .IN4(n20412), .Q(
        n5567) );
  OA22X1 U28591 ( .IN1(n1954), .IN2(n20463), .IN3(n1868), .IN4(n20437), .Q(
        n5568) );
  OA22X1 U28592 ( .IN1(n2126), .IN2(n20497), .IN3(n2040), .IN4(n20478), .Q(
        n5569) );
  NAND4X0 U28593 ( .IN1(n5563), .IN2(n5564), .IN3(n5565), .IN4(n5566), .QN(
        s6_addr_o[8]) );
  OA22X1 U28594 ( .IN1(n1781), .IN2(n20430), .IN3(n1677), .IN4(n20413), .Q(
        n5563) );
  OA22X1 U28595 ( .IN1(n1953), .IN2(n20463), .IN3(n1867), .IN4(n20446), .Q(
        n5564) );
  OA22X1 U28596 ( .IN1(n2125), .IN2(n20497), .IN3(n2039), .IN4(n20479), .Q(
        n5565) );
  NAND4X0 U28597 ( .IN1(n5559), .IN2(n5560), .IN3(n5561), .IN4(n5562), .QN(
        s6_addr_o[9]) );
  OA22X1 U28598 ( .IN1(n1780), .IN2(n20430), .IN3(n1676), .IN4(n20413), .Q(
        n5559) );
  OA22X1 U28599 ( .IN1(n1952), .IN2(n20463), .IN3(n1866), .IN4(n20446), .Q(
        n5560) );
  OA22X1 U28600 ( .IN1(n2124), .IN2(n20497), .IN3(n2038), .IN4(n20479), .Q(
        n5561) );
  NAND4X0 U28601 ( .IN1(n5679), .IN2(n5680), .IN3(n5681), .IN4(n5682), .QN(
        s6_addr_o[10]) );
  OA22X1 U28602 ( .IN1(n1779), .IN2(n20430), .IN3(n1675), .IN4(n20404), .Q(
        n5679) );
  OA22X1 U28603 ( .IN1(n1951), .IN2(n20460), .IN3(n1865), .IN4(n20437), .Q(
        n5680) );
  OA22X1 U28604 ( .IN1(n2123), .IN2(n20493), .IN3(n2037), .IN4(n20470), .Q(
        n5681) );
  NAND4X0 U28605 ( .IN1(n5675), .IN2(n5676), .IN3(n5677), .IN4(n5678), .QN(
        s6_addr_o[11]) );
  OA22X1 U28606 ( .IN1(n1778), .IN2(n20428), .IN3(n1674), .IN4(n20404), .Q(
        n5675) );
  OA22X1 U28607 ( .IN1(n1950), .IN2(n20460), .IN3(n1864), .IN4(n20437), .Q(
        n5676) );
  OA22X1 U28608 ( .IN1(n2122), .IN2(n20493), .IN3(n2036), .IN4(n20470), .Q(
        n5677) );
  NAND4X0 U28609 ( .IN1(n5671), .IN2(n5672), .IN3(n5673), .IN4(n5674), .QN(
        s6_addr_o[12]) );
  OA22X1 U28610 ( .IN1(n1777), .IN2(n20427), .IN3(n1673), .IN4(n20405), .Q(
        n5671) );
  OA22X1 U28611 ( .IN1(n1949), .IN2(n20460), .IN3(n1863), .IN4(n20438), .Q(
        n5672) );
  OA22X1 U28612 ( .IN1(n2121), .IN2(n20493), .IN3(n2035), .IN4(n20471), .Q(
        n5673) );
  NAND4X0 U28613 ( .IN1(n5667), .IN2(n5668), .IN3(n5669), .IN4(n5670), .QN(
        s6_addr_o[13]) );
  OA22X1 U28614 ( .IN1(n1776), .IN2(n20427), .IN3(n1672), .IN4(n20405), .Q(
        n5667) );
  OA22X1 U28615 ( .IN1(n1948), .IN2(n20461), .IN3(n1862), .IN4(n20438), .Q(
        n5668) );
  OA22X1 U28616 ( .IN1(n2120), .IN2(n20494), .IN3(n2034), .IN4(n20471), .Q(
        n5669) );
  NAND4X0 U28617 ( .IN1(n5663), .IN2(n5664), .IN3(n5665), .IN4(n5666), .QN(
        s6_addr_o[14]) );
  OA22X1 U28618 ( .IN1(n1775), .IN2(n20427), .IN3(n1671), .IN4(n20405), .Q(
        n5663) );
  OA22X1 U28619 ( .IN1(n1947), .IN2(n20461), .IN3(n1861), .IN4(n20438), .Q(
        n5664) );
  OA22X1 U28620 ( .IN1(n2119), .IN2(n20494), .IN3(n2033), .IN4(n20471), .Q(
        n5665) );
  NAND4X0 U28621 ( .IN1(n5659), .IN2(n5660), .IN3(n5661), .IN4(n5662), .QN(
        s6_addr_o[15]) );
  OA22X1 U28622 ( .IN1(n1774), .IN2(n20427), .IN3(n1670), .IN4(n20406), .Q(
        n5659) );
  OA22X1 U28623 ( .IN1(n1946), .IN2(n20461), .IN3(n1860), .IN4(n20439), .Q(
        n5660) );
  OA22X1 U28624 ( .IN1(n2118), .IN2(n20494), .IN3(n2032), .IN4(n20472), .Q(
        n5661) );
  NAND4X0 U28625 ( .IN1(n5655), .IN2(n5656), .IN3(n5657), .IN4(n5658), .QN(
        s6_addr_o[16]) );
  OA22X1 U28626 ( .IN1(n1773), .IN2(n20427), .IN3(n1669), .IN4(n20406), .Q(
        n5655) );
  OA22X1 U28627 ( .IN1(n1945), .IN2(n20461), .IN3(n1859), .IN4(n20439), .Q(
        n5656) );
  OA22X1 U28628 ( .IN1(n2117), .IN2(n20494), .IN3(n2031), .IN4(n20472), .Q(
        n5657) );
  NAND4X0 U28629 ( .IN1(n5651), .IN2(n5652), .IN3(n5653), .IN4(n5654), .QN(
        s6_addr_o[17]) );
  OA22X1 U28630 ( .IN1(n1772), .IN2(n20428), .IN3(n1668), .IN4(n20406), .Q(
        n5651) );
  OA22X1 U28631 ( .IN1(n1944), .IN2(n20462), .IN3(n1858), .IN4(n20439), .Q(
        n5652) );
  OA22X1 U28632 ( .IN1(n2116), .IN2(n20495), .IN3(n2030), .IN4(n20472), .Q(
        n5653) );
  NAND4X0 U28633 ( .IN1(n5647), .IN2(n5648), .IN3(n5649), .IN4(n5650), .QN(
        s6_addr_o[18]) );
  OA22X1 U28634 ( .IN1(n1771), .IN2(n20428), .IN3(n1667), .IN4(n20407), .Q(
        n5647) );
  OA22X1 U28635 ( .IN1(n1943), .IN2(n20462), .IN3(n1857), .IN4(n20440), .Q(
        n5648) );
  OA22X1 U28636 ( .IN1(n2115), .IN2(n20495), .IN3(n2029), .IN4(n20473), .Q(
        n5649) );
  NAND4X0 U28637 ( .IN1(n5643), .IN2(n5644), .IN3(n5645), .IN4(n5646), .QN(
        s6_addr_o[19]) );
  OA22X1 U28638 ( .IN1(n1770), .IN2(n20428), .IN3(n1666), .IN4(n20407), .Q(
        n5643) );
  OA22X1 U28639 ( .IN1(n1942), .IN2(n20462), .IN3(n1856), .IN4(n20440), .Q(
        n5644) );
  OA22X1 U28640 ( .IN1(n2114), .IN2(n20495), .IN3(n2028), .IN4(n20473), .Q(
        n5645) );
  NAND4X0 U28641 ( .IN1(n5635), .IN2(n5636), .IN3(n5637), .IN4(n5638), .QN(
        s6_addr_o[20]) );
  OA22X1 U28642 ( .IN1(n1769), .IN2(n20427), .IN3(n1665), .IN4(n20408), .Q(
        n5635) );
  OA22X1 U28643 ( .IN1(n1941), .IN2(n20461), .IN3(n1855), .IN4(n20441), .Q(
        n5636) );
  OA22X1 U28644 ( .IN1(n2113), .IN2(n20494), .IN3(n2027), .IN4(n20474), .Q(
        n5637) );
  NAND4X0 U28645 ( .IN1(n5631), .IN2(n5632), .IN3(n5633), .IN4(n5634), .QN(
        s6_addr_o[21]) );
  OA22X1 U28646 ( .IN1(n1768), .IN2(n20427), .IN3(n1664), .IN4(n20408), .Q(
        n5631) );
  OA22X1 U28647 ( .IN1(n1940), .IN2(n20461), .IN3(n1854), .IN4(n20441), .Q(
        n5632) );
  OA22X1 U28648 ( .IN1(n2112), .IN2(n20494), .IN3(n2026), .IN4(n20474), .Q(
        n5633) );
  NAND4X0 U28649 ( .IN1(n5627), .IN2(n5628), .IN3(n5629), .IN4(n5630), .QN(
        s6_addr_o[22]) );
  OA22X1 U28650 ( .IN1(n1767), .IN2(n20429), .IN3(n1663), .IN4(n20408), .Q(
        n5627) );
  OA22X1 U28651 ( .IN1(n1939), .IN2(n20460), .IN3(n1853), .IN4(n20441), .Q(
        n5628) );
  OA22X1 U28652 ( .IN1(n2111), .IN2(n20493), .IN3(n2025), .IN4(n20474), .Q(
        n5629) );
  NAND4X0 U28653 ( .IN1(n5623), .IN2(n5624), .IN3(n5625), .IN4(n5626), .QN(
        s6_addr_o[23]) );
  OA22X1 U28654 ( .IN1(n1766), .IN2(n20427), .IN3(n1662), .IN4(n20409), .Q(
        n5623) );
  OA22X1 U28655 ( .IN1(n1938), .IN2(n20461), .IN3(n1852), .IN4(n20442), .Q(
        n5624) );
  OA22X1 U28656 ( .IN1(n2110), .IN2(n20494), .IN3(n2024), .IN4(n20475), .Q(
        n5625) );
  NAND4X0 U28657 ( .IN1(n5619), .IN2(n5620), .IN3(n5621), .IN4(n5622), .QN(
        s6_addr_o[24]) );
  OA22X1 U28658 ( .IN1(n1765), .IN2(n20429), .IN3(n1661), .IN4(n20409), .Q(
        n5619) );
  OA22X1 U28659 ( .IN1(n1937), .IN2(n20467), .IN3(n1851), .IN4(n20442), .Q(
        n5620) );
  OA22X1 U28660 ( .IN1(n2109), .IN2(n20496), .IN3(n2023), .IN4(n20475), .Q(
        n5621) );
  NAND4X0 U28661 ( .IN1(n5615), .IN2(n5616), .IN3(n5617), .IN4(n5618), .QN(
        s6_addr_o[25]) );
  OA22X1 U28662 ( .IN1(n1764), .IN2(n20429), .IN3(n1660), .IN4(n20409), .Q(
        n5615) );
  OA22X1 U28663 ( .IN1(n1936), .IN2(n20463), .IN3(n1850), .IN4(n20442), .Q(
        n5616) );
  OA22X1 U28664 ( .IN1(n2108), .IN2(n20496), .IN3(n2022), .IN4(n20475), .Q(
        n5617) );
  NAND4X0 U28665 ( .IN1(n5611), .IN2(n5612), .IN3(n5613), .IN4(n5614), .QN(
        s6_addr_o[26]) );
  OA22X1 U28666 ( .IN1(n1763), .IN2(n20429), .IN3(n1659), .IN4(n20410), .Q(
        n5611) );
  OA22X1 U28667 ( .IN1(n1935), .IN2(n20462), .IN3(n1849), .IN4(n20443), .Q(
        n5612) );
  OA22X1 U28668 ( .IN1(n2107), .IN2(n20496), .IN3(n2021), .IN4(n20476), .Q(
        n5613) );
  NAND4X0 U28669 ( .IN1(n5607), .IN2(n5608), .IN3(n5609), .IN4(n5610), .QN(
        s6_addr_o[27]) );
  OA22X1 U28670 ( .IN1(n1762), .IN2(n20429), .IN3(n1658), .IN4(n20410), .Q(
        n5607) );
  OA22X1 U28671 ( .IN1(n1934), .IN2(n20461), .IN3(n1848), .IN4(n20443), .Q(
        n5608) );
  OA22X1 U28672 ( .IN1(n2106), .IN2(n20496), .IN3(n2020), .IN4(n20476), .Q(
        n5609) );
  NAND4X0 U28673 ( .IN1(n5603), .IN2(n5604), .IN3(n5605), .IN4(n5606), .QN(
        s6_addr_o[28]) );
  OA22X1 U28674 ( .IN1(n1761), .IN2(n20427), .IN3(n1657), .IN4(n20410), .Q(
        n5603) );
  OA22X1 U28675 ( .IN1(n1933), .IN2(n20461), .IN3(n1847), .IN4(n20443), .Q(
        n5604) );
  OA22X1 U28676 ( .IN1(n2105), .IN2(n20500), .IN3(n2019), .IN4(n20476), .Q(
        n5605) );
  NAND4X0 U28677 ( .IN1(n5599), .IN2(n5600), .IN3(n5601), .IN4(n5602), .QN(
        s6_addr_o[29]) );
  OA22X1 U28678 ( .IN1(n1760), .IN2(n20433), .IN3(n1656), .IN4(n20411), .Q(
        n5599) );
  OA22X1 U28679 ( .IN1(n1932), .IN2(n20465), .IN3(n1846), .IN4(n20444), .Q(
        n5600) );
  OA22X1 U28680 ( .IN1(n2104), .IN2(n20496), .IN3(n2018), .IN4(n20477), .Q(
        n5601) );
  NAND4X0 U28681 ( .IN1(n5591), .IN2(n5592), .IN3(n5593), .IN4(n5594), .QN(
        s6_addr_o[30]) );
  OA22X1 U28682 ( .IN1(n1759), .IN2(n20432), .IN3(n1655), .IN4(n20411), .Q(
        n5591) );
  OA22X1 U28683 ( .IN1(n1931), .IN2(n20466), .IN3(n1845), .IN4(n20444), .Q(
        n5592) );
  OA22X1 U28684 ( .IN1(n2103), .IN2(n20496), .IN3(n2017), .IN4(n20477), .Q(
        n5593) );
  NAND4X0 U28685 ( .IN1(n5587), .IN2(n5588), .IN3(n5589), .IN4(n5590), .QN(
        s6_addr_o[31]) );
  OA22X1 U28686 ( .IN1(n1758), .IN2(n20431), .IN3(n1650), .IN4(n20411), .Q(
        n5587) );
  OA22X1 U28687 ( .IN1(n1930), .IN2(n20464), .IN3(n1844), .IN4(n20445), .Q(
        n5588) );
  OA22X1 U28688 ( .IN1(n2102), .IN2(n20500), .IN3(n2016), .IN4(n20488), .Q(
        n5589) );
  NAND4X0 U28689 ( .IN1(n5555), .IN2(n5556), .IN3(n5557), .IN4(n5558), .QN(
        s6_data_o[0]) );
  OA22X1 U28690 ( .IN1(n1741), .IN2(n20430), .IN3(n1636), .IN4(n20413), .Q(
        n5555) );
  OA22X1 U28691 ( .IN1(n1913), .IN2(n20463), .IN3(n1827), .IN4(n20446), .Q(
        n5556) );
  OA22X1 U28692 ( .IN1(n2085), .IN2(n20497), .IN3(n1999), .IN4(n20479), .Q(
        n5557) );
  NAND4X0 U28693 ( .IN1(n5511), .IN2(n5512), .IN3(n5513), .IN4(n5514), .QN(
        s6_data_o[1]) );
  OA22X1 U28694 ( .IN1(n1740), .IN2(n20428), .IN3(n1635), .IN4(n20415), .Q(
        n5511) );
  OA22X1 U28695 ( .IN1(n1912), .IN2(n20465), .IN3(n1826), .IN4(n20444), .Q(
        n5512) );
  OA22X1 U28696 ( .IN1(n2084), .IN2(n20499), .IN3(n1998), .IN4(n20471), .Q(
        n5513) );
  NAND4X0 U28697 ( .IN1(n5467), .IN2(n5468), .IN3(n5469), .IN4(n5470), .QN(
        s6_data_o[2]) );
  OA22X1 U28698 ( .IN1(n1739), .IN2(n20432), .IN3(n1634), .IN4(n20419), .Q(
        n5467) );
  OA22X1 U28699 ( .IN1(n1911), .IN2(n20466), .IN3(n1825), .IN4(n20437), .Q(
        n5468) );
  OA22X1 U28700 ( .IN1(n2083), .IN2(n20494), .IN3(n1997), .IN4(n20486), .Q(
        n5469) );
  NAND4X0 U28701 ( .IN1(n5455), .IN2(n5456), .IN3(n5457), .IN4(n5458), .QN(
        s6_data_o[3]) );
  OA22X1 U28702 ( .IN1(n1738), .IN2(n20431), .IN3(n1633), .IN4(n20419), .Q(
        n5455) );
  OA22X1 U28703 ( .IN1(n1910), .IN2(n20464), .IN3(n1824), .IN4(n20439), .Q(
        n5456) );
  OA22X1 U28704 ( .IN1(n2082), .IN2(n20498), .IN3(n1996), .IN4(n20486), .Q(
        n5457) );
  NAND4X0 U28705 ( .IN1(n5451), .IN2(n5452), .IN3(n5453), .IN4(n5454), .QN(
        s6_data_o[4]) );
  OA22X1 U28706 ( .IN1(n1737), .IN2(n20433), .IN3(n1632), .IN4(n20419), .Q(
        n5451) );
  OA22X1 U28707 ( .IN1(n1909), .IN2(n20465), .IN3(n1823), .IN4(n20454), .Q(
        n5452) );
  OA22X1 U28708 ( .IN1(n2081), .IN2(n20498), .IN3(n1995), .IN4(n20486), .Q(
        n5453) );
  NAND4X0 U28709 ( .IN1(n5447), .IN2(n5448), .IN3(n5449), .IN4(n5450), .QN(
        s6_data_o[5]) );
  OA22X1 U28710 ( .IN1(n1736), .IN2(n20432), .IN3(n1631), .IN4(n20419), .Q(
        n5447) );
  OA22X1 U28711 ( .IN1(n1908), .IN2(n20466), .IN3(n1822), .IN4(n20452), .Q(
        n5448) );
  OA22X1 U28712 ( .IN1(n2080), .IN2(n20498), .IN3(n1994), .IN4(n20486), .Q(
        n5449) );
  NAND4X0 U28713 ( .IN1(n5443), .IN2(n5444), .IN3(n5445), .IN4(n5446), .QN(
        s6_data_o[6]) );
  OA22X1 U28714 ( .IN1(n1735), .IN2(n20433), .IN3(n1630), .IN4(n20421), .Q(
        n5443) );
  OA22X1 U28715 ( .IN1(n1907), .IN2(n20462), .IN3(n1821), .IN4(n20452), .Q(
        n5444) );
  OA22X1 U28716 ( .IN1(n2079), .IN2(n20499), .IN3(n1993), .IN4(n20487), .Q(
        n5445) );
  NAND4X0 U28717 ( .IN1(n5439), .IN2(n5440), .IN3(n5441), .IN4(n5442), .QN(
        s6_data_o[7]) );
  OA22X1 U28718 ( .IN1(n1734), .IN2(n20433), .IN3(n1629), .IN4(n20421), .Q(
        n5439) );
  OA22X1 U28719 ( .IN1(n1906), .IN2(n20460), .IN3(n1820), .IN4(n20452), .Q(
        n5440) );
  OA22X1 U28720 ( .IN1(n2078), .IN2(n20499), .IN3(n1992), .IN4(n20487), .Q(
        n5441) );
  NAND4X0 U28721 ( .IN1(n5435), .IN2(n5436), .IN3(n5437), .IN4(n5438), .QN(
        s6_data_o[8]) );
  OA22X1 U28722 ( .IN1(n1733), .IN2(n20433), .IN3(n1628), .IN4(n20421), .Q(
        n5435) );
  OA22X1 U28723 ( .IN1(n1905), .IN2(n20467), .IN3(n1819), .IN4(n20452), .Q(
        n5436) );
  OA22X1 U28724 ( .IN1(n2077), .IN2(n20499), .IN3(n1991), .IN4(n20487), .Q(
        n5437) );
  NAND4X0 U28725 ( .IN1(n5431), .IN2(n5432), .IN3(n5433), .IN4(n5434), .QN(
        s6_data_o[9]) );
  OA22X1 U28726 ( .IN1(n1732), .IN2(n20433), .IN3(n1627), .IN4(n20420), .Q(
        n5431) );
  OA22X1 U28727 ( .IN1(n1904), .IN2(n20460), .IN3(n1818), .IN4(n20453), .Q(
        n5432) );
  OA22X1 U28728 ( .IN1(n2076), .IN2(n20499), .IN3(n1990), .IN4(n20470), .Q(
        n5433) );
  NAND4X0 U28729 ( .IN1(n5551), .IN2(n5552), .IN3(n5553), .IN4(n5554), .QN(
        s6_data_o[10]) );
  OA22X1 U28730 ( .IN1(n1731), .IN2(n20428), .IN3(n1626), .IN4(n20414), .Q(
        n5551) );
  OA22X1 U28731 ( .IN1(n1903), .IN2(n20462), .IN3(n1817), .IN4(n20447), .Q(
        n5552) );
  OA22X1 U28732 ( .IN1(n2075), .IN2(n20495), .IN3(n1989), .IN4(n20480), .Q(
        n5553) );
  NAND4X0 U28733 ( .IN1(n5547), .IN2(n5548), .IN3(n5549), .IN4(n5550), .QN(
        s6_data_o[11]) );
  OA22X1 U28734 ( .IN1(n1730), .IN2(n20429), .IN3(n1625), .IN4(n20414), .Q(
        n5547) );
  OA22X1 U28735 ( .IN1(n1902), .IN2(n20467), .IN3(n1816), .IN4(n20447), .Q(
        n5548) );
  OA22X1 U28736 ( .IN1(n2074), .IN2(n20496), .IN3(n1988), .IN4(n20480), .Q(
        n5549) );
  NAND4X0 U28737 ( .IN1(n5543), .IN2(n5544), .IN3(n5545), .IN4(n5546), .QN(
        s6_data_o[12]) );
  OA22X1 U28738 ( .IN1(n1729), .IN2(n20430), .IN3(n1624), .IN4(n20414), .Q(
        n5543) );
  OA22X1 U28739 ( .IN1(n1901), .IN2(n20463), .IN3(n1815), .IN4(n20447), .Q(
        n5544) );
  OA22X1 U28740 ( .IN1(n2073), .IN2(n20498), .IN3(n1987), .IN4(n20480), .Q(
        n5545) );
  NAND4X0 U28741 ( .IN1(n5539), .IN2(n5540), .IN3(n5541), .IN4(n5542), .QN(
        s6_data_o[13]) );
  OA22X1 U28742 ( .IN1(n1728), .IN2(n20431), .IN3(n1623), .IN4(n20415), .Q(
        n5539) );
  OA22X1 U28743 ( .IN1(n1900), .IN2(n20464), .IN3(n1814), .IN4(n20441), .Q(
        n5540) );
  OA22X1 U28744 ( .IN1(n2072), .IN2(n20498), .IN3(n1986), .IN4(n20481), .Q(
        n5541) );
  NAND4X0 U28745 ( .IN1(n5535), .IN2(n5536), .IN3(n5537), .IN4(n5538), .QN(
        s6_data_o[14]) );
  OA22X1 U28746 ( .IN1(n1727), .IN2(n20431), .IN3(n1622), .IN4(n20415), .Q(
        n5535) );
  OA22X1 U28747 ( .IN1(n1899), .IN2(n20464), .IN3(n1813), .IN4(n20446), .Q(
        n5536) );
  OA22X1 U28748 ( .IN1(n2071), .IN2(n20498), .IN3(n1985), .IN4(n20481), .Q(
        n5537) );
  NAND4X0 U28749 ( .IN1(n5531), .IN2(n5532), .IN3(n5533), .IN4(n5534), .QN(
        s6_data_o[15]) );
  OA22X1 U28750 ( .IN1(n1726), .IN2(n20431), .IN3(n1621), .IN4(n20415), .Q(
        n5531) );
  OA22X1 U28751 ( .IN1(n1898), .IN2(n20464), .IN3(n1812), .IN4(n20447), .Q(
        n5532) );
  OA22X1 U28752 ( .IN1(n2070), .IN2(n20498), .IN3(n1984), .IN4(n20481), .Q(
        n5533) );
  NAND4X0 U28753 ( .IN1(n5527), .IN2(n5528), .IN3(n5529), .IN4(n5530), .QN(
        s6_data_o[16]) );
  OA22X1 U28754 ( .IN1(n1725), .IN2(n20431), .IN3(n1620), .IN4(n20416), .Q(
        n5527) );
  OA22X1 U28755 ( .IN1(n1897), .IN2(n20464), .IN3(n1811), .IN4(n20448), .Q(
        n5528) );
  OA22X1 U28756 ( .IN1(n2069), .IN2(n20498), .IN3(n1983), .IN4(n20482), .Q(
        n5529) );
  NAND4X0 U28757 ( .IN1(n5523), .IN2(n5524), .IN3(n5525), .IN4(n5526), .QN(
        s6_data_o[17]) );
  OA22X1 U28758 ( .IN1(n1724), .IN2(n20434), .IN3(n1619), .IN4(n20416), .Q(
        n5523) );
  OA22X1 U28759 ( .IN1(n1896), .IN2(n20465), .IN3(n1810), .IN4(n20448), .Q(
        n5524) );
  OA22X1 U28760 ( .IN1(n2068), .IN2(n20497), .IN3(n1982), .IN4(n20482), .Q(
        n5525) );
  NAND4X0 U28761 ( .IN1(n5519), .IN2(n5520), .IN3(n5521), .IN4(n5522), .QN(
        s6_data_o[18]) );
  OA22X1 U28762 ( .IN1(n1723), .IN2(n20434), .IN3(n1618), .IN4(n20416), .Q(
        n5519) );
  OA22X1 U28763 ( .IN1(n1895), .IN2(n20465), .IN3(n1809), .IN4(n20448), .Q(
        n5520) );
  OA22X1 U28764 ( .IN1(n2067), .IN2(n20495), .IN3(n1981), .IN4(n20482), .Q(
        n5521) );
  NAND4X0 U28765 ( .IN1(n5515), .IN2(n5516), .IN3(n5517), .IN4(n5518), .QN(
        s6_data_o[19]) );
  OA22X1 U28766 ( .IN1(n1722), .IN2(n20429), .IN3(n1617), .IN4(n20416), .Q(
        n5515) );
  OA22X1 U28767 ( .IN1(n1894), .IN2(n20465), .IN3(n1808), .IN4(n20448), .Q(
        n5516) );
  OA22X1 U28768 ( .IN1(n2066), .IN2(n20493), .IN3(n1980), .IN4(n20472), .Q(
        n5517) );
  NAND4X0 U28769 ( .IN1(n5507), .IN2(n5508), .IN3(n5509), .IN4(n5510), .QN(
        s6_data_o[20]) );
  OA22X1 U28770 ( .IN1(n1721), .IN2(n20432), .IN3(n1616), .IN4(n20415), .Q(
        n5507) );
  OA22X1 U28771 ( .IN1(n1893), .IN2(n20466), .IN3(n1807), .IN4(n20445), .Q(
        n5508) );
  OA22X1 U28772 ( .IN1(n2065), .IN2(n20495), .IN3(n1979), .IN4(n20471), .Q(
        n5509) );
  NAND4X0 U28773 ( .IN1(n5503), .IN2(n5504), .IN3(n5505), .IN4(n5506), .QN(
        s6_data_o[21]) );
  OA22X1 U28774 ( .IN1(n1720), .IN2(n20432), .IN3(n1615), .IN4(n20417), .Q(
        n5503) );
  OA22X1 U28775 ( .IN1(n1892), .IN2(n20466), .IN3(n1806), .IN4(n20449), .Q(
        n5504) );
  OA22X1 U28776 ( .IN1(n2064), .IN2(n20493), .IN3(n1978), .IN4(n20483), .Q(
        n5505) );
  NAND4X0 U28777 ( .IN1(n5499), .IN2(n5500), .IN3(n5501), .IN4(n5502), .QN(
        s6_data_o[22]) );
  OA22X1 U28778 ( .IN1(n1719), .IN2(n20431), .IN3(n1614), .IN4(n20417), .Q(
        n5499) );
  OA22X1 U28779 ( .IN1(n1891), .IN2(n20464), .IN3(n1805), .IN4(n20449), .Q(
        n5500) );
  OA22X1 U28780 ( .IN1(n2063), .IN2(n20500), .IN3(n1977), .IN4(n20483), .Q(
        n5501) );
  NAND4X0 U28781 ( .IN1(n5495), .IN2(n5496), .IN3(n5497), .IN4(n5498), .QN(
        s6_data_o[23]) );
  OA22X1 U28782 ( .IN1(n1718), .IN2(n20430), .IN3(n1613), .IN4(n20417), .Q(
        n5495) );
  OA22X1 U28783 ( .IN1(n1890), .IN2(n20465), .IN3(n1804), .IN4(n20449), .Q(
        n5496) );
  OA22X1 U28784 ( .IN1(n2062), .IN2(n20496), .IN3(n1976), .IN4(n20483), .Q(
        n5497) );
  NAND4X0 U28785 ( .IN1(n5491), .IN2(n5492), .IN3(n5493), .IN4(n5494), .QN(
        s6_data_o[24]) );
  OA22X1 U28786 ( .IN1(n1717), .IN2(n20433), .IN3(n1612), .IN4(n20418), .Q(
        n5491) );
  OA22X1 U28787 ( .IN1(n1889), .IN2(n20463), .IN3(n1803), .IN4(n20450), .Q(
        n5492) );
  OA22X1 U28788 ( .IN1(n2061), .IN2(n20499), .IN3(n1975), .IN4(n20484), .Q(
        n5493) );
  NAND4X0 U28789 ( .IN1(n5487), .IN2(n5488), .IN3(n5489), .IN4(n5490), .QN(
        s6_data_o[25]) );
  OA22X1 U28790 ( .IN1(n1716), .IN2(n20430), .IN3(n1611), .IN4(n20418), .Q(
        n5487) );
  OA22X1 U28791 ( .IN1(n1888), .IN2(n20463), .IN3(n1802), .IN4(n20450), .Q(
        n5488) );
  OA22X1 U28792 ( .IN1(n2060), .IN2(n20497), .IN3(n1974), .IN4(n20484), .Q(
        n5489) );
  NAND4X0 U28793 ( .IN1(n5483), .IN2(n5484), .IN3(n5485), .IN4(n5486), .QN(
        s6_data_o[26]) );
  OA22X1 U28794 ( .IN1(n1715), .IN2(n20428), .IN3(n1610), .IN4(n20418), .Q(
        n5483) );
  OA22X1 U28795 ( .IN1(n1887), .IN2(n20462), .IN3(n1801), .IN4(n20450), .Q(
        n5484) );
  OA22X1 U28796 ( .IN1(n2059), .IN2(n20495), .IN3(n1973), .IN4(n20484), .Q(
        n5485) );
  NAND4X0 U28797 ( .IN1(n5479), .IN2(n5480), .IN3(n5481), .IN4(n5482), .QN(
        s6_data_o[27]) );
  OA22X1 U28798 ( .IN1(n1714), .IN2(n20433), .IN3(n1609), .IN4(n20417), .Q(
        n5479) );
  OA22X1 U28799 ( .IN1(n1886), .IN2(n20465), .IN3(n1800), .IN4(n20451), .Q(
        n5480) );
  OA22X1 U28800 ( .IN1(n2058), .IN2(n20499), .IN3(n1972), .IN4(n20485), .Q(
        n5481) );
  NAND4X0 U28801 ( .IN1(n5475), .IN2(n5476), .IN3(n5477), .IN4(n5478), .QN(
        s6_data_o[28]) );
  OA22X1 U28802 ( .IN1(n1713), .IN2(n20432), .IN3(n1608), .IN4(n20418), .Q(
        n5475) );
  OA22X1 U28803 ( .IN1(n1885), .IN2(n20466), .IN3(n1799), .IN4(n20451), .Q(
        n5476) );
  OA22X1 U28804 ( .IN1(n2057), .IN2(n20499), .IN3(n1971), .IN4(n20485), .Q(
        n5477) );
  NAND4X0 U28805 ( .IN1(n5471), .IN2(n5472), .IN3(n5473), .IN4(n5474), .QN(
        s6_data_o[29]) );
  OA22X1 U28806 ( .IN1(n1712), .IN2(n20432), .IN3(n1607), .IN4(n20417), .Q(
        n5471) );
  OA22X1 U28807 ( .IN1(n1884), .IN2(n20466), .IN3(n1798), .IN4(n20451), .Q(
        n5472) );
  OA22X1 U28808 ( .IN1(n2056), .IN2(n20498), .IN3(n1970), .IN4(n20485), .Q(
        n5473) );
  NAND4X0 U28809 ( .IN1(n5463), .IN2(n5464), .IN3(n5465), .IN4(n5466), .QN(
        s6_data_o[30]) );
  OA22X1 U28810 ( .IN1(n1711), .IN2(n20432), .IN3(n1606), .IN4(n20420), .Q(
        n5463) );
  OA22X1 U28811 ( .IN1(n1883), .IN2(n20466), .IN3(n1797), .IN4(n20453), .Q(
        n5464) );
  OA22X1 U28812 ( .IN1(n2055), .IN2(n20494), .IN3(n1969), .IN4(n20486), .Q(
        n5465) );
  NAND4X0 U28813 ( .IN1(n5459), .IN2(n5460), .IN3(n5461), .IN4(n5462), .QN(
        s6_data_o[31]) );
  OA22X1 U28814 ( .IN1(n1710), .IN2(n20431), .IN3(n1605), .IN4(n20419), .Q(
        n5459) );
  OA22X1 U28815 ( .IN1(n1882), .IN2(n20464), .IN3(n1796), .IN4(n20438), .Q(
        n5460) );
  OA22X1 U28816 ( .IN1(n2054), .IN2(n20497), .IN3(n1968), .IN4(n20486), .Q(
        n5461) );
  NAND4X0 U28817 ( .IN1(n5699), .IN2(n5700), .IN3(n5701), .IN4(n5702), .QN(
        s5_stb_o) );
  OA22X1 U28818 ( .IN1(n1795), .IN2(n5709), .IN3(n1709), .IN4(n5710), .Q(n5699) );
  OA22X1 U28819 ( .IN1(n1967), .IN2(n5707), .IN3(n1881), .IN4(n5708), .Q(n5700) );
  OA22X1 U28820 ( .IN1(n2139), .IN2(n5705), .IN3(n2053), .IN4(n5706), .Q(n5701) );
  NAND4X0 U28821 ( .IN1(n5687), .IN2(n5688), .IN3(n5689), .IN4(n5690), .QN(
        s5_we_o) );
  OA22X1 U28822 ( .IN1(n1794), .IN2(n20302), .IN3(n1708), .IN4(n20289), .Q(
        n5687) );
  OA22X1 U28823 ( .IN1(n1966), .IN2(n20328), .IN3(n1880), .IN4(n20322), .Q(
        n5688) );
  OA22X1 U28824 ( .IN1(n2138), .IN2(n20361), .IN3(n2052), .IN4(n20355), .Q(
        n5689) );
  NAND4X0 U28825 ( .IN1(n5723), .IN2(n5724), .IN3(n5725), .IN4(n5726), .QN(
        s5_sel_o[0]) );
  OA22X1 U28826 ( .IN1(n1793), .IN2(n20302), .IN3(n1707), .IN4(n20288), .Q(
        n5723) );
  OA22X1 U28827 ( .IN1(n1965), .IN2(n20335), .IN3(n1879), .IN4(n20321), .Q(
        n5724) );
  OA22X1 U28828 ( .IN1(n2137), .IN2(n20368), .IN3(n2051), .IN4(n20354), .Q(
        n5725) );
  NAND4X0 U28829 ( .IN1(n5719), .IN2(n5720), .IN3(n5721), .IN4(n5722), .QN(
        s5_sel_o[1]) );
  OA22X1 U28830 ( .IN1(n1792), .IN2(n20302), .IN3(n1706), .IN4(n20288), .Q(
        n5719) );
  OA22X1 U28831 ( .IN1(n1964), .IN2(n20335), .IN3(n1878), .IN4(n20321), .Q(
        n5720) );
  OA22X1 U28832 ( .IN1(n2136), .IN2(n20368), .IN3(n2050), .IN4(n20354), .Q(
        n5721) );
  NAND4X0 U28833 ( .IN1(n5715), .IN2(n5716), .IN3(n5717), .IN4(n5718), .QN(
        s5_sel_o[2]) );
  OA22X1 U28834 ( .IN1(n1791), .IN2(n20302), .IN3(n1705), .IN4(n20289), .Q(
        n5715) );
  OA22X1 U28835 ( .IN1(n1963), .IN2(n20335), .IN3(n1877), .IN4(n20322), .Q(
        n5716) );
  OA22X1 U28836 ( .IN1(n2135), .IN2(n20368), .IN3(n2049), .IN4(n20355), .Q(
        n5717) );
  NAND4X0 U28837 ( .IN1(n5711), .IN2(n5712), .IN3(n5713), .IN4(n5714), .QN(
        s5_sel_o[3]) );
  OA22X1 U28838 ( .IN1(n1790), .IN2(n20302), .IN3(n1704), .IN4(n20289), .Q(
        n5711) );
  OA22X1 U28839 ( .IN1(n1962), .IN2(n20335), .IN3(n1876), .IN4(n20322), .Q(
        n5712) );
  OA22X1 U28840 ( .IN1(n2134), .IN2(n20368), .IN3(n2048), .IN4(n20355), .Q(
        n5713) );
  NAND4X0 U28841 ( .IN1(n5979), .IN2(n5980), .IN3(n5981), .IN4(n5982), .QN(
        s5_addr_o[0]) );
  OA22X1 U28842 ( .IN1(n1789), .IN2(n20297), .IN3(n1703), .IN4(n20272), .Q(
        n5979) );
  OA22X1 U28843 ( .IN1(n1961), .IN2(n20328), .IN3(n1875), .IN4(n20305), .Q(
        n5980) );
  OA22X1 U28844 ( .IN1(n2133), .IN2(n20361), .IN3(n2047), .IN4(n20338), .Q(
        n5981) );
  NAND4X0 U28845 ( .IN1(n5935), .IN2(n5936), .IN3(n5937), .IN4(n5938), .QN(
        s5_addr_o[1]) );
  OA22X1 U28846 ( .IN1(n1788), .IN2(n20296), .IN3(n1702), .IN4(n20275), .Q(
        n5935) );
  OA22X1 U28847 ( .IN1(n1960), .IN2(n20330), .IN3(n1874), .IN4(n20308), .Q(
        n5936) );
  OA22X1 U28848 ( .IN1(n2132), .IN2(n20363), .IN3(n2046), .IN4(n20341), .Q(
        n5937) );
  NAND4X0 U28849 ( .IN1(n5891), .IN2(n5892), .IN3(n5893), .IN4(n5894), .QN(
        s5_addr_o[2]) );
  OA22X1 U28850 ( .IN1(n1787), .IN2(n20296), .IN3(n1701), .IN4(n20279), .Q(
        n5891) );
  OA22X1 U28851 ( .IN1(n1959), .IN2(n20330), .IN3(n1873), .IN4(n20312), .Q(
        n5892) );
  OA22X1 U28852 ( .IN1(n2131), .IN2(n20363), .IN3(n2045), .IN4(n20345), .Q(
        n5893) );
  NAND4X0 U28853 ( .IN1(n5879), .IN2(n5880), .IN3(n5881), .IN4(n5882), .QN(
        s5_addr_o[3]) );
  OA22X1 U28854 ( .IN1(n1786), .IN2(n20302), .IN3(n1699), .IN4(n20280), .Q(
        n5879) );
  OA22X1 U28855 ( .IN1(n1958), .IN2(n20335), .IN3(n1872), .IN4(n20313), .Q(
        n5880) );
  OA22X1 U28856 ( .IN1(n2130), .IN2(n20368), .IN3(n2044), .IN4(n20346), .Q(
        n5881) );
  NAND4X0 U28857 ( .IN1(n5875), .IN2(n5876), .IN3(n5877), .IN4(n5878), .QN(
        s5_addr_o[4]) );
  OA22X1 U28858 ( .IN1(n1785), .IN2(n20297), .IN3(n1697), .IN4(n20280), .Q(
        n5875) );
  OA22X1 U28859 ( .IN1(n1957), .IN2(n20328), .IN3(n1871), .IN4(n20313), .Q(
        n5876) );
  OA22X1 U28860 ( .IN1(n2129), .IN2(n20361), .IN3(n2043), .IN4(n20346), .Q(
        n5877) );
  NAND4X0 U28861 ( .IN1(n5871), .IN2(n5872), .IN3(n5873), .IN4(n5874), .QN(
        s5_addr_o[5]) );
  OA22X1 U28862 ( .IN1(n1784), .IN2(n20302), .IN3(n1696), .IN4(n20280), .Q(
        n5871) );
  OA22X1 U28863 ( .IN1(n1956), .IN2(n20335), .IN3(n1870), .IN4(n20312), .Q(
        n5872) );
  OA22X1 U28864 ( .IN1(n2128), .IN2(n20368), .IN3(n2042), .IN4(n20345), .Q(
        n5873) );
  NAND4X0 U28865 ( .IN1(n5867), .IN2(n5868), .IN3(n5869), .IN4(n5870), .QN(
        s5_addr_o[6]) );
  OA22X1 U28866 ( .IN1(n1783), .IN2(n20298), .IN3(n1679), .IN4(n20280), .Q(
        n5867) );
  OA22X1 U28867 ( .IN1(n1955), .IN2(n20331), .IN3(n1869), .IN4(n20313), .Q(
        n5868) );
  OA22X1 U28868 ( .IN1(n2127), .IN2(n20364), .IN3(n2041), .IN4(n20346), .Q(
        n5869) );
  NAND4X0 U28869 ( .IN1(n5863), .IN2(n5864), .IN3(n5865), .IN4(n5866), .QN(
        s5_addr_o[7]) );
  OA22X1 U28870 ( .IN1(n1782), .IN2(n20298), .IN3(n1678), .IN4(n20280), .Q(
        n5863) );
  OA22X1 U28871 ( .IN1(n1954), .IN2(n20331), .IN3(n1868), .IN4(n20305), .Q(
        n5864) );
  OA22X1 U28872 ( .IN1(n2126), .IN2(n20364), .IN3(n2040), .IN4(n20345), .Q(
        n5865) );
  NAND4X0 U28873 ( .IN1(n5859), .IN2(n5860), .IN3(n5861), .IN4(n5862), .QN(
        s5_addr_o[8]) );
  OA22X1 U28874 ( .IN1(n1781), .IN2(n20298), .IN3(n1677), .IN4(n20281), .Q(
        n5859) );
  OA22X1 U28875 ( .IN1(n1953), .IN2(n20331), .IN3(n1867), .IN4(n20314), .Q(
        n5860) );
  OA22X1 U28876 ( .IN1(n2125), .IN2(n20364), .IN3(n2039), .IN4(n20347), .Q(
        n5861) );
  NAND4X0 U28877 ( .IN1(n5855), .IN2(n5856), .IN3(n5857), .IN4(n5858), .QN(
        s5_addr_o[9]) );
  OA22X1 U28878 ( .IN1(n1780), .IN2(n20298), .IN3(n1676), .IN4(n20281), .Q(
        n5855) );
  OA22X1 U28879 ( .IN1(n1952), .IN2(n20331), .IN3(n1866), .IN4(n20314), .Q(
        n5856) );
  OA22X1 U28880 ( .IN1(n2124), .IN2(n20364), .IN3(n2038), .IN4(n20347), .Q(
        n5857) );
  NAND4X0 U28881 ( .IN1(n5975), .IN2(n5976), .IN3(n5977), .IN4(n5978), .QN(
        s5_addr_o[10]) );
  OA22X1 U28882 ( .IN1(n1779), .IN2(n20298), .IN3(n1675), .IN4(n20272), .Q(
        n5975) );
  OA22X1 U28883 ( .IN1(n1951), .IN2(n20328), .IN3(n1865), .IN4(n20305), .Q(
        n5976) );
  OA22X1 U28884 ( .IN1(n2123), .IN2(n20361), .IN3(n2037), .IN4(n20338), .Q(
        n5977) );
  NAND4X0 U28885 ( .IN1(n5971), .IN2(n5972), .IN3(n5973), .IN4(n5974), .QN(
        s5_addr_o[11]) );
  OA22X1 U28886 ( .IN1(n1778), .IN2(n20296), .IN3(n1674), .IN4(n20272), .Q(
        n5971) );
  OA22X1 U28887 ( .IN1(n1950), .IN2(n20328), .IN3(n1864), .IN4(n20305), .Q(
        n5972) );
  OA22X1 U28888 ( .IN1(n2122), .IN2(n20361), .IN3(n2036), .IN4(n20338), .Q(
        n5973) );
  NAND4X0 U28889 ( .IN1(n5967), .IN2(n5968), .IN3(n5969), .IN4(n5970), .QN(
        s5_addr_o[12]) );
  OA22X1 U28890 ( .IN1(n1777), .IN2(n20295), .IN3(n1673), .IN4(n20273), .Q(
        n5967) );
  OA22X1 U28891 ( .IN1(n1949), .IN2(n20328), .IN3(n1863), .IN4(n20306), .Q(
        n5968) );
  OA22X1 U28892 ( .IN1(n2121), .IN2(n20361), .IN3(n2035), .IN4(n20339), .Q(
        n5969) );
  NAND4X0 U28893 ( .IN1(n5963), .IN2(n5964), .IN3(n5965), .IN4(n5966), .QN(
        s5_addr_o[13]) );
  OA22X1 U28894 ( .IN1(n1776), .IN2(n20295), .IN3(n1672), .IN4(n20273), .Q(
        n5963) );
  OA22X1 U28895 ( .IN1(n1948), .IN2(n20329), .IN3(n1862), .IN4(n20306), .Q(
        n5964) );
  OA22X1 U28896 ( .IN1(n2120), .IN2(n20362), .IN3(n2034), .IN4(n20339), .Q(
        n5965) );
  NAND4X0 U28897 ( .IN1(n5959), .IN2(n5960), .IN3(n5961), .IN4(n5962), .QN(
        s5_addr_o[14]) );
  OA22X1 U28898 ( .IN1(n1775), .IN2(n20295), .IN3(n1671), .IN4(n20273), .Q(
        n5959) );
  OA22X1 U28899 ( .IN1(n1947), .IN2(n20329), .IN3(n1861), .IN4(n20306), .Q(
        n5960) );
  OA22X1 U28900 ( .IN1(n2119), .IN2(n20362), .IN3(n2033), .IN4(n20339), .Q(
        n5961) );
  NAND4X0 U28901 ( .IN1(n5955), .IN2(n5956), .IN3(n5957), .IN4(n5958), .QN(
        s5_addr_o[15]) );
  OA22X1 U28902 ( .IN1(n1774), .IN2(n20295), .IN3(n1670), .IN4(n20274), .Q(
        n5955) );
  OA22X1 U28903 ( .IN1(n1946), .IN2(n20329), .IN3(n1860), .IN4(n20307), .Q(
        n5956) );
  OA22X1 U28904 ( .IN1(n2118), .IN2(n20362), .IN3(n2032), .IN4(n20340), .Q(
        n5957) );
  NAND4X0 U28905 ( .IN1(n5951), .IN2(n5952), .IN3(n5953), .IN4(n5954), .QN(
        s5_addr_o[16]) );
  OA22X1 U28906 ( .IN1(n1773), .IN2(n20295), .IN3(n1669), .IN4(n20274), .Q(
        n5951) );
  OA22X1 U28907 ( .IN1(n1945), .IN2(n20329), .IN3(n1859), .IN4(n20307), .Q(
        n5952) );
  OA22X1 U28908 ( .IN1(n2117), .IN2(n20362), .IN3(n2031), .IN4(n20340), .Q(
        n5953) );
  NAND4X0 U28909 ( .IN1(n5947), .IN2(n5948), .IN3(n5949), .IN4(n5950), .QN(
        s5_addr_o[17]) );
  OA22X1 U28910 ( .IN1(n1772), .IN2(n20296), .IN3(n1668), .IN4(n20274), .Q(
        n5947) );
  OA22X1 U28911 ( .IN1(n1944), .IN2(n20330), .IN3(n1858), .IN4(n20307), .Q(
        n5948) );
  OA22X1 U28912 ( .IN1(n2116), .IN2(n20363), .IN3(n2030), .IN4(n20340), .Q(
        n5949) );
  NAND4X0 U28913 ( .IN1(n5943), .IN2(n5944), .IN3(n5945), .IN4(n5946), .QN(
        s5_addr_o[18]) );
  OA22X1 U28914 ( .IN1(n1771), .IN2(n20296), .IN3(n1667), .IN4(n20275), .Q(
        n5943) );
  OA22X1 U28915 ( .IN1(n1943), .IN2(n20330), .IN3(n1857), .IN4(n20308), .Q(
        n5944) );
  OA22X1 U28916 ( .IN1(n2115), .IN2(n20363), .IN3(n2029), .IN4(n20341), .Q(
        n5945) );
  NAND4X0 U28917 ( .IN1(n5939), .IN2(n5940), .IN3(n5941), .IN4(n5942), .QN(
        s5_addr_o[19]) );
  OA22X1 U28918 ( .IN1(n1770), .IN2(n20296), .IN3(n1666), .IN4(n20275), .Q(
        n5939) );
  OA22X1 U28919 ( .IN1(n1942), .IN2(n20330), .IN3(n1856), .IN4(n20308), .Q(
        n5940) );
  OA22X1 U28920 ( .IN1(n2114), .IN2(n20363), .IN3(n2028), .IN4(n20341), .Q(
        n5941) );
  NAND4X0 U28921 ( .IN1(n5931), .IN2(n5932), .IN3(n5933), .IN4(n5934), .QN(
        s5_addr_o[20]) );
  OA22X1 U28922 ( .IN1(n1769), .IN2(n20295), .IN3(n1665), .IN4(n20276), .Q(
        n5931) );
  OA22X1 U28923 ( .IN1(n1941), .IN2(n20329), .IN3(n1855), .IN4(n20309), .Q(
        n5932) );
  OA22X1 U28924 ( .IN1(n2113), .IN2(n20362), .IN3(n2027), .IN4(n20342), .Q(
        n5933) );
  NAND4X0 U28925 ( .IN1(n5927), .IN2(n5928), .IN3(n5929), .IN4(n5930), .QN(
        s5_addr_o[21]) );
  OA22X1 U28926 ( .IN1(n1768), .IN2(n20295), .IN3(n1664), .IN4(n20276), .Q(
        n5927) );
  OA22X1 U28927 ( .IN1(n1940), .IN2(n20329), .IN3(n1854), .IN4(n20309), .Q(
        n5928) );
  OA22X1 U28928 ( .IN1(n2112), .IN2(n20362), .IN3(n2026), .IN4(n20342), .Q(
        n5929) );
  NAND4X0 U28929 ( .IN1(n5923), .IN2(n5924), .IN3(n5925), .IN4(n5926), .QN(
        s5_addr_o[22]) );
  OA22X1 U28930 ( .IN1(n1767), .IN2(n20297), .IN3(n1663), .IN4(n20276), .Q(
        n5923) );
  OA22X1 U28931 ( .IN1(n1939), .IN2(n20328), .IN3(n1853), .IN4(n20309), .Q(
        n5924) );
  OA22X1 U28932 ( .IN1(n2111), .IN2(n20361), .IN3(n2025), .IN4(n20342), .Q(
        n5925) );
  NAND4X0 U28933 ( .IN1(n5919), .IN2(n5920), .IN3(n5921), .IN4(n5922), .QN(
        s5_addr_o[23]) );
  OA22X1 U28934 ( .IN1(n1766), .IN2(n20295), .IN3(n1662), .IN4(n20277), .Q(
        n5919) );
  OA22X1 U28935 ( .IN1(n1938), .IN2(n20329), .IN3(n1852), .IN4(n20310), .Q(
        n5920) );
  OA22X1 U28936 ( .IN1(n2110), .IN2(n20362), .IN3(n2024), .IN4(n20343), .Q(
        n5921) );
  NAND4X0 U28937 ( .IN1(n5915), .IN2(n5916), .IN3(n5917), .IN4(n5918), .QN(
        s5_addr_o[24]) );
  OA22X1 U28938 ( .IN1(n1765), .IN2(n20297), .IN3(n1661), .IN4(n20277), .Q(
        n5915) );
  OA22X1 U28939 ( .IN1(n1937), .IN2(n20335), .IN3(n1851), .IN4(n20310), .Q(
        n5916) );
  OA22X1 U28940 ( .IN1(n2109), .IN2(n20368), .IN3(n2023), .IN4(n20343), .Q(
        n5917) );
  NAND4X0 U28941 ( .IN1(n5911), .IN2(n5912), .IN3(n5913), .IN4(n5914), .QN(
        s5_addr_o[25]) );
  OA22X1 U28942 ( .IN1(n1764), .IN2(n20297), .IN3(n1660), .IN4(n20277), .Q(
        n5911) );
  OA22X1 U28943 ( .IN1(n1936), .IN2(n20331), .IN3(n1850), .IN4(n20310), .Q(
        n5912) );
  OA22X1 U28944 ( .IN1(n2108), .IN2(n20364), .IN3(n2022), .IN4(n20343), .Q(
        n5913) );
  NAND4X0 U28945 ( .IN1(n5907), .IN2(n5908), .IN3(n5909), .IN4(n5910), .QN(
        s5_addr_o[26]) );
  OA22X1 U28946 ( .IN1(n1763), .IN2(n20297), .IN3(n1659), .IN4(n20278), .Q(
        n5907) );
  OA22X1 U28947 ( .IN1(n1935), .IN2(n20330), .IN3(n1849), .IN4(n20311), .Q(
        n5908) );
  OA22X1 U28948 ( .IN1(n2107), .IN2(n20363), .IN3(n2021), .IN4(n20344), .Q(
        n5909) );
  NAND4X0 U28949 ( .IN1(n5903), .IN2(n5904), .IN3(n5905), .IN4(n5906), .QN(
        s5_addr_o[27]) );
  OA22X1 U28950 ( .IN1(n1762), .IN2(n20297), .IN3(n1658), .IN4(n20278), .Q(
        n5903) );
  OA22X1 U28951 ( .IN1(n1934), .IN2(n20329), .IN3(n1848), .IN4(n20311), .Q(
        n5904) );
  OA22X1 U28952 ( .IN1(n2106), .IN2(n20362), .IN3(n2020), .IN4(n20344), .Q(
        n5905) );
  NAND4X0 U28953 ( .IN1(n5899), .IN2(n5900), .IN3(n5901), .IN4(n5902), .QN(
        s5_addr_o[28]) );
  OA22X1 U28954 ( .IN1(n1761), .IN2(n20295), .IN3(n1657), .IN4(n20278), .Q(
        n5899) );
  OA22X1 U28955 ( .IN1(n1933), .IN2(n20329), .IN3(n1847), .IN4(n20311), .Q(
        n5900) );
  OA22X1 U28956 ( .IN1(n2105), .IN2(n20362), .IN3(n2019), .IN4(n20344), .Q(
        n5901) );
  NAND4X0 U28957 ( .IN1(n5895), .IN2(n5896), .IN3(n5897), .IN4(n5898), .QN(
        s5_addr_o[29]) );
  OA22X1 U28958 ( .IN1(n1760), .IN2(n20301), .IN3(n1656), .IN4(n20279), .Q(
        n5895) );
  OA22X1 U28959 ( .IN1(n1932), .IN2(n20333), .IN3(n1846), .IN4(n20312), .Q(
        n5896) );
  OA22X1 U28960 ( .IN1(n2104), .IN2(n20366), .IN3(n2018), .IN4(n20345), .Q(
        n5897) );
  NAND4X0 U28961 ( .IN1(n5887), .IN2(n5888), .IN3(n5889), .IN4(n5890), .QN(
        s5_addr_o[30]) );
  OA22X1 U28962 ( .IN1(n1759), .IN2(n20300), .IN3(n1655), .IN4(n20279), .Q(
        n5887) );
  OA22X1 U28963 ( .IN1(n1931), .IN2(n20334), .IN3(n1845), .IN4(n20312), .Q(
        n5888) );
  OA22X1 U28964 ( .IN1(n2103), .IN2(n20367), .IN3(n2017), .IN4(n20345), .Q(
        n5889) );
  NAND4X0 U28965 ( .IN1(n5883), .IN2(n5884), .IN3(n5885), .IN4(n5886), .QN(
        s5_addr_o[31]) );
  OA22X1 U28966 ( .IN1(n1758), .IN2(n20299), .IN3(n1650), .IN4(n20279), .Q(
        n5883) );
  OA22X1 U28967 ( .IN1(n1930), .IN2(n20332), .IN3(n1844), .IN4(n20313), .Q(
        n5884) );
  OA22X1 U28968 ( .IN1(n2102), .IN2(n20365), .IN3(n2016), .IN4(n20346), .Q(
        n5885) );
  NAND4X0 U28969 ( .IN1(n5851), .IN2(n5852), .IN3(n5853), .IN4(n5854), .QN(
        s5_data_o[0]) );
  OA22X1 U28970 ( .IN1(n1741), .IN2(n20298), .IN3(n1636), .IN4(n20281), .Q(
        n5851) );
  OA22X1 U28971 ( .IN1(n1913), .IN2(n20331), .IN3(n1827), .IN4(n20314), .Q(
        n5852) );
  OA22X1 U28972 ( .IN1(n2085), .IN2(n20364), .IN3(n1999), .IN4(n20347), .Q(
        n5853) );
  NAND4X0 U28973 ( .IN1(n5807), .IN2(n5808), .IN3(n5809), .IN4(n5810), .QN(
        s5_data_o[1]) );
  OA22X1 U28974 ( .IN1(n1740), .IN2(n20296), .IN3(n1635), .IN4(n20283), .Q(
        n5807) );
  OA22X1 U28975 ( .IN1(n1912), .IN2(n20333), .IN3(n1826), .IN4(n20312), .Q(
        n5808) );
  OA22X1 U28976 ( .IN1(n2084), .IN2(n20366), .IN3(n1998), .IN4(n20345), .Q(
        n5809) );
  NAND4X0 U28977 ( .IN1(n5763), .IN2(n5764), .IN3(n5765), .IN4(n5766), .QN(
        s5_data_o[2]) );
  OA22X1 U28978 ( .IN1(n1739), .IN2(n20300), .IN3(n1634), .IN4(n20287), .Q(
        n5763) );
  OA22X1 U28979 ( .IN1(n1911), .IN2(n20334), .IN3(n1825), .IN4(n20305), .Q(
        n5764) );
  OA22X1 U28980 ( .IN1(n2083), .IN2(n20367), .IN3(n1997), .IN4(n20338), .Q(
        n5765) );
  NAND4X0 U28981 ( .IN1(n5751), .IN2(n5752), .IN3(n5753), .IN4(n5754), .QN(
        s5_data_o[3]) );
  OA22X1 U28982 ( .IN1(n1738), .IN2(n20299), .IN3(n1633), .IN4(n20287), .Q(
        n5751) );
  OA22X1 U28983 ( .IN1(n1910), .IN2(n20332), .IN3(n1824), .IN4(n20307), .Q(
        n5752) );
  OA22X1 U28984 ( .IN1(n2082), .IN2(n20365), .IN3(n1996), .IN4(n20340), .Q(
        n5753) );
  NAND4X0 U28985 ( .IN1(n5747), .IN2(n5748), .IN3(n5749), .IN4(n5750), .QN(
        s5_data_o[4]) );
  OA22X1 U28986 ( .IN1(n1737), .IN2(n20301), .IN3(n1632), .IN4(n20287), .Q(
        n5747) );
  OA22X1 U28987 ( .IN1(n1909), .IN2(n20333), .IN3(n1823), .IN4(n20322), .Q(
        n5748) );
  OA22X1 U28988 ( .IN1(n2081), .IN2(n20366), .IN3(n1995), .IN4(n20355), .Q(
        n5749) );
  NAND4X0 U28989 ( .IN1(n5743), .IN2(n5744), .IN3(n5745), .IN4(n5746), .QN(
        s5_data_o[5]) );
  OA22X1 U28990 ( .IN1(n1736), .IN2(n20300), .IN3(n1631), .IN4(n20287), .Q(
        n5743) );
  OA22X1 U28991 ( .IN1(n1908), .IN2(n20334), .IN3(n1822), .IN4(n20320), .Q(
        n5744) );
  OA22X1 U28992 ( .IN1(n2080), .IN2(n20367), .IN3(n1994), .IN4(n20353), .Q(
        n5745) );
  NAND4X0 U28993 ( .IN1(n5739), .IN2(n5740), .IN3(n5741), .IN4(n5742), .QN(
        s5_data_o[6]) );
  OA22X1 U28994 ( .IN1(n1735), .IN2(n20301), .IN3(n1630), .IN4(n20289), .Q(
        n5739) );
  OA22X1 U28995 ( .IN1(n1907), .IN2(n20330), .IN3(n1821), .IN4(n20320), .Q(
        n5740) );
  OA22X1 U28996 ( .IN1(n2079), .IN2(n20363), .IN3(n1993), .IN4(n20353), .Q(
        n5741) );
  NAND4X0 U28997 ( .IN1(n5735), .IN2(n5736), .IN3(n5737), .IN4(n5738), .QN(
        s5_data_o[7]) );
  OA22X1 U28998 ( .IN1(n1734), .IN2(n20301), .IN3(n1629), .IN4(n20289), .Q(
        n5735) );
  OA22X1 U28999 ( .IN1(n1906), .IN2(n20328), .IN3(n1820), .IN4(n20320), .Q(
        n5736) );
  OA22X1 U29000 ( .IN1(n2078), .IN2(n20361), .IN3(n1992), .IN4(n20353), .Q(
        n5737) );
  NAND4X0 U29001 ( .IN1(n5731), .IN2(n5732), .IN3(n5733), .IN4(n5734), .QN(
        s5_data_o[8]) );
  OA22X1 U29002 ( .IN1(n1733), .IN2(n20301), .IN3(n1628), .IN4(n20289), .Q(
        n5731) );
  OA22X1 U29003 ( .IN1(n1905), .IN2(n20335), .IN3(n1819), .IN4(n20320), .Q(
        n5732) );
  OA22X1 U29004 ( .IN1(n2077), .IN2(n20368), .IN3(n1991), .IN4(n20353), .Q(
        n5733) );
  NAND4X0 U29005 ( .IN1(n5727), .IN2(n5728), .IN3(n5729), .IN4(n5730), .QN(
        s5_data_o[9]) );
  OA22X1 U29006 ( .IN1(n1732), .IN2(n20301), .IN3(n1627), .IN4(n20288), .Q(
        n5727) );
  OA22X1 U29007 ( .IN1(n1904), .IN2(n20328), .IN3(n1818), .IN4(n20321), .Q(
        n5728) );
  OA22X1 U29008 ( .IN1(n2076), .IN2(n20361), .IN3(n1990), .IN4(n20354), .Q(
        n5729) );
  NAND4X0 U29009 ( .IN1(n5847), .IN2(n5848), .IN3(n5849), .IN4(n5850), .QN(
        s5_data_o[10]) );
  OA22X1 U29010 ( .IN1(n1731), .IN2(n20296), .IN3(n1626), .IN4(n20282), .Q(
        n5847) );
  OA22X1 U29011 ( .IN1(n1903), .IN2(n20330), .IN3(n1817), .IN4(n20315), .Q(
        n5848) );
  OA22X1 U29012 ( .IN1(n2075), .IN2(n20363), .IN3(n1989), .IN4(n20348), .Q(
        n5849) );
  NAND4X0 U29013 ( .IN1(n5843), .IN2(n5844), .IN3(n5845), .IN4(n5846), .QN(
        s5_data_o[11]) );
  OA22X1 U29014 ( .IN1(n1730), .IN2(n20297), .IN3(n1625), .IN4(n20282), .Q(
        n5843) );
  OA22X1 U29015 ( .IN1(n1902), .IN2(n20335), .IN3(n1816), .IN4(n20315), .Q(
        n5844) );
  OA22X1 U29016 ( .IN1(n2074), .IN2(n20368), .IN3(n1988), .IN4(n20348), .Q(
        n5845) );
  NAND4X0 U29017 ( .IN1(n5839), .IN2(n5840), .IN3(n5841), .IN4(n5842), .QN(
        s5_data_o[12]) );
  OA22X1 U29018 ( .IN1(n1729), .IN2(n20298), .IN3(n1624), .IN4(n20282), .Q(
        n5839) );
  OA22X1 U29019 ( .IN1(n1901), .IN2(n20331), .IN3(n1815), .IN4(n20315), .Q(
        n5840) );
  OA22X1 U29020 ( .IN1(n2073), .IN2(n20364), .IN3(n1987), .IN4(n20348), .Q(
        n5841) );
  NAND4X0 U29021 ( .IN1(n5835), .IN2(n5836), .IN3(n5837), .IN4(n5838), .QN(
        s5_data_o[13]) );
  OA22X1 U29022 ( .IN1(n1728), .IN2(n20299), .IN3(n1623), .IN4(n20283), .Q(
        n5835) );
  OA22X1 U29023 ( .IN1(n1900), .IN2(n20332), .IN3(n1814), .IN4(n20309), .Q(
        n5836) );
  OA22X1 U29024 ( .IN1(n2072), .IN2(n20365), .IN3(n1986), .IN4(n20342), .Q(
        n5837) );
  NAND4X0 U29025 ( .IN1(n5831), .IN2(n5832), .IN3(n5833), .IN4(n5834), .QN(
        s5_data_o[14]) );
  OA22X1 U29026 ( .IN1(n1727), .IN2(n20299), .IN3(n1622), .IN4(n20283), .Q(
        n5831) );
  OA22X1 U29027 ( .IN1(n1899), .IN2(n20332), .IN3(n1813), .IN4(n20314), .Q(
        n5832) );
  OA22X1 U29028 ( .IN1(n2071), .IN2(n20365), .IN3(n1985), .IN4(n20347), .Q(
        n5833) );
  NAND4X0 U29029 ( .IN1(n5827), .IN2(n5828), .IN3(n5829), .IN4(n5830), .QN(
        s5_data_o[15]) );
  OA22X1 U29030 ( .IN1(n1726), .IN2(n20299), .IN3(n1621), .IN4(n20283), .Q(
        n5827) );
  OA22X1 U29031 ( .IN1(n1898), .IN2(n20332), .IN3(n1812), .IN4(n20315), .Q(
        n5828) );
  OA22X1 U29032 ( .IN1(n2070), .IN2(n20365), .IN3(n1984), .IN4(n20348), .Q(
        n5829) );
  NAND4X0 U29033 ( .IN1(n5823), .IN2(n5824), .IN3(n5825), .IN4(n5826), .QN(
        s5_data_o[16]) );
  OA22X1 U29034 ( .IN1(n1725), .IN2(n20299), .IN3(n1620), .IN4(n20284), .Q(
        n5823) );
  OA22X1 U29035 ( .IN1(n1897), .IN2(n20332), .IN3(n1811), .IN4(n20316), .Q(
        n5824) );
  OA22X1 U29036 ( .IN1(n2069), .IN2(n20365), .IN3(n1983), .IN4(n20349), .Q(
        n5825) );
  NAND4X0 U29037 ( .IN1(n5819), .IN2(n5820), .IN3(n5821), .IN4(n5822), .QN(
        s5_data_o[17]) );
  OA22X1 U29038 ( .IN1(n1724), .IN2(n20302), .IN3(n1619), .IN4(n20284), .Q(
        n5819) );
  OA22X1 U29039 ( .IN1(n1896), .IN2(n20333), .IN3(n1810), .IN4(n20316), .Q(
        n5820) );
  OA22X1 U29040 ( .IN1(n2068), .IN2(n20366), .IN3(n1982), .IN4(n20349), .Q(
        n5821) );
  NAND4X0 U29041 ( .IN1(n5815), .IN2(n5816), .IN3(n5817), .IN4(n5818), .QN(
        s5_data_o[18]) );
  OA22X1 U29042 ( .IN1(n1723), .IN2(n20302), .IN3(n1618), .IN4(n20284), .Q(
        n5815) );
  OA22X1 U29043 ( .IN1(n1895), .IN2(n20333), .IN3(n1809), .IN4(n20316), .Q(
        n5816) );
  OA22X1 U29044 ( .IN1(n2067), .IN2(n20366), .IN3(n1981), .IN4(n20349), .Q(
        n5817) );
  NAND4X0 U29045 ( .IN1(n5811), .IN2(n5812), .IN3(n5813), .IN4(n5814), .QN(
        s5_data_o[19]) );
  OA22X1 U29046 ( .IN1(n1722), .IN2(n20297), .IN3(n1617), .IN4(n20284), .Q(
        n5811) );
  OA22X1 U29047 ( .IN1(n1894), .IN2(n20333), .IN3(n1808), .IN4(n20316), .Q(
        n5812) );
  OA22X1 U29048 ( .IN1(n2066), .IN2(n20366), .IN3(n1980), .IN4(n20349), .Q(
        n5813) );
  NAND4X0 U29049 ( .IN1(n5803), .IN2(n5804), .IN3(n5805), .IN4(n5806), .QN(
        s5_data_o[20]) );
  OA22X1 U29050 ( .IN1(n1721), .IN2(n20300), .IN3(n1616), .IN4(n20283), .Q(
        n5803) );
  OA22X1 U29051 ( .IN1(n1893), .IN2(n20334), .IN3(n1807), .IN4(n20313), .Q(
        n5804) );
  OA22X1 U29052 ( .IN1(n2065), .IN2(n20367), .IN3(n1979), .IN4(n20346), .Q(
        n5805) );
  NAND4X0 U29053 ( .IN1(n5799), .IN2(n5800), .IN3(n5801), .IN4(n5802), .QN(
        s5_data_o[21]) );
  OA22X1 U29054 ( .IN1(n1720), .IN2(n20300), .IN3(n1615), .IN4(n20285), .Q(
        n5799) );
  OA22X1 U29055 ( .IN1(n1892), .IN2(n20334), .IN3(n1806), .IN4(n20317), .Q(
        n5800) );
  OA22X1 U29056 ( .IN1(n2064), .IN2(n20367), .IN3(n1978), .IN4(n20350), .Q(
        n5801) );
  NAND4X0 U29057 ( .IN1(n5795), .IN2(n5796), .IN3(n5797), .IN4(n5798), .QN(
        s5_data_o[22]) );
  OA22X1 U29058 ( .IN1(n1719), .IN2(n20299), .IN3(n1614), .IN4(n20285), .Q(
        n5795) );
  OA22X1 U29059 ( .IN1(n1891), .IN2(n20332), .IN3(n1805), .IN4(n20317), .Q(
        n5796) );
  OA22X1 U29060 ( .IN1(n2063), .IN2(n20365), .IN3(n1977), .IN4(n20350), .Q(
        n5797) );
  NAND4X0 U29061 ( .IN1(n5791), .IN2(n5792), .IN3(n5793), .IN4(n5794), .QN(
        s5_data_o[23]) );
  OA22X1 U29062 ( .IN1(n1718), .IN2(n20298), .IN3(n1613), .IN4(n20285), .Q(
        n5791) );
  OA22X1 U29063 ( .IN1(n1890), .IN2(n20333), .IN3(n1804), .IN4(n20317), .Q(
        n5792) );
  OA22X1 U29064 ( .IN1(n2062), .IN2(n20366), .IN3(n1976), .IN4(n20350), .Q(
        n5793) );
  NAND4X0 U29065 ( .IN1(n5787), .IN2(n5788), .IN3(n5789), .IN4(n5790), .QN(
        s5_data_o[24]) );
  OA22X1 U29066 ( .IN1(n1717), .IN2(n20301), .IN3(n1612), .IN4(n20286), .Q(
        n5787) );
  OA22X1 U29067 ( .IN1(n1889), .IN2(n20331), .IN3(n1803), .IN4(n20318), .Q(
        n5788) );
  OA22X1 U29068 ( .IN1(n2061), .IN2(n20364), .IN3(n1975), .IN4(n20351), .Q(
        n5789) );
  NAND4X0 U29069 ( .IN1(n5783), .IN2(n5784), .IN3(n5785), .IN4(n5786), .QN(
        s5_data_o[25]) );
  OA22X1 U29070 ( .IN1(n1716), .IN2(n20298), .IN3(n1611), .IN4(n20286), .Q(
        n5783) );
  OA22X1 U29071 ( .IN1(n1888), .IN2(n20331), .IN3(n1802), .IN4(n20318), .Q(
        n5784) );
  OA22X1 U29072 ( .IN1(n2060), .IN2(n20364), .IN3(n1974), .IN4(n20351), .Q(
        n5785) );
  NAND4X0 U29073 ( .IN1(n5779), .IN2(n5780), .IN3(n5781), .IN4(n5782), .QN(
        s5_data_o[26]) );
  OA22X1 U29074 ( .IN1(n1715), .IN2(n20296), .IN3(n1610), .IN4(n20286), .Q(
        n5779) );
  OA22X1 U29075 ( .IN1(n1887), .IN2(n20330), .IN3(n1801), .IN4(n20318), .Q(
        n5780) );
  OA22X1 U29076 ( .IN1(n2059), .IN2(n20363), .IN3(n1973), .IN4(n20351), .Q(
        n5781) );
  NAND4X0 U29077 ( .IN1(n5775), .IN2(n5776), .IN3(n5777), .IN4(n5778), .QN(
        s5_data_o[27]) );
  OA22X1 U29078 ( .IN1(n1714), .IN2(n20301), .IN3(n1609), .IN4(n20285), .Q(
        n5775) );
  OA22X1 U29079 ( .IN1(n1886), .IN2(n20333), .IN3(n1800), .IN4(n20319), .Q(
        n5776) );
  OA22X1 U29080 ( .IN1(n2058), .IN2(n20366), .IN3(n1972), .IN4(n20352), .Q(
        n5777) );
  NAND4X0 U29081 ( .IN1(n5771), .IN2(n5772), .IN3(n5773), .IN4(n5774), .QN(
        s5_data_o[28]) );
  OA22X1 U29082 ( .IN1(n1713), .IN2(n20300), .IN3(n1608), .IN4(n20286), .Q(
        n5771) );
  OA22X1 U29083 ( .IN1(n1885), .IN2(n20334), .IN3(n1799), .IN4(n20319), .Q(
        n5772) );
  OA22X1 U29084 ( .IN1(n2057), .IN2(n20367), .IN3(n1971), .IN4(n20352), .Q(
        n5773) );
  NAND4X0 U29085 ( .IN1(n5767), .IN2(n5768), .IN3(n5769), .IN4(n5770), .QN(
        s5_data_o[29]) );
  OA22X1 U29086 ( .IN1(n1712), .IN2(n20300), .IN3(n1607), .IN4(n20285), .Q(
        n5767) );
  OA22X1 U29087 ( .IN1(n1884), .IN2(n20334), .IN3(n1798), .IN4(n20319), .Q(
        n5768) );
  OA22X1 U29088 ( .IN1(n2056), .IN2(n20367), .IN3(n1970), .IN4(n20352), .Q(
        n5769) );
  NAND4X0 U29089 ( .IN1(n5759), .IN2(n5760), .IN3(n5761), .IN4(n5762), .QN(
        s5_data_o[30]) );
  OA22X1 U29090 ( .IN1(n1711), .IN2(n20300), .IN3(n1606), .IN4(n20288), .Q(
        n5759) );
  OA22X1 U29091 ( .IN1(n1883), .IN2(n20334), .IN3(n1797), .IN4(n20321), .Q(
        n5760) );
  OA22X1 U29092 ( .IN1(n2055), .IN2(n20367), .IN3(n1969), .IN4(n20354), .Q(
        n5761) );
  NAND4X0 U29093 ( .IN1(n5755), .IN2(n5756), .IN3(n5757), .IN4(n5758), .QN(
        s5_data_o[31]) );
  OA22X1 U29094 ( .IN1(n1710), .IN2(n20299), .IN3(n1605), .IN4(n20287), .Q(
        n5755) );
  OA22X1 U29095 ( .IN1(n1882), .IN2(n20332), .IN3(n1796), .IN4(n20306), .Q(
        n5756) );
  OA22X1 U29096 ( .IN1(n2054), .IN2(n20365), .IN3(n1968), .IN4(n20339), .Q(
        n5757) );
  NAND4X0 U29097 ( .IN1(n5995), .IN2(n5996), .IN3(n5997), .IN4(n5998), .QN(
        s4_stb_o) );
  OA22X1 U29098 ( .IN1(n1795), .IN2(n6005), .IN3(n1709), .IN4(n6006), .Q(n5995) );
  OA22X1 U29099 ( .IN1(n1967), .IN2(n6003), .IN3(n1881), .IN4(n6004), .Q(n5996) );
  OA22X1 U29100 ( .IN1(n2139), .IN2(n6001), .IN3(n2053), .IN4(n6002), .Q(n5997) );
  NAND4X0 U29101 ( .IN1(n5983), .IN2(n5984), .IN3(n5985), .IN4(n5986), .QN(
        s4_we_o) );
  OA22X1 U29102 ( .IN1(n1794), .IN2(n20163), .IN3(n1708), .IN4(n20157), .Q(
        n5983) );
  OA22X1 U29103 ( .IN1(n1966), .IN2(n20196), .IN3(n1880), .IN4(n20190), .Q(
        n5984) );
  OA22X1 U29104 ( .IN1(n2138), .IN2(n20229), .IN3(n2052), .IN4(n20223), .Q(
        n5985) );
  NAND4X0 U29105 ( .IN1(n6019), .IN2(n6020), .IN3(n6021), .IN4(n6022), .QN(
        s4_sel_o[0]) );
  OA22X1 U29106 ( .IN1(n1793), .IN2(n20170), .IN3(n1707), .IN4(n20156), .Q(
        n6019) );
  OA22X1 U29107 ( .IN1(n1965), .IN2(n20203), .IN3(n1879), .IN4(n20189), .Q(
        n6020) );
  OA22X1 U29108 ( .IN1(n2137), .IN2(n20236), .IN3(n2051), .IN4(n20222), .Q(
        n6021) );
  NAND4X0 U29109 ( .IN1(n6015), .IN2(n6016), .IN3(n6017), .IN4(n6018), .QN(
        s4_sel_o[1]) );
  OA22X1 U29110 ( .IN1(n1792), .IN2(n20170), .IN3(n1706), .IN4(n20156), .Q(
        n6015) );
  OA22X1 U29111 ( .IN1(n1964), .IN2(n20203), .IN3(n1878), .IN4(n20189), .Q(
        n6016) );
  OA22X1 U29112 ( .IN1(n2136), .IN2(n20236), .IN3(n2050), .IN4(n20222), .Q(
        n6017) );
  NAND4X0 U29113 ( .IN1(n6011), .IN2(n6012), .IN3(n6013), .IN4(n6014), .QN(
        s4_sel_o[2]) );
  OA22X1 U29114 ( .IN1(n1791), .IN2(n20170), .IN3(n1705), .IN4(n20157), .Q(
        n6011) );
  OA22X1 U29115 ( .IN1(n1963), .IN2(n20203), .IN3(n1877), .IN4(n20190), .Q(
        n6012) );
  OA22X1 U29116 ( .IN1(n2135), .IN2(n20236), .IN3(n2049), .IN4(n20223), .Q(
        n6013) );
  NAND4X0 U29117 ( .IN1(n6007), .IN2(n6008), .IN3(n6009), .IN4(n6010), .QN(
        s4_sel_o[3]) );
  OA22X1 U29118 ( .IN1(n1790), .IN2(n20170), .IN3(n1704), .IN4(n20157), .Q(
        n6007) );
  OA22X1 U29119 ( .IN1(n1962), .IN2(n20203), .IN3(n1876), .IN4(n20190), .Q(
        n6008) );
  OA22X1 U29120 ( .IN1(n2134), .IN2(n20236), .IN3(n2048), .IN4(n20223), .Q(
        n6009) );
  NAND4X0 U29121 ( .IN1(n6275), .IN2(n6276), .IN3(n6277), .IN4(n6278), .QN(
        s4_addr_o[0]) );
  OA22X1 U29122 ( .IN1(n1789), .IN2(n20163), .IN3(n1703), .IN4(n20140), .Q(
        n6275) );
  OA22X1 U29123 ( .IN1(n1961), .IN2(n20196), .IN3(n1875), .IN4(n20173), .Q(
        n6276) );
  OA22X1 U29124 ( .IN1(n2133), .IN2(n20229), .IN3(n2047), .IN4(n20206), .Q(
        n6277) );
  NAND4X0 U29125 ( .IN1(n6231), .IN2(n6232), .IN3(n6233), .IN4(n6234), .QN(
        s4_addr_o[1]) );
  OA22X1 U29126 ( .IN1(n1788), .IN2(n20165), .IN3(n1702), .IN4(n20143), .Q(
        n6231) );
  OA22X1 U29127 ( .IN1(n1960), .IN2(n20198), .IN3(n1874), .IN4(n20176), .Q(
        n6232) );
  OA22X1 U29128 ( .IN1(n2132), .IN2(n20231), .IN3(n2046), .IN4(n20209), .Q(
        n6233) );
  NAND4X0 U29129 ( .IN1(n6187), .IN2(n6188), .IN3(n6189), .IN4(n6190), .QN(
        s4_addr_o[2]) );
  OA22X1 U29130 ( .IN1(n1787), .IN2(n20165), .IN3(n1701), .IN4(n20147), .Q(
        n6187) );
  OA22X1 U29131 ( .IN1(n1959), .IN2(n20198), .IN3(n1873), .IN4(n20180), .Q(
        n6188) );
  OA22X1 U29132 ( .IN1(n2131), .IN2(n20231), .IN3(n2045), .IN4(n20213), .Q(
        n6189) );
  NAND4X0 U29133 ( .IN1(n6175), .IN2(n6176), .IN3(n6177), .IN4(n6178), .QN(
        s4_addr_o[3]) );
  OA22X1 U29134 ( .IN1(n1786), .IN2(n20170), .IN3(n1699), .IN4(n20148), .Q(
        n6175) );
  OA22X1 U29135 ( .IN1(n1958), .IN2(n20203), .IN3(n1872), .IN4(n20181), .Q(
        n6176) );
  OA22X1 U29136 ( .IN1(n2130), .IN2(n20236), .IN3(n2044), .IN4(n20214), .Q(
        n6177) );
  NAND4X0 U29137 ( .IN1(n6171), .IN2(n6172), .IN3(n6173), .IN4(n6174), .QN(
        s4_addr_o[4]) );
  OA22X1 U29138 ( .IN1(n1785), .IN2(n20163), .IN3(n1697), .IN4(n20148), .Q(
        n6171) );
  OA22X1 U29139 ( .IN1(n1957), .IN2(n20196), .IN3(n1871), .IN4(n20181), .Q(
        n6172) );
  OA22X1 U29140 ( .IN1(n2129), .IN2(n20229), .IN3(n2043), .IN4(n20214), .Q(
        n6173) );
  NAND4X0 U29141 ( .IN1(n6167), .IN2(n6168), .IN3(n6169), .IN4(n6170), .QN(
        s4_addr_o[5]) );
  OA22X1 U29142 ( .IN1(n1784), .IN2(n20170), .IN3(n1696), .IN4(n20147), .Q(
        n6167) );
  OA22X1 U29143 ( .IN1(n1956), .IN2(n20203), .IN3(n1870), .IN4(n20180), .Q(
        n6168) );
  OA22X1 U29144 ( .IN1(n2128), .IN2(n20236), .IN3(n2042), .IN4(n20213), .Q(
        n6169) );
  NAND4X0 U29145 ( .IN1(n6163), .IN2(n6164), .IN3(n6165), .IN4(n6166), .QN(
        s4_addr_o[6]) );
  OA22X1 U29146 ( .IN1(n1783), .IN2(n20166), .IN3(n1679), .IN4(n20148), .Q(
        n6163) );
  OA22X1 U29147 ( .IN1(n1955), .IN2(n20199), .IN3(n1869), .IN4(n20181), .Q(
        n6164) );
  OA22X1 U29148 ( .IN1(n2127), .IN2(n20232), .IN3(n2041), .IN4(n20214), .Q(
        n6165) );
  NAND4X0 U29149 ( .IN1(n6159), .IN2(n6160), .IN3(n6161), .IN4(n6162), .QN(
        s4_addr_o[7]) );
  OA22X1 U29150 ( .IN1(n1782), .IN2(n20166), .IN3(n1678), .IN4(n20140), .Q(
        n6159) );
  OA22X1 U29151 ( .IN1(n1954), .IN2(n20199), .IN3(n1868), .IN4(n20173), .Q(
        n6160) );
  OA22X1 U29152 ( .IN1(n2126), .IN2(n20232), .IN3(n2040), .IN4(n20213), .Q(
        n6161) );
  NAND4X0 U29153 ( .IN1(n6155), .IN2(n6156), .IN3(n6157), .IN4(n6158), .QN(
        s4_addr_o[8]) );
  OA22X1 U29154 ( .IN1(n1781), .IN2(n20166), .IN3(n1677), .IN4(n20149), .Q(
        n6155) );
  OA22X1 U29155 ( .IN1(n1953), .IN2(n20199), .IN3(n1867), .IN4(n20182), .Q(
        n6156) );
  OA22X1 U29156 ( .IN1(n2125), .IN2(n20232), .IN3(n2039), .IN4(n20215), .Q(
        n6157) );
  NAND4X0 U29157 ( .IN1(n6151), .IN2(n6152), .IN3(n6153), .IN4(n6154), .QN(
        s4_addr_o[9]) );
  OA22X1 U29158 ( .IN1(n1780), .IN2(n20166), .IN3(n1676), .IN4(n20149), .Q(
        n6151) );
  OA22X1 U29159 ( .IN1(n1952), .IN2(n20199), .IN3(n1866), .IN4(n20182), .Q(
        n6152) );
  OA22X1 U29160 ( .IN1(n2124), .IN2(n20232), .IN3(n2038), .IN4(n20215), .Q(
        n6153) );
  NAND4X0 U29161 ( .IN1(n6271), .IN2(n6272), .IN3(n6273), .IN4(n6274), .QN(
        s4_addr_o[10]) );
  OA22X1 U29162 ( .IN1(n1779), .IN2(n20163), .IN3(n1675), .IN4(n20140), .Q(
        n6271) );
  OA22X1 U29163 ( .IN1(n1951), .IN2(n20196), .IN3(n1865), .IN4(n20173), .Q(
        n6272) );
  OA22X1 U29164 ( .IN1(n2123), .IN2(n20229), .IN3(n2037), .IN4(n20206), .Q(
        n6273) );
  NAND4X0 U29165 ( .IN1(n6267), .IN2(n6268), .IN3(n6269), .IN4(n6270), .QN(
        s4_addr_o[11]) );
  OA22X1 U29166 ( .IN1(n1778), .IN2(n20163), .IN3(n1674), .IN4(n20140), .Q(
        n6267) );
  OA22X1 U29167 ( .IN1(n1950), .IN2(n20196), .IN3(n1864), .IN4(n20173), .Q(
        n6268) );
  OA22X1 U29168 ( .IN1(n2122), .IN2(n20229), .IN3(n2036), .IN4(n20206), .Q(
        n6269) );
  NAND4X0 U29169 ( .IN1(n6263), .IN2(n6264), .IN3(n6265), .IN4(n6266), .QN(
        s4_addr_o[12]) );
  OA22X1 U29170 ( .IN1(n1777), .IN2(n20163), .IN3(n1673), .IN4(n20141), .Q(
        n6263) );
  OA22X1 U29171 ( .IN1(n1949), .IN2(n20196), .IN3(n1863), .IN4(n20174), .Q(
        n6264) );
  OA22X1 U29172 ( .IN1(n2121), .IN2(n20229), .IN3(n2035), .IN4(n20207), .Q(
        n6265) );
  NAND4X0 U29173 ( .IN1(n6259), .IN2(n6260), .IN3(n6261), .IN4(n6262), .QN(
        s4_addr_o[13]) );
  OA22X1 U29174 ( .IN1(n1776), .IN2(n20164), .IN3(n1672), .IN4(n20141), .Q(
        n6259) );
  OA22X1 U29175 ( .IN1(n1948), .IN2(n20197), .IN3(n1862), .IN4(n20174), .Q(
        n6260) );
  OA22X1 U29176 ( .IN1(n2120), .IN2(n20230), .IN3(n2034), .IN4(n20207), .Q(
        n6261) );
  NAND4X0 U29177 ( .IN1(n6255), .IN2(n6256), .IN3(n6257), .IN4(n6258), .QN(
        s4_addr_o[14]) );
  OA22X1 U29178 ( .IN1(n1775), .IN2(n20164), .IN3(n1671), .IN4(n20141), .Q(
        n6255) );
  OA22X1 U29179 ( .IN1(n1947), .IN2(n20197), .IN3(n1861), .IN4(n20174), .Q(
        n6256) );
  OA22X1 U29180 ( .IN1(n2119), .IN2(n20230), .IN3(n2033), .IN4(n20207), .Q(
        n6257) );
  NAND4X0 U29181 ( .IN1(n6251), .IN2(n6252), .IN3(n6253), .IN4(n6254), .QN(
        s4_addr_o[15]) );
  OA22X1 U29182 ( .IN1(n1774), .IN2(n20164), .IN3(n1670), .IN4(n20142), .Q(
        n6251) );
  OA22X1 U29183 ( .IN1(n1946), .IN2(n20197), .IN3(n1860), .IN4(n20175), .Q(
        n6252) );
  OA22X1 U29184 ( .IN1(n2118), .IN2(n20230), .IN3(n2032), .IN4(n20208), .Q(
        n6253) );
  NAND4X0 U29185 ( .IN1(n6247), .IN2(n6248), .IN3(n6249), .IN4(n6250), .QN(
        s4_addr_o[16]) );
  OA22X1 U29186 ( .IN1(n1773), .IN2(n20164), .IN3(n1669), .IN4(n20142), .Q(
        n6247) );
  OA22X1 U29187 ( .IN1(n1945), .IN2(n20197), .IN3(n1859), .IN4(n20175), .Q(
        n6248) );
  OA22X1 U29188 ( .IN1(n2117), .IN2(n20230), .IN3(n2031), .IN4(n20208), .Q(
        n6249) );
  NAND4X0 U29189 ( .IN1(n6243), .IN2(n6244), .IN3(n6245), .IN4(n6246), .QN(
        s4_addr_o[17]) );
  OA22X1 U29190 ( .IN1(n1772), .IN2(n20165), .IN3(n1668), .IN4(n20142), .Q(
        n6243) );
  OA22X1 U29191 ( .IN1(n1944), .IN2(n20198), .IN3(n1858), .IN4(n20175), .Q(
        n6244) );
  OA22X1 U29192 ( .IN1(n2116), .IN2(n20231), .IN3(n2030), .IN4(n20208), .Q(
        n6245) );
  NAND4X0 U29193 ( .IN1(n6239), .IN2(n6240), .IN3(n6241), .IN4(n6242), .QN(
        s4_addr_o[18]) );
  OA22X1 U29194 ( .IN1(n1771), .IN2(n20165), .IN3(n1667), .IN4(n20143), .Q(
        n6239) );
  OA22X1 U29195 ( .IN1(n1943), .IN2(n20198), .IN3(n1857), .IN4(n20176), .Q(
        n6240) );
  OA22X1 U29196 ( .IN1(n2115), .IN2(n20231), .IN3(n2029), .IN4(n20209), .Q(
        n6241) );
  NAND4X0 U29197 ( .IN1(n6235), .IN2(n6236), .IN3(n6237), .IN4(n6238), .QN(
        s4_addr_o[19]) );
  OA22X1 U29198 ( .IN1(n1770), .IN2(n20165), .IN3(n1666), .IN4(n20143), .Q(
        n6235) );
  OA22X1 U29199 ( .IN1(n1942), .IN2(n20198), .IN3(n1856), .IN4(n20176), .Q(
        n6236) );
  OA22X1 U29200 ( .IN1(n2114), .IN2(n20231), .IN3(n2028), .IN4(n20209), .Q(
        n6237) );
  NAND4X0 U29201 ( .IN1(n6227), .IN2(n6228), .IN3(n6229), .IN4(n6230), .QN(
        s4_addr_o[20]) );
  OA22X1 U29202 ( .IN1(n1769), .IN2(n20164), .IN3(n1665), .IN4(n20144), .Q(
        n6227) );
  OA22X1 U29203 ( .IN1(n1941), .IN2(n20197), .IN3(n1855), .IN4(n20177), .Q(
        n6228) );
  OA22X1 U29204 ( .IN1(n2113), .IN2(n20230), .IN3(n2027), .IN4(n20210), .Q(
        n6229) );
  NAND4X0 U29205 ( .IN1(n6223), .IN2(n6224), .IN3(n6225), .IN4(n6226), .QN(
        s4_addr_o[21]) );
  OA22X1 U29206 ( .IN1(n1768), .IN2(n20164), .IN3(n1664), .IN4(n20144), .Q(
        n6223) );
  OA22X1 U29207 ( .IN1(n1940), .IN2(n20197), .IN3(n1854), .IN4(n20177), .Q(
        n6224) );
  OA22X1 U29208 ( .IN1(n2112), .IN2(n20230), .IN3(n2026), .IN4(n20210), .Q(
        n6225) );
  NAND4X0 U29209 ( .IN1(n6219), .IN2(n6220), .IN3(n6221), .IN4(n6222), .QN(
        s4_addr_o[22]) );
  OA22X1 U29210 ( .IN1(n1767), .IN2(n20163), .IN3(n1663), .IN4(n20144), .Q(
        n6219) );
  OA22X1 U29211 ( .IN1(n1939), .IN2(n20196), .IN3(n1853), .IN4(n20177), .Q(
        n6220) );
  OA22X1 U29212 ( .IN1(n2111), .IN2(n20229), .IN3(n2025), .IN4(n20210), .Q(
        n6221) );
  NAND4X0 U29213 ( .IN1(n6215), .IN2(n6216), .IN3(n6217), .IN4(n6218), .QN(
        s4_addr_o[23]) );
  OA22X1 U29214 ( .IN1(n1766), .IN2(n20164), .IN3(n1662), .IN4(n20145), .Q(
        n6215) );
  OA22X1 U29215 ( .IN1(n1938), .IN2(n20197), .IN3(n1852), .IN4(n20178), .Q(
        n6216) );
  OA22X1 U29216 ( .IN1(n2110), .IN2(n20230), .IN3(n2024), .IN4(n20211), .Q(
        n6217) );
  NAND4X0 U29217 ( .IN1(n6211), .IN2(n6212), .IN3(n6213), .IN4(n6214), .QN(
        s4_addr_o[24]) );
  OA22X1 U29218 ( .IN1(n1765), .IN2(n20170), .IN3(n1661), .IN4(n20145), .Q(
        n6211) );
  OA22X1 U29219 ( .IN1(n1937), .IN2(n20203), .IN3(n1851), .IN4(n20178), .Q(
        n6212) );
  OA22X1 U29220 ( .IN1(n2109), .IN2(n20236), .IN3(n2023), .IN4(n20211), .Q(
        n6213) );
  NAND4X0 U29221 ( .IN1(n6207), .IN2(n6208), .IN3(n6209), .IN4(n6210), .QN(
        s4_addr_o[25]) );
  OA22X1 U29222 ( .IN1(n1764), .IN2(n20166), .IN3(n1660), .IN4(n20145), .Q(
        n6207) );
  OA22X1 U29223 ( .IN1(n1936), .IN2(n20199), .IN3(n1850), .IN4(n20178), .Q(
        n6208) );
  OA22X1 U29224 ( .IN1(n2108), .IN2(n20232), .IN3(n2022), .IN4(n20211), .Q(
        n6209) );
  NAND4X0 U29225 ( .IN1(n6203), .IN2(n6204), .IN3(n6205), .IN4(n6206), .QN(
        s4_addr_o[26]) );
  OA22X1 U29226 ( .IN1(n1763), .IN2(n20165), .IN3(n1659), .IN4(n20146), .Q(
        n6203) );
  OA22X1 U29227 ( .IN1(n1935), .IN2(n20198), .IN3(n1849), .IN4(n20179), .Q(
        n6204) );
  OA22X1 U29228 ( .IN1(n2107), .IN2(n20231), .IN3(n2021), .IN4(n20212), .Q(
        n6205) );
  NAND4X0 U29229 ( .IN1(n6199), .IN2(n6200), .IN3(n6201), .IN4(n6202), .QN(
        s4_addr_o[27]) );
  OA22X1 U29230 ( .IN1(n1762), .IN2(n20164), .IN3(n1658), .IN4(n20146), .Q(
        n6199) );
  OA22X1 U29231 ( .IN1(n1934), .IN2(n20197), .IN3(n1848), .IN4(n20179), .Q(
        n6200) );
  OA22X1 U29232 ( .IN1(n2106), .IN2(n20230), .IN3(n2020), .IN4(n20212), .Q(
        n6201) );
  NAND4X0 U29233 ( .IN1(n6195), .IN2(n6196), .IN3(n6197), .IN4(n6198), .QN(
        s4_addr_o[28]) );
  OA22X1 U29234 ( .IN1(n1761), .IN2(n20164), .IN3(n1657), .IN4(n20146), .Q(
        n6195) );
  OA22X1 U29235 ( .IN1(n1933), .IN2(n20197), .IN3(n1847), .IN4(n20179), .Q(
        n6196) );
  OA22X1 U29236 ( .IN1(n2105), .IN2(n20230), .IN3(n2019), .IN4(n20212), .Q(
        n6197) );
  NAND4X0 U29237 ( .IN1(n6191), .IN2(n6192), .IN3(n6193), .IN4(n6194), .QN(
        s4_addr_o[29]) );
  OA22X1 U29238 ( .IN1(n1760), .IN2(n20168), .IN3(n1656), .IN4(n20147), .Q(
        n6191) );
  OA22X1 U29239 ( .IN1(n1932), .IN2(n20201), .IN3(n1846), .IN4(n20180), .Q(
        n6192) );
  OA22X1 U29240 ( .IN1(n2104), .IN2(n20234), .IN3(n2018), .IN4(n20213), .Q(
        n6193) );
  NAND4X0 U29241 ( .IN1(n6183), .IN2(n6184), .IN3(n6185), .IN4(n6186), .QN(
        s4_addr_o[30]) );
  OA22X1 U29242 ( .IN1(n1759), .IN2(n20169), .IN3(n1655), .IN4(n20147), .Q(
        n6183) );
  OA22X1 U29243 ( .IN1(n1931), .IN2(n20202), .IN3(n1845), .IN4(n20180), .Q(
        n6184) );
  OA22X1 U29244 ( .IN1(n2103), .IN2(n20235), .IN3(n2017), .IN4(n20213), .Q(
        n6185) );
  NAND4X0 U29245 ( .IN1(n6179), .IN2(n6180), .IN3(n6181), .IN4(n6182), .QN(
        s4_addr_o[31]) );
  OA22X1 U29246 ( .IN1(n1758), .IN2(n20167), .IN3(n1650), .IN4(n20148), .Q(
        n6179) );
  OA22X1 U29247 ( .IN1(n1930), .IN2(n20200), .IN3(n1844), .IN4(n20181), .Q(
        n6180) );
  OA22X1 U29248 ( .IN1(n2102), .IN2(n20233), .IN3(n2016), .IN4(n20214), .Q(
        n6181) );
  NAND4X0 U29249 ( .IN1(n6147), .IN2(n6148), .IN3(n6149), .IN4(n6150), .QN(
        s4_data_o[0]) );
  OA22X1 U29250 ( .IN1(n1741), .IN2(n20166), .IN3(n1636), .IN4(n20149), .Q(
        n6147) );
  OA22X1 U29251 ( .IN1(n1913), .IN2(n20199), .IN3(n1827), .IN4(n20182), .Q(
        n6148) );
  OA22X1 U29252 ( .IN1(n2085), .IN2(n20232), .IN3(n1999), .IN4(n20215), .Q(
        n6149) );
  NAND4X0 U29253 ( .IN1(n6103), .IN2(n6104), .IN3(n6105), .IN4(n6106), .QN(
        s4_data_o[1]) );
  OA22X1 U29254 ( .IN1(n1740), .IN2(n20168), .IN3(n1635), .IN4(n20147), .Q(
        n6103) );
  OA22X1 U29255 ( .IN1(n1912), .IN2(n20201), .IN3(n1826), .IN4(n20180), .Q(
        n6104) );
  OA22X1 U29256 ( .IN1(n2084), .IN2(n20234), .IN3(n1998), .IN4(n20213), .Q(
        n6105) );
  NAND4X0 U29257 ( .IN1(n6059), .IN2(n6060), .IN3(n6061), .IN4(n6062), .QN(
        s4_data_o[2]) );
  OA22X1 U29258 ( .IN1(n1739), .IN2(n20169), .IN3(n1634), .IN4(n20140), .Q(
        n6059) );
  OA22X1 U29259 ( .IN1(n1911), .IN2(n20202), .IN3(n1825), .IN4(n20173), .Q(
        n6060) );
  OA22X1 U29260 ( .IN1(n2083), .IN2(n20235), .IN3(n1997), .IN4(n20206), .Q(
        n6061) );
  NAND4X0 U29261 ( .IN1(n6047), .IN2(n6048), .IN3(n6049), .IN4(n6050), .QN(
        s4_data_o[3]) );
  OA22X1 U29262 ( .IN1(n1738), .IN2(n20167), .IN3(n1633), .IN4(n20142), .Q(
        n6047) );
  OA22X1 U29263 ( .IN1(n1910), .IN2(n20200), .IN3(n1824), .IN4(n20175), .Q(
        n6048) );
  OA22X1 U29264 ( .IN1(n2082), .IN2(n20233), .IN3(n1996), .IN4(n20208), .Q(
        n6049) );
  NAND4X0 U29265 ( .IN1(n6043), .IN2(n6044), .IN3(n6045), .IN4(n6046), .QN(
        s4_data_o[4]) );
  OA22X1 U29266 ( .IN1(n1737), .IN2(n20168), .IN3(n1632), .IN4(n20157), .Q(
        n6043) );
  OA22X1 U29267 ( .IN1(n1909), .IN2(n20201), .IN3(n1823), .IN4(n20190), .Q(
        n6044) );
  OA22X1 U29268 ( .IN1(n2081), .IN2(n20234), .IN3(n1995), .IN4(n20223), .Q(
        n6045) );
  NAND4X0 U29269 ( .IN1(n6039), .IN2(n6040), .IN3(n6041), .IN4(n6042), .QN(
        s4_data_o[5]) );
  OA22X1 U29270 ( .IN1(n1736), .IN2(n20169), .IN3(n1631), .IN4(n20155), .Q(
        n6039) );
  OA22X1 U29271 ( .IN1(n1908), .IN2(n20202), .IN3(n1822), .IN4(n20188), .Q(
        n6040) );
  OA22X1 U29272 ( .IN1(n2080), .IN2(n20235), .IN3(n1994), .IN4(n20221), .Q(
        n6041) );
  NAND4X0 U29273 ( .IN1(n6035), .IN2(n6036), .IN3(n6037), .IN4(n6038), .QN(
        s4_data_o[6]) );
  OA22X1 U29274 ( .IN1(n1735), .IN2(n20165), .IN3(n1630), .IN4(n20155), .Q(
        n6035) );
  OA22X1 U29275 ( .IN1(n1907), .IN2(n20198), .IN3(n1821), .IN4(n20188), .Q(
        n6036) );
  OA22X1 U29276 ( .IN1(n2079), .IN2(n20231), .IN3(n1993), .IN4(n20221), .Q(
        n6037) );
  NAND4X0 U29277 ( .IN1(n6031), .IN2(n6032), .IN3(n6033), .IN4(n6034), .QN(
        s4_data_o[7]) );
  OA22X1 U29278 ( .IN1(n1734), .IN2(n20163), .IN3(n1629), .IN4(n20155), .Q(
        n6031) );
  OA22X1 U29279 ( .IN1(n1906), .IN2(n20196), .IN3(n1820), .IN4(n20188), .Q(
        n6032) );
  OA22X1 U29280 ( .IN1(n2078), .IN2(n20229), .IN3(n1992), .IN4(n20221), .Q(
        n6033) );
  NAND4X0 U29281 ( .IN1(n6027), .IN2(n6028), .IN3(n6029), .IN4(n6030), .QN(
        s4_data_o[8]) );
  OA22X1 U29282 ( .IN1(n1733), .IN2(n20170), .IN3(n1628), .IN4(n20155), .Q(
        n6027) );
  OA22X1 U29283 ( .IN1(n1905), .IN2(n20203), .IN3(n1819), .IN4(n20188), .Q(
        n6028) );
  OA22X1 U29284 ( .IN1(n2077), .IN2(n20236), .IN3(n1991), .IN4(n20221), .Q(
        n6029) );
  NAND4X0 U29285 ( .IN1(n6023), .IN2(n6024), .IN3(n6025), .IN4(n6026), .QN(
        s4_data_o[9]) );
  OA22X1 U29286 ( .IN1(n1732), .IN2(n20163), .IN3(n1627), .IN4(n20156), .Q(
        n6023) );
  OA22X1 U29287 ( .IN1(n1904), .IN2(n20196), .IN3(n1818), .IN4(n20189), .Q(
        n6024) );
  OA22X1 U29288 ( .IN1(n2076), .IN2(n20229), .IN3(n1990), .IN4(n20222), .Q(
        n6025) );
  NAND4X0 U29289 ( .IN1(n6143), .IN2(n6144), .IN3(n6145), .IN4(n6146), .QN(
        s4_data_o[10]) );
  OA22X1 U29290 ( .IN1(n1731), .IN2(n20165), .IN3(n1626), .IN4(n20150), .Q(
        n6143) );
  OA22X1 U29291 ( .IN1(n1903), .IN2(n20198), .IN3(n1817), .IN4(n20183), .Q(
        n6144) );
  OA22X1 U29292 ( .IN1(n2075), .IN2(n20231), .IN3(n1989), .IN4(n20216), .Q(
        n6145) );
  NAND4X0 U29293 ( .IN1(n6139), .IN2(n6140), .IN3(n6141), .IN4(n6142), .QN(
        s4_data_o[11]) );
  OA22X1 U29294 ( .IN1(n1730), .IN2(n20170), .IN3(n1625), .IN4(n20150), .Q(
        n6139) );
  OA22X1 U29295 ( .IN1(n1902), .IN2(n20203), .IN3(n1816), .IN4(n20183), .Q(
        n6140) );
  OA22X1 U29296 ( .IN1(n2074), .IN2(n20236), .IN3(n1988), .IN4(n20216), .Q(
        n6141) );
  NAND4X0 U29297 ( .IN1(n6135), .IN2(n6136), .IN3(n6137), .IN4(n6138), .QN(
        s4_data_o[12]) );
  OA22X1 U29298 ( .IN1(n1729), .IN2(n20166), .IN3(n1624), .IN4(n20150), .Q(
        n6135) );
  OA22X1 U29299 ( .IN1(n1901), .IN2(n20199), .IN3(n1815), .IN4(n20183), .Q(
        n6136) );
  OA22X1 U29300 ( .IN1(n2073), .IN2(n20232), .IN3(n1987), .IN4(n20216), .Q(
        n6137) );
  NAND4X0 U29301 ( .IN1(n6131), .IN2(n6132), .IN3(n6133), .IN4(n6134), .QN(
        s4_data_o[13]) );
  OA22X1 U29302 ( .IN1(n1728), .IN2(n20167), .IN3(n1623), .IN4(n20144), .Q(
        n6131) );
  OA22X1 U29303 ( .IN1(n1900), .IN2(n20200), .IN3(n1814), .IN4(n20177), .Q(
        n6132) );
  OA22X1 U29304 ( .IN1(n2072), .IN2(n20233), .IN3(n1986), .IN4(n20210), .Q(
        n6133) );
  NAND4X0 U29305 ( .IN1(n6127), .IN2(n6128), .IN3(n6129), .IN4(n6130), .QN(
        s4_data_o[14]) );
  OA22X1 U29306 ( .IN1(n1727), .IN2(n20167), .IN3(n1622), .IN4(n20149), .Q(
        n6127) );
  OA22X1 U29307 ( .IN1(n1899), .IN2(n20200), .IN3(n1813), .IN4(n20182), .Q(
        n6128) );
  OA22X1 U29308 ( .IN1(n2071), .IN2(n20233), .IN3(n1985), .IN4(n20215), .Q(
        n6129) );
  NAND4X0 U29309 ( .IN1(n6123), .IN2(n6124), .IN3(n6125), .IN4(n6126), .QN(
        s4_data_o[15]) );
  OA22X1 U29310 ( .IN1(n1726), .IN2(n20167), .IN3(n1621), .IN4(n20150), .Q(
        n6123) );
  OA22X1 U29311 ( .IN1(n1898), .IN2(n20200), .IN3(n1812), .IN4(n20183), .Q(
        n6124) );
  OA22X1 U29312 ( .IN1(n2070), .IN2(n20233), .IN3(n1984), .IN4(n20216), .Q(
        n6125) );
  NAND4X0 U29313 ( .IN1(n6119), .IN2(n6120), .IN3(n6121), .IN4(n6122), .QN(
        s4_data_o[16]) );
  OA22X1 U29314 ( .IN1(n1725), .IN2(n20167), .IN3(n1620), .IN4(n20151), .Q(
        n6119) );
  OA22X1 U29315 ( .IN1(n1897), .IN2(n20200), .IN3(n1811), .IN4(n20184), .Q(
        n6120) );
  OA22X1 U29316 ( .IN1(n2069), .IN2(n20233), .IN3(n1983), .IN4(n20217), .Q(
        n6121) );
  NAND4X0 U29317 ( .IN1(n6115), .IN2(n6116), .IN3(n6117), .IN4(n6118), .QN(
        s4_data_o[17]) );
  OA22X1 U29318 ( .IN1(n1724), .IN2(n20168), .IN3(n1619), .IN4(n20151), .Q(
        n6115) );
  OA22X1 U29319 ( .IN1(n1896), .IN2(n20201), .IN3(n1810), .IN4(n20184), .Q(
        n6116) );
  OA22X1 U29320 ( .IN1(n2068), .IN2(n20234), .IN3(n1982), .IN4(n20217), .Q(
        n6117) );
  NAND4X0 U29321 ( .IN1(n6111), .IN2(n6112), .IN3(n6113), .IN4(n6114), .QN(
        s4_data_o[18]) );
  OA22X1 U29322 ( .IN1(n1723), .IN2(n20168), .IN3(n1618), .IN4(n20151), .Q(
        n6111) );
  OA22X1 U29323 ( .IN1(n1895), .IN2(n20201), .IN3(n1809), .IN4(n20184), .Q(
        n6112) );
  OA22X1 U29324 ( .IN1(n2067), .IN2(n20234), .IN3(n1981), .IN4(n20217), .Q(
        n6113) );
  NAND4X0 U29325 ( .IN1(n6107), .IN2(n6108), .IN3(n6109), .IN4(n6110), .QN(
        s4_data_o[19]) );
  OA22X1 U29326 ( .IN1(n1722), .IN2(n20168), .IN3(n1617), .IN4(n20151), .Q(
        n6107) );
  OA22X1 U29327 ( .IN1(n1894), .IN2(n20201), .IN3(n1808), .IN4(n20184), .Q(
        n6108) );
  OA22X1 U29328 ( .IN1(n2066), .IN2(n20234), .IN3(n1980), .IN4(n20217), .Q(
        n6109) );
  NAND4X0 U29329 ( .IN1(n6099), .IN2(n6100), .IN3(n6101), .IN4(n6102), .QN(
        s4_data_o[20]) );
  OA22X1 U29330 ( .IN1(n1721), .IN2(n20169), .IN3(n1616), .IN4(n20148), .Q(
        n6099) );
  OA22X1 U29331 ( .IN1(n1893), .IN2(n20202), .IN3(n1807), .IN4(n20181), .Q(
        n6100) );
  OA22X1 U29332 ( .IN1(n2065), .IN2(n20235), .IN3(n1979), .IN4(n20214), .Q(
        n6101) );
  NAND4X0 U29333 ( .IN1(n6095), .IN2(n6096), .IN3(n6097), .IN4(n6098), .QN(
        s4_data_o[21]) );
  OA22X1 U29334 ( .IN1(n1720), .IN2(n20169), .IN3(n1615), .IN4(n20152), .Q(
        n6095) );
  OA22X1 U29335 ( .IN1(n1892), .IN2(n20202), .IN3(n1806), .IN4(n20185), .Q(
        n6096) );
  OA22X1 U29336 ( .IN1(n2064), .IN2(n20235), .IN3(n1978), .IN4(n20218), .Q(
        n6097) );
  NAND4X0 U29337 ( .IN1(n6091), .IN2(n6092), .IN3(n6093), .IN4(n6094), .QN(
        s4_data_o[22]) );
  OA22X1 U29338 ( .IN1(n1719), .IN2(n20167), .IN3(n1614), .IN4(n20152), .Q(
        n6091) );
  OA22X1 U29339 ( .IN1(n1891), .IN2(n20200), .IN3(n1805), .IN4(n20185), .Q(
        n6092) );
  OA22X1 U29340 ( .IN1(n2063), .IN2(n20233), .IN3(n1977), .IN4(n20218), .Q(
        n6093) );
  NAND4X0 U29341 ( .IN1(n6087), .IN2(n6088), .IN3(n6089), .IN4(n6090), .QN(
        s4_data_o[23]) );
  OA22X1 U29342 ( .IN1(n1718), .IN2(n20168), .IN3(n1613), .IN4(n20152), .Q(
        n6087) );
  OA22X1 U29343 ( .IN1(n1890), .IN2(n20201), .IN3(n1804), .IN4(n20185), .Q(
        n6088) );
  OA22X1 U29344 ( .IN1(n2062), .IN2(n20234), .IN3(n1976), .IN4(n20218), .Q(
        n6089) );
  NAND4X0 U29345 ( .IN1(n6083), .IN2(n6084), .IN3(n6085), .IN4(n6086), .QN(
        s4_data_o[24]) );
  OA22X1 U29346 ( .IN1(n1717), .IN2(n20166), .IN3(n1612), .IN4(n20153), .Q(
        n6083) );
  OA22X1 U29347 ( .IN1(n1889), .IN2(n20199), .IN3(n1803), .IN4(n20186), .Q(
        n6084) );
  OA22X1 U29348 ( .IN1(n2061), .IN2(n20232), .IN3(n1975), .IN4(n20219), .Q(
        n6085) );
  NAND4X0 U29349 ( .IN1(n6079), .IN2(n6080), .IN3(n6081), .IN4(n6082), .QN(
        s4_data_o[25]) );
  OA22X1 U29350 ( .IN1(n1716), .IN2(n20166), .IN3(n1611), .IN4(n20153), .Q(
        n6079) );
  OA22X1 U29351 ( .IN1(n1888), .IN2(n20199), .IN3(n1802), .IN4(n20186), .Q(
        n6080) );
  OA22X1 U29352 ( .IN1(n2060), .IN2(n20232), .IN3(n1974), .IN4(n20219), .Q(
        n6081) );
  NAND4X0 U29353 ( .IN1(n6075), .IN2(n6076), .IN3(n6077), .IN4(n6078), .QN(
        s4_data_o[26]) );
  OA22X1 U29354 ( .IN1(n1715), .IN2(n20165), .IN3(n1610), .IN4(n20153), .Q(
        n6075) );
  OA22X1 U29355 ( .IN1(n1887), .IN2(n20198), .IN3(n1801), .IN4(n20186), .Q(
        n6076) );
  OA22X1 U29356 ( .IN1(n2059), .IN2(n20231), .IN3(n1973), .IN4(n20219), .Q(
        n6077) );
  NAND4X0 U29357 ( .IN1(n6071), .IN2(n6072), .IN3(n6073), .IN4(n6074), .QN(
        s4_data_o[27]) );
  OA22X1 U29358 ( .IN1(n1714), .IN2(n20168), .IN3(n1609), .IN4(n20154), .Q(
        n6071) );
  OA22X1 U29359 ( .IN1(n1886), .IN2(n20201), .IN3(n1800), .IN4(n20187), .Q(
        n6072) );
  OA22X1 U29360 ( .IN1(n2058), .IN2(n20234), .IN3(n1972), .IN4(n20220), .Q(
        n6073) );
  NAND4X0 U29361 ( .IN1(n6067), .IN2(n6068), .IN3(n6069), .IN4(n6070), .QN(
        s4_data_o[28]) );
  OA22X1 U29362 ( .IN1(n1713), .IN2(n20169), .IN3(n1608), .IN4(n20154), .Q(
        n6067) );
  OA22X1 U29363 ( .IN1(n1885), .IN2(n20202), .IN3(n1799), .IN4(n20187), .Q(
        n6068) );
  OA22X1 U29364 ( .IN1(n2057), .IN2(n20235), .IN3(n1971), .IN4(n20220), .Q(
        n6069) );
  NAND4X0 U29365 ( .IN1(n6063), .IN2(n6064), .IN3(n6065), .IN4(n6066), .QN(
        s4_data_o[29]) );
  OA22X1 U29366 ( .IN1(n1712), .IN2(n20169), .IN3(n1607), .IN4(n20154), .Q(
        n6063) );
  OA22X1 U29367 ( .IN1(n1884), .IN2(n20202), .IN3(n1798), .IN4(n20187), .Q(
        n6064) );
  OA22X1 U29368 ( .IN1(n2056), .IN2(n20235), .IN3(n1970), .IN4(n20220), .Q(
        n6065) );
  NAND4X0 U29369 ( .IN1(n6055), .IN2(n6056), .IN3(n6057), .IN4(n6058), .QN(
        s4_data_o[30]) );
  OA22X1 U29370 ( .IN1(n1711), .IN2(n20169), .IN3(n1606), .IN4(n20156), .Q(
        n6055) );
  OA22X1 U29371 ( .IN1(n1883), .IN2(n20202), .IN3(n1797), .IN4(n20189), .Q(
        n6056) );
  OA22X1 U29372 ( .IN1(n2055), .IN2(n20235), .IN3(n1969), .IN4(n20222), .Q(
        n6057) );
  NAND4X0 U29373 ( .IN1(n6051), .IN2(n6052), .IN3(n6053), .IN4(n6054), .QN(
        s4_data_o[31]) );
  OA22X1 U29374 ( .IN1(n1710), .IN2(n20167), .IN3(n1605), .IN4(n20141), .Q(
        n6051) );
  OA22X1 U29375 ( .IN1(n1882), .IN2(n20200), .IN3(n1796), .IN4(n20174), .Q(
        n6052) );
  OA22X1 U29376 ( .IN1(n2054), .IN2(n20233), .IN3(n1968), .IN4(n20207), .Q(
        n6053) );
  NAND4X0 U29377 ( .IN1(n6291), .IN2(n6292), .IN3(n6293), .IN4(n6294), .QN(
        s3_stb_o) );
  OA22X1 U29378 ( .IN1(n1795), .IN2(n6301), .IN3(n1709), .IN4(n6302), .Q(n6291) );
  OA22X1 U29379 ( .IN1(n1967), .IN2(n6299), .IN3(n1881), .IN4(n6300), .Q(n6292) );
  OA22X1 U29380 ( .IN1(n2139), .IN2(n6297), .IN3(n2053), .IN4(n6298), .Q(n6293) );
  NAND4X0 U29381 ( .IN1(n6279), .IN2(n6280), .IN3(n6281), .IN4(n6282), .QN(
        s3_we_o) );
  OA22X1 U29382 ( .IN1(n1794), .IN2(n20032), .IN3(n1708), .IN4(n20026), .Q(
        n6279) );
  OA22X1 U29383 ( .IN1(n1966), .IN2(n20065), .IN3(n1880), .IN4(n20042), .Q(
        n6280) );
  OA22X1 U29384 ( .IN1(n2138), .IN2(n20097), .IN3(n2052), .IN4(n20091), .Q(
        n6281) );
  NAND4X0 U29385 ( .IN1(n6315), .IN2(n6316), .IN3(n6317), .IN4(n6318), .QN(
        s3_sel_o[0]) );
  OA22X1 U29386 ( .IN1(n1793), .IN2(n6289), .IN3(n1707), .IN4(n20024), .Q(
        n6315) );
  OA22X1 U29387 ( .IN1(n1965), .IN2(n20072), .IN3(n1879), .IN4(n20059), .Q(
        n6316) );
  OA22X1 U29388 ( .IN1(n2137), .IN2(n6285), .IN3(n2051), .IN4(n20092), .Q(
        n6317) );
  NAND4X0 U29389 ( .IN1(n6311), .IN2(n6312), .IN3(n6313), .IN4(n6314), .QN(
        s3_sel_o[1]) );
  OA22X1 U29390 ( .IN1(n1792), .IN2(n6289), .IN3(n1706), .IN4(n20024), .Q(
        n6311) );
  OA22X1 U29391 ( .IN1(n1964), .IN2(n20072), .IN3(n1878), .IN4(n20059), .Q(
        n6312) );
  OA22X1 U29392 ( .IN1(n2136), .IN2(n6285), .IN3(n2050), .IN4(n20092), .Q(
        n6313) );
  NAND4X0 U29393 ( .IN1(n6307), .IN2(n6308), .IN3(n6309), .IN4(n6310), .QN(
        s3_sel_o[2]) );
  OA22X1 U29394 ( .IN1(n1791), .IN2(n6289), .IN3(n1705), .IN4(n20026), .Q(
        n6307) );
  OA22X1 U29395 ( .IN1(n1963), .IN2(n20072), .IN3(n1877), .IN4(n20043), .Q(
        n6308) );
  OA22X1 U29396 ( .IN1(n2135), .IN2(n6285), .IN3(n2049), .IN4(n20091), .Q(
        n6309) );
  NAND4X0 U29397 ( .IN1(n6303), .IN2(n6304), .IN3(n6305), .IN4(n6306), .QN(
        s3_sel_o[3]) );
  OA22X1 U29398 ( .IN1(n1790), .IN2(n6289), .IN3(n1704), .IN4(n20026), .Q(
        n6303) );
  OA22X1 U29399 ( .IN1(n1962), .IN2(n20072), .IN3(n1876), .IN4(n20044), .Q(
        n6304) );
  OA22X1 U29400 ( .IN1(n2134), .IN2(n6285), .IN3(n2048), .IN4(n20091), .Q(
        n6305) );
  NAND4X0 U29401 ( .IN1(n6571), .IN2(n6572), .IN3(n6573), .IN4(n6574), .QN(
        s3_addr_o[0]) );
  OA22X1 U29402 ( .IN1(n1789), .IN2(n20032), .IN3(n1703), .IN4(n20009), .Q(
        n6571) );
  OA22X1 U29403 ( .IN1(n1961), .IN2(n20065), .IN3(n1875), .IN4(n20042), .Q(
        n6572) );
  OA22X1 U29404 ( .IN1(n2133), .IN2(n20097), .IN3(n2047), .IN4(n20075), .Q(
        n6573) );
  NAND4X0 U29405 ( .IN1(n6527), .IN2(n6528), .IN3(n6529), .IN4(n6530), .QN(
        s3_addr_o[1]) );
  OA22X1 U29406 ( .IN1(n1788), .IN2(n20034), .IN3(n1702), .IN4(n20012), .Q(
        n6527) );
  OA22X1 U29407 ( .IN1(n1960), .IN2(n20067), .IN3(n1874), .IN4(n20045), .Q(
        n6528) );
  OA22X1 U29408 ( .IN1(n2132), .IN2(n20099), .IN3(n2046), .IN4(n20078), .Q(
        n6529) );
  NAND4X0 U29409 ( .IN1(n6483), .IN2(n6484), .IN3(n6485), .IN4(n6486), .QN(
        s3_addr_o[2]) );
  OA22X1 U29410 ( .IN1(n1787), .IN2(n20032), .IN3(n1701), .IN4(n20016), .Q(
        n6483) );
  OA22X1 U29411 ( .IN1(n1959), .IN2(n20065), .IN3(n1873), .IN4(n20049), .Q(
        n6484) );
  OA22X1 U29412 ( .IN1(n2131), .IN2(n20101), .IN3(n2045), .IN4(n20091), .Q(
        n6485) );
  NAND4X0 U29413 ( .IN1(n6471), .IN2(n6472), .IN3(n6473), .IN4(n6474), .QN(
        s3_addr_o[3]) );
  OA22X1 U29414 ( .IN1(n1786), .IN2(n6289), .IN3(n1699), .IN4(n20017), .Q(
        n6471) );
  OA22X1 U29415 ( .IN1(n1958), .IN2(n20072), .IN3(n1872), .IN4(n20050), .Q(
        n6472) );
  OA22X1 U29416 ( .IN1(n2130), .IN2(n6285), .IN3(n2044), .IN4(n20082), .Q(
        n6473) );
  NAND4X0 U29417 ( .IN1(n6467), .IN2(n6468), .IN3(n6469), .IN4(n6470), .QN(
        s3_addr_o[4]) );
  OA22X1 U29418 ( .IN1(n1785), .IN2(n20035), .IN3(n1697), .IN4(n20017), .Q(
        n6467) );
  OA22X1 U29419 ( .IN1(n1957), .IN2(n20068), .IN3(n1871), .IN4(n20050), .Q(
        n6468) );
  OA22X1 U29420 ( .IN1(n2129), .IN2(n20100), .IN3(n2043), .IN4(n20082), .Q(
        n6469) );
  NAND4X0 U29421 ( .IN1(n6463), .IN2(n6464), .IN3(n6465), .IN4(n6466), .QN(
        s3_addr_o[5]) );
  OA22X1 U29422 ( .IN1(n1784), .IN2(n6289), .IN3(n1696), .IN4(n20018), .Q(
        n6463) );
  OA22X1 U29423 ( .IN1(n1956), .IN2(n20072), .IN3(n1870), .IN4(n20051), .Q(
        n6464) );
  OA22X1 U29424 ( .IN1(n2128), .IN2(n6285), .IN3(n2042), .IN4(n20082), .Q(
        n6465) );
  NAND4X0 U29425 ( .IN1(n6459), .IN2(n6460), .IN3(n6461), .IN4(n6462), .QN(
        s3_addr_o[6]) );
  OA22X1 U29426 ( .IN1(n1783), .IN2(n20036), .IN3(n1679), .IN4(n20018), .Q(
        n6459) );
  OA22X1 U29427 ( .IN1(n1955), .IN2(n20069), .IN3(n1869), .IN4(n20051), .Q(
        n6460) );
  OA22X1 U29428 ( .IN1(n2127), .IN2(n20102), .IN3(n2041), .IN4(n20082), .Q(
        n6461) );
  NAND4X0 U29429 ( .IN1(n6455), .IN2(n6456), .IN3(n6457), .IN4(n6458), .QN(
        s3_addr_o[7]) );
  OA22X1 U29430 ( .IN1(n1782), .IN2(n20036), .IN3(n1678), .IN4(n20018), .Q(
        n6455) );
  OA22X1 U29431 ( .IN1(n1954), .IN2(n20069), .IN3(n1868), .IN4(n20051), .Q(
        n6456) );
  OA22X1 U29432 ( .IN1(n2126), .IN2(n20102), .IN3(n2040), .IN4(n20082), .Q(
        n6457) );
  NAND4X0 U29433 ( .IN1(n6451), .IN2(n6452), .IN3(n6453), .IN4(n6454), .QN(
        s3_addr_o[8]) );
  OA22X1 U29434 ( .IN1(n1781), .IN2(n20036), .IN3(n1677), .IN4(n20019), .Q(
        n6451) );
  OA22X1 U29435 ( .IN1(n1953), .IN2(n20069), .IN3(n1867), .IN4(n20052), .Q(
        n6452) );
  OA22X1 U29436 ( .IN1(n2125), .IN2(n20102), .IN3(n2039), .IN4(n20083), .Q(
        n6453) );
  NAND4X0 U29437 ( .IN1(n6447), .IN2(n6448), .IN3(n6449), .IN4(n6450), .QN(
        s3_addr_o[9]) );
  OA22X1 U29438 ( .IN1(n1780), .IN2(n20036), .IN3(n1676), .IN4(n20019), .Q(
        n6447) );
  OA22X1 U29439 ( .IN1(n1952), .IN2(n20069), .IN3(n1866), .IN4(n20052), .Q(
        n6448) );
  OA22X1 U29440 ( .IN1(n2124), .IN2(n20102), .IN3(n2038), .IN4(n20083), .Q(
        n6449) );
  NAND4X0 U29441 ( .IN1(n6567), .IN2(n6568), .IN3(n6569), .IN4(n6570), .QN(
        s3_addr_o[10]) );
  OA22X1 U29442 ( .IN1(n1779), .IN2(n20032), .IN3(n1675), .IN4(n20009), .Q(
        n6567) );
  OA22X1 U29443 ( .IN1(n1951), .IN2(n20065), .IN3(n1865), .IN4(n20042), .Q(
        n6568) );
  OA22X1 U29444 ( .IN1(n2123), .IN2(n20097), .IN3(n2037), .IN4(n20075), .Q(
        n6569) );
  NAND4X0 U29445 ( .IN1(n6563), .IN2(n6564), .IN3(n6565), .IN4(n6566), .QN(
        s3_addr_o[11]) );
  OA22X1 U29446 ( .IN1(n1778), .IN2(n20032), .IN3(n1674), .IN4(n20009), .Q(
        n6563) );
  OA22X1 U29447 ( .IN1(n1950), .IN2(n20065), .IN3(n1864), .IN4(n20042), .Q(
        n6564) );
  OA22X1 U29448 ( .IN1(n2122), .IN2(n20097), .IN3(n2036), .IN4(n20075), .Q(
        n6565) );
  NAND4X0 U29449 ( .IN1(n6559), .IN2(n6560), .IN3(n6561), .IN4(n6562), .QN(
        s3_addr_o[12]) );
  OA22X1 U29450 ( .IN1(n1777), .IN2(n20032), .IN3(n1673), .IN4(n20010), .Q(
        n6559) );
  OA22X1 U29451 ( .IN1(n1949), .IN2(n20065), .IN3(n1863), .IN4(n20043), .Q(
        n6560) );
  OA22X1 U29452 ( .IN1(n2121), .IN2(n20097), .IN3(n2035), .IN4(n20076), .Q(
        n6561) );
  NAND4X0 U29453 ( .IN1(n6555), .IN2(n6556), .IN3(n6557), .IN4(n6558), .QN(
        s3_addr_o[13]) );
  OA22X1 U29454 ( .IN1(n1776), .IN2(n20033), .IN3(n1672), .IN4(n20010), .Q(
        n6555) );
  OA22X1 U29455 ( .IN1(n1948), .IN2(n20066), .IN3(n1862), .IN4(n20043), .Q(
        n6556) );
  OA22X1 U29456 ( .IN1(n2120), .IN2(n20098), .IN3(n2034), .IN4(n20076), .Q(
        n6557) );
  NAND4X0 U29457 ( .IN1(n6551), .IN2(n6552), .IN3(n6553), .IN4(n6554), .QN(
        s3_addr_o[14]) );
  OA22X1 U29458 ( .IN1(n1775), .IN2(n20033), .IN3(n1671), .IN4(n20010), .Q(
        n6551) );
  OA22X1 U29459 ( .IN1(n1947), .IN2(n20066), .IN3(n1861), .IN4(n20043), .Q(
        n6552) );
  OA22X1 U29460 ( .IN1(n2119), .IN2(n20098), .IN3(n2033), .IN4(n20076), .Q(
        n6553) );
  NAND4X0 U29461 ( .IN1(n6547), .IN2(n6548), .IN3(n6549), .IN4(n6550), .QN(
        s3_addr_o[15]) );
  OA22X1 U29462 ( .IN1(n1774), .IN2(n20033), .IN3(n1670), .IN4(n20011), .Q(
        n6547) );
  OA22X1 U29463 ( .IN1(n1946), .IN2(n20066), .IN3(n1860), .IN4(n20044), .Q(
        n6548) );
  OA22X1 U29464 ( .IN1(n2118), .IN2(n20098), .IN3(n2032), .IN4(n20077), .Q(
        n6549) );
  NAND4X0 U29465 ( .IN1(n6543), .IN2(n6544), .IN3(n6545), .IN4(n6546), .QN(
        s3_addr_o[16]) );
  OA22X1 U29466 ( .IN1(n1773), .IN2(n20033), .IN3(n1669), .IN4(n20011), .Q(
        n6543) );
  OA22X1 U29467 ( .IN1(n1945), .IN2(n20066), .IN3(n1859), .IN4(n20044), .Q(
        n6544) );
  OA22X1 U29468 ( .IN1(n2117), .IN2(n20098), .IN3(n2031), .IN4(n20077), .Q(
        n6545) );
  NAND4X0 U29469 ( .IN1(n6539), .IN2(n6540), .IN3(n6541), .IN4(n6542), .QN(
        s3_addr_o[17]) );
  OA22X1 U29470 ( .IN1(n1772), .IN2(n20034), .IN3(n1668), .IN4(n20011), .Q(
        n6539) );
  OA22X1 U29471 ( .IN1(n1944), .IN2(n20067), .IN3(n1858), .IN4(n20044), .Q(
        n6540) );
  OA22X1 U29472 ( .IN1(n2116), .IN2(n20099), .IN3(n2030), .IN4(n20077), .Q(
        n6541) );
  NAND4X0 U29473 ( .IN1(n6535), .IN2(n6536), .IN3(n6537), .IN4(n6538), .QN(
        s3_addr_o[18]) );
  OA22X1 U29474 ( .IN1(n1771), .IN2(n20034), .IN3(n1667), .IN4(n20012), .Q(
        n6535) );
  OA22X1 U29475 ( .IN1(n1943), .IN2(n20067), .IN3(n1857), .IN4(n20045), .Q(
        n6536) );
  OA22X1 U29476 ( .IN1(n2115), .IN2(n20099), .IN3(n2029), .IN4(n20078), .Q(
        n6537) );
  NAND4X0 U29477 ( .IN1(n6531), .IN2(n6532), .IN3(n6533), .IN4(n6534), .QN(
        s3_addr_o[19]) );
  OA22X1 U29478 ( .IN1(n1770), .IN2(n20034), .IN3(n1666), .IN4(n20012), .Q(
        n6531) );
  OA22X1 U29479 ( .IN1(n1942), .IN2(n20067), .IN3(n1856), .IN4(n20045), .Q(
        n6532) );
  OA22X1 U29480 ( .IN1(n2114), .IN2(n20099), .IN3(n2028), .IN4(n20078), .Q(
        n6533) );
  NAND4X0 U29481 ( .IN1(n6523), .IN2(n6524), .IN3(n6525), .IN4(n6526), .QN(
        s3_addr_o[20]) );
  OA22X1 U29482 ( .IN1(n1769), .IN2(n20033), .IN3(n1665), .IN4(n20013), .Q(
        n6523) );
  OA22X1 U29483 ( .IN1(n1941), .IN2(n20066), .IN3(n1855), .IN4(n20046), .Q(
        n6524) );
  OA22X1 U29484 ( .IN1(n2113), .IN2(n20098), .IN3(n2027), .IN4(n20079), .Q(
        n6525) );
  NAND4X0 U29485 ( .IN1(n6519), .IN2(n6520), .IN3(n6521), .IN4(n6522), .QN(
        s3_addr_o[21]) );
  OA22X1 U29486 ( .IN1(n1768), .IN2(n20033), .IN3(n1664), .IN4(n20013), .Q(
        n6519) );
  OA22X1 U29487 ( .IN1(n1940), .IN2(n20066), .IN3(n1854), .IN4(n20046), .Q(
        n6520) );
  OA22X1 U29488 ( .IN1(n2112), .IN2(n20098), .IN3(n2026), .IN4(n20079), .Q(
        n6521) );
  NAND4X0 U29489 ( .IN1(n6515), .IN2(n6516), .IN3(n6517), .IN4(n6518), .QN(
        s3_addr_o[22]) );
  OA22X1 U29490 ( .IN1(n1767), .IN2(n20032), .IN3(n1663), .IN4(n20013), .Q(
        n6515) );
  OA22X1 U29491 ( .IN1(n1939), .IN2(n20065), .IN3(n1853), .IN4(n20046), .Q(
        n6516) );
  OA22X1 U29492 ( .IN1(n2111), .IN2(n20097), .IN3(n2025), .IN4(n20079), .Q(
        n6517) );
  NAND4X0 U29493 ( .IN1(n6511), .IN2(n6512), .IN3(n6513), .IN4(n6514), .QN(
        s3_addr_o[23]) );
  OA22X1 U29494 ( .IN1(n1766), .IN2(n20033), .IN3(n1662), .IN4(n20014), .Q(
        n6511) );
  OA22X1 U29495 ( .IN1(n1938), .IN2(n20066), .IN3(n1852), .IN4(n20047), .Q(
        n6512) );
  OA22X1 U29496 ( .IN1(n2110), .IN2(n20098), .IN3(n2024), .IN4(n20080), .Q(
        n6513) );
  NAND4X0 U29497 ( .IN1(n6507), .IN2(n6508), .IN3(n6509), .IN4(n6510), .QN(
        s3_addr_o[24]) );
  OA22X1 U29498 ( .IN1(n1765), .IN2(n20035), .IN3(n1661), .IN4(n20014), .Q(
        n6507) );
  OA22X1 U29499 ( .IN1(n1937), .IN2(n20068), .IN3(n1851), .IN4(n20047), .Q(
        n6508) );
  OA22X1 U29500 ( .IN1(n2109), .IN2(n20100), .IN3(n2023), .IN4(n20080), .Q(
        n6509) );
  NAND4X0 U29501 ( .IN1(n6503), .IN2(n6504), .IN3(n6505), .IN4(n6506), .QN(
        s3_addr_o[25]) );
  OA22X1 U29502 ( .IN1(n1764), .IN2(n20035), .IN3(n1660), .IN4(n20014), .Q(
        n6503) );
  OA22X1 U29503 ( .IN1(n1936), .IN2(n20068), .IN3(n1850), .IN4(n20047), .Q(
        n6504) );
  OA22X1 U29504 ( .IN1(n2108), .IN2(n20100), .IN3(n2022), .IN4(n20080), .Q(
        n6505) );
  NAND4X0 U29505 ( .IN1(n6499), .IN2(n6500), .IN3(n6501), .IN4(n6502), .QN(
        s3_addr_o[26]) );
  OA22X1 U29506 ( .IN1(n1763), .IN2(n20035), .IN3(n1659), .IN4(n20015), .Q(
        n6499) );
  OA22X1 U29507 ( .IN1(n1935), .IN2(n20068), .IN3(n1849), .IN4(n20048), .Q(
        n6500) );
  OA22X1 U29508 ( .IN1(n2107), .IN2(n20100), .IN3(n2021), .IN4(n20081), .Q(
        n6501) );
  NAND4X0 U29509 ( .IN1(n6495), .IN2(n6496), .IN3(n6497), .IN4(n6498), .QN(
        s3_addr_o[27]) );
  OA22X1 U29510 ( .IN1(n1762), .IN2(n20035), .IN3(n1658), .IN4(n20015), .Q(
        n6495) );
  OA22X1 U29511 ( .IN1(n1934), .IN2(n20068), .IN3(n1848), .IN4(n20048), .Q(
        n6496) );
  OA22X1 U29512 ( .IN1(n2106), .IN2(n20100), .IN3(n2020), .IN4(n20081), .Q(
        n6497) );
  NAND4X0 U29513 ( .IN1(n6491), .IN2(n6492), .IN3(n6493), .IN4(n6494), .QN(
        s3_addr_o[28]) );
  OA22X1 U29514 ( .IN1(n1761), .IN2(n20035), .IN3(n1657), .IN4(n20015), .Q(
        n6491) );
  OA22X1 U29515 ( .IN1(n1933), .IN2(n20069), .IN3(n1847), .IN4(n20048), .Q(
        n6492) );
  OA22X1 U29516 ( .IN1(n2105), .IN2(n20101), .IN3(n2019), .IN4(n20081), .Q(
        n6493) );
  NAND4X0 U29517 ( .IN1(n6487), .IN2(n6488), .IN3(n6489), .IN4(n6490), .QN(
        s3_addr_o[29]) );
  OA22X1 U29518 ( .IN1(n1760), .IN2(n20036), .IN3(n1656), .IN4(n20016), .Q(
        n6487) );
  OA22X1 U29519 ( .IN1(n1932), .IN2(n20068), .IN3(n1846), .IN4(n20049), .Q(
        n6488) );
  OA22X1 U29520 ( .IN1(n2104), .IN2(n20101), .IN3(n2018), .IN4(n20082), .Q(
        n6489) );
  NAND4X0 U29521 ( .IN1(n6479), .IN2(n6480), .IN3(n6481), .IN4(n6482), .QN(
        s3_addr_o[30]) );
  OA22X1 U29522 ( .IN1(n1759), .IN2(n20035), .IN3(n1655), .IN4(n20016), .Q(
        n6479) );
  OA22X1 U29523 ( .IN1(n1931), .IN2(n20068), .IN3(n1845), .IN4(n20049), .Q(
        n6480) );
  OA22X1 U29524 ( .IN1(n2103), .IN2(n20101), .IN3(n2017), .IN4(n20082), .Q(
        n6481) );
  NAND4X0 U29525 ( .IN1(n6475), .IN2(n6476), .IN3(n6477), .IN4(n6478), .QN(
        s3_addr_o[31]) );
  OA22X1 U29526 ( .IN1(n1758), .IN2(n20039), .IN3(n1650), .IN4(n20017), .Q(
        n6475) );
  OA22X1 U29527 ( .IN1(n1930), .IN2(n20069), .IN3(n1844), .IN4(n20050), .Q(
        n6476) );
  OA22X1 U29528 ( .IN1(n2102), .IN2(n20101), .IN3(n2016), .IN4(n20082), .Q(
        n6477) );
  NAND4X0 U29529 ( .IN1(n6443), .IN2(n6444), .IN3(n6445), .IN4(n6446), .QN(
        s3_data_o[0]) );
  OA22X1 U29530 ( .IN1(n1741), .IN2(n20037), .IN3(n1636), .IN4(n20019), .Q(
        n6443) );
  OA22X1 U29531 ( .IN1(n1913), .IN2(n20067), .IN3(n1827), .IN4(n20052), .Q(
        n6444) );
  OA22X1 U29532 ( .IN1(n2085), .IN2(n20103), .IN3(n1999), .IN4(n20083), .Q(
        n6445) );
  NAND4X0 U29533 ( .IN1(n6399), .IN2(n6400), .IN3(n6401), .IN4(n6402), .QN(
        s3_data_o[1]) );
  OA22X1 U29534 ( .IN1(n1740), .IN2(n20038), .IN3(n1635), .IN4(n20021), .Q(
        n6399) );
  OA22X1 U29535 ( .IN1(n1912), .IN2(n20070), .IN3(n1826), .IN4(n20056), .Q(
        n6400) );
  OA22X1 U29536 ( .IN1(n2084), .IN2(n20099), .IN3(n1998), .IN4(n20086), .Q(
        n6401) );
  NAND4X0 U29537 ( .IN1(n6355), .IN2(n6356), .IN3(n6357), .IN4(n6358), .QN(
        s3_data_o[2]) );
  OA22X1 U29538 ( .IN1(n1739), .IN2(n20038), .IN3(n1634), .IN4(n20024), .Q(
        n6355) );
  OA22X1 U29539 ( .IN1(n1911), .IN2(n6287), .IN3(n1825), .IN4(n20059), .Q(
        n6356) );
  OA22X1 U29540 ( .IN1(n2083), .IN2(n20104), .IN3(n1997), .IN4(n20089), .Q(
        n6357) );
  NAND4X0 U29541 ( .IN1(n6343), .IN2(n6344), .IN3(n6345), .IN4(n6346), .QN(
        s3_data_o[3]) );
  OA22X1 U29542 ( .IN1(n1738), .IN2(n20033), .IN3(n1633), .IN4(n20024), .Q(
        n6343) );
  OA22X1 U29543 ( .IN1(n1910), .IN2(n20067), .IN3(n1824), .IN4(n20059), .Q(
        n6344) );
  OA22X1 U29544 ( .IN1(n2082), .IN2(n20104), .IN3(n1996), .IN4(n20090), .Q(
        n6345) );
  NAND4X0 U29545 ( .IN1(n6339), .IN2(n6340), .IN3(n6341), .IN4(n6342), .QN(
        s3_data_o[4]) );
  OA22X1 U29546 ( .IN1(n1737), .IN2(n20037), .IN3(n1632), .IN4(n20024), .Q(
        n6339) );
  OA22X1 U29547 ( .IN1(n1909), .IN2(n6287), .IN3(n1823), .IN4(n20059), .Q(
        n6340) );
  OA22X1 U29548 ( .IN1(n2081), .IN2(n20098), .IN3(n1995), .IN4(n20090), .Q(
        n6341) );
  NAND4X0 U29549 ( .IN1(n6335), .IN2(n6336), .IN3(n6337), .IN4(n6338), .QN(
        s3_data_o[5]) );
  OA22X1 U29550 ( .IN1(n1736), .IN2(n20038), .IN3(n1631), .IN4(n20024), .Q(
        n6335) );
  OA22X1 U29551 ( .IN1(n1908), .IN2(n20070), .IN3(n1822), .IN4(n20059), .Q(
        n6336) );
  OA22X1 U29552 ( .IN1(n2080), .IN2(n20102), .IN3(n1994), .IN4(n20090), .Q(
        n6337) );
  NAND4X0 U29553 ( .IN1(n6331), .IN2(n6332), .IN3(n6333), .IN4(n6334), .QN(
        s3_data_o[6]) );
  OA22X1 U29554 ( .IN1(n1735), .IN2(n20039), .IN3(n1630), .IN4(n20025), .Q(
        n6331) );
  OA22X1 U29555 ( .IN1(n1907), .IN2(n20071), .IN3(n1821), .IN4(n20057), .Q(
        n6332) );
  OA22X1 U29556 ( .IN1(n2079), .IN2(n20104), .IN3(n1993), .IN4(n20091), .Q(
        n6333) );
  NAND4X0 U29557 ( .IN1(n6327), .IN2(n6328), .IN3(n6329), .IN4(n6330), .QN(
        s3_data_o[7]) );
  OA22X1 U29558 ( .IN1(n1734), .IN2(n20039), .IN3(n1629), .IN4(n20025), .Q(
        n6327) );
  OA22X1 U29559 ( .IN1(n1906), .IN2(n20071), .IN3(n1820), .IN4(n20057), .Q(
        n6328) );
  OA22X1 U29560 ( .IN1(n2078), .IN2(n20104), .IN3(n1992), .IN4(n20091), .Q(
        n6329) );
  NAND4X0 U29561 ( .IN1(n6323), .IN2(n6324), .IN3(n6325), .IN4(n6326), .QN(
        s3_data_o[8]) );
  OA22X1 U29562 ( .IN1(n1733), .IN2(n20039), .IN3(n1628), .IN4(n20025), .Q(
        n6323) );
  OA22X1 U29563 ( .IN1(n1905), .IN2(n20071), .IN3(n1819), .IN4(n20057), .Q(
        n6324) );
  OA22X1 U29564 ( .IN1(n2077), .IN2(n20104), .IN3(n1991), .IN4(n20091), .Q(
        n6325) );
  NAND4X0 U29565 ( .IN1(n6319), .IN2(n6320), .IN3(n6321), .IN4(n6322), .QN(
        s3_data_o[9]) );
  OA22X1 U29566 ( .IN1(n1732), .IN2(n20039), .IN3(n1627), .IN4(n20024), .Q(
        n6319) );
  OA22X1 U29567 ( .IN1(n1904), .IN2(n20071), .IN3(n1818), .IN4(n20057), .Q(
        n6320) );
  OA22X1 U29568 ( .IN1(n2076), .IN2(n20104), .IN3(n1990), .IN4(n20092), .Q(
        n6321) );
  NAND4X0 U29569 ( .IN1(n6439), .IN2(n6440), .IN3(n6441), .IN4(n6442), .QN(
        s3_data_o[10]) );
  OA22X1 U29570 ( .IN1(n1731), .IN2(n20038), .IN3(n1626), .IN4(n20020), .Q(
        n6439) );
  OA22X1 U29571 ( .IN1(n1903), .IN2(n20072), .IN3(n1817), .IN4(n20053), .Q(
        n6440) );
  OA22X1 U29572 ( .IN1(n2075), .IN2(n20103), .IN3(n1989), .IN4(n20086), .Q(
        n6441) );
  NAND4X0 U29573 ( .IN1(n6435), .IN2(n6436), .IN3(n6437), .IN4(n6438), .QN(
        s3_data_o[11]) );
  OA22X1 U29574 ( .IN1(n1730), .IN2(n20039), .IN3(n1625), .IN4(n20020), .Q(
        n6435) );
  OA22X1 U29575 ( .IN1(n1902), .IN2(n20070), .IN3(n1816), .IN4(n20053), .Q(
        n6436) );
  OA22X1 U29576 ( .IN1(n2074), .IN2(n20103), .IN3(n1988), .IN4(n20087), .Q(
        n6437) );
  NAND4X0 U29577 ( .IN1(n6431), .IN2(n6432), .IN3(n6433), .IN4(n6434), .QN(
        s3_data_o[12]) );
  OA22X1 U29578 ( .IN1(n1729), .IN2(n20036), .IN3(n1624), .IN4(n20020), .Q(
        n6431) );
  OA22X1 U29579 ( .IN1(n1901), .IN2(n20071), .IN3(n1815), .IN4(n20053), .Q(
        n6432) );
  OA22X1 U29580 ( .IN1(n2073), .IN2(n20103), .IN3(n1987), .IN4(n20088), .Q(
        n6433) );
  NAND4X0 U29581 ( .IN1(n6427), .IN2(n6428), .IN3(n6429), .IN4(n6430), .QN(
        s3_data_o[13]) );
  OA22X1 U29582 ( .IN1(n1728), .IN2(n20037), .IN3(n1623), .IN4(n20021), .Q(
        n6427) );
  OA22X1 U29583 ( .IN1(n1900), .IN2(n20070), .IN3(n1814), .IN4(n20054), .Q(
        n6428) );
  OA22X1 U29584 ( .IN1(n2072), .IN2(n20104), .IN3(n1986), .IN4(n20084), .Q(
        n6429) );
  NAND4X0 U29585 ( .IN1(n6423), .IN2(n6424), .IN3(n6425), .IN4(n6426), .QN(
        s3_data_o[14]) );
  OA22X1 U29586 ( .IN1(n1727), .IN2(n20037), .IN3(n1622), .IN4(n20021), .Q(
        n6423) );
  OA22X1 U29587 ( .IN1(n1899), .IN2(n20070), .IN3(n1813), .IN4(n20054), .Q(
        n6424) );
  OA22X1 U29588 ( .IN1(n2071), .IN2(n20102), .IN3(n1985), .IN4(n20084), .Q(
        n6425) );
  NAND4X0 U29589 ( .IN1(n6419), .IN2(n6420), .IN3(n6421), .IN4(n6422), .QN(
        s3_data_o[15]) );
  OA22X1 U29590 ( .IN1(n1726), .IN2(n20037), .IN3(n1621), .IN4(n20021), .Q(
        n6419) );
  OA22X1 U29591 ( .IN1(n1898), .IN2(n20070), .IN3(n1812), .IN4(n20054), .Q(
        n6420) );
  OA22X1 U29592 ( .IN1(n2070), .IN2(n20099), .IN3(n1984), .IN4(n20084), .Q(
        n6421) );
  NAND4X0 U29593 ( .IN1(n6415), .IN2(n6416), .IN3(n6417), .IN4(n6418), .QN(
        s3_data_o[16]) );
  OA22X1 U29594 ( .IN1(n1725), .IN2(n20037), .IN3(n1620), .IN4(n20022), .Q(
        n6415) );
  OA22X1 U29595 ( .IN1(n1897), .IN2(n20070), .IN3(n1811), .IN4(n20055), .Q(
        n6416) );
  OA22X1 U29596 ( .IN1(n2069), .IN2(n20103), .IN3(n1983), .IN4(n20085), .Q(
        n6417) );
  NAND4X0 U29597 ( .IN1(n6411), .IN2(n6412), .IN3(n6413), .IN4(n6414), .QN(
        s3_data_o[17]) );
  OA22X1 U29598 ( .IN1(n1724), .IN2(n20038), .IN3(n1619), .IN4(n20022), .Q(
        n6411) );
  OA22X1 U29599 ( .IN1(n1896), .IN2(n20065), .IN3(n1810), .IN4(n20055), .Q(
        n6412) );
  OA22X1 U29600 ( .IN1(n2068), .IN2(n20103), .IN3(n1982), .IN4(n20085), .Q(
        n6413) );
  NAND4X0 U29601 ( .IN1(n6407), .IN2(n6408), .IN3(n6409), .IN4(n6410), .QN(
        s3_data_o[18]) );
  OA22X1 U29602 ( .IN1(n1723), .IN2(n20038), .IN3(n1618), .IN4(n20022), .Q(
        n6407) );
  OA22X1 U29603 ( .IN1(n1895), .IN2(n20072), .IN3(n1809), .IN4(n20055), .Q(
        n6408) );
  OA22X1 U29604 ( .IN1(n2067), .IN2(n20097), .IN3(n1981), .IN4(n20085), .Q(
        n6409) );
  NAND4X0 U29605 ( .IN1(n6403), .IN2(n6404), .IN3(n6405), .IN4(n6406), .QN(
        s3_data_o[19]) );
  OA22X1 U29606 ( .IN1(n1722), .IN2(n20038), .IN3(n1617), .IN4(n20022), .Q(
        n6403) );
  OA22X1 U29607 ( .IN1(n1894), .IN2(n6287), .IN3(n1808), .IN4(n20056), .Q(
        n6404) );
  OA22X1 U29608 ( .IN1(n2066), .IN2(n20100), .IN3(n1980), .IN4(n20087), .Q(
        n6405) );
  NAND4X0 U29609 ( .IN1(n6395), .IN2(n6396), .IN3(n6397), .IN4(n6398), .QN(
        s3_data_o[20]) );
  OA22X1 U29610 ( .IN1(n1721), .IN2(n20034), .IN3(n1616), .IN4(n20021), .Q(
        n6395) );
  OA22X1 U29611 ( .IN1(n1893), .IN2(n20071), .IN3(n1807), .IN4(n20056), .Q(
        n6396) );
  OA22X1 U29612 ( .IN1(n2065), .IN2(n20101), .IN3(n1979), .IN4(n20088), .Q(
        n6397) );
  NAND4X0 U29613 ( .IN1(n6391), .IN2(n6392), .IN3(n6393), .IN4(n6394), .QN(
        s3_data_o[21]) );
  OA22X1 U29614 ( .IN1(n1720), .IN2(n20037), .IN3(n1615), .IN4(n20024), .Q(
        n6391) );
  OA22X1 U29615 ( .IN1(n1892), .IN2(n6287), .IN3(n1806), .IN4(n20057), .Q(
        n6392) );
  OA22X1 U29616 ( .IN1(n2064), .IN2(n20100), .IN3(n1978), .IN4(n20086), .Q(
        n6393) );
  NAND4X0 U29617 ( .IN1(n6387), .IN2(n6388), .IN3(n6389), .IN4(n6390), .QN(
        s3_data_o[22]) );
  OA22X1 U29618 ( .IN1(n1719), .IN2(n20037), .IN3(n1614), .IN4(n20008), .Q(
        n6387) );
  OA22X1 U29619 ( .IN1(n1891), .IN2(n20070), .IN3(n1805), .IN4(n20057), .Q(
        n6388) );
  OA22X1 U29620 ( .IN1(n2063), .IN2(n20101), .IN3(n1977), .IN4(n20086), .Q(
        n6389) );
  NAND4X0 U29621 ( .IN1(n6383), .IN2(n6384), .IN3(n6385), .IN4(n6386), .QN(
        s3_data_o[23]) );
  OA22X1 U29622 ( .IN1(n1718), .IN2(n20038), .IN3(n1613), .IN4(n20026), .Q(
        n6383) );
  OA22X1 U29623 ( .IN1(n1890), .IN2(n20066), .IN3(n1804), .IN4(n20057), .Q(
        n6384) );
  OA22X1 U29624 ( .IN1(n2062), .IN2(n20097), .IN3(n1976), .IN4(n20086), .Q(
        n6385) );
  NAND4X0 U29625 ( .IN1(n6379), .IN2(n6380), .IN3(n6381), .IN4(n6382), .QN(
        s3_data_o[24]) );
  OA22X1 U29626 ( .IN1(n1717), .IN2(n20039), .IN3(n1612), .IN4(n20023), .Q(
        n6379) );
  OA22X1 U29627 ( .IN1(n1889), .IN2(n20071), .IN3(n1803), .IN4(n20058), .Q(
        n6380) );
  OA22X1 U29628 ( .IN1(n2061), .IN2(n20104), .IN3(n1975), .IN4(n20087), .Q(
        n6381) );
  NAND4X0 U29629 ( .IN1(n6375), .IN2(n6376), .IN3(n6377), .IN4(n6378), .QN(
        s3_data_o[25]) );
  OA22X1 U29630 ( .IN1(n1716), .IN2(n20036), .IN3(n1611), .IN4(n20023), .Q(
        n6375) );
  OA22X1 U29631 ( .IN1(n1888), .IN2(n20069), .IN3(n1802), .IN4(n20058), .Q(
        n6376) );
  OA22X1 U29632 ( .IN1(n2060), .IN2(n20102), .IN3(n1974), .IN4(n20087), .Q(
        n6377) );
  NAND4X0 U29633 ( .IN1(n6371), .IN2(n6372), .IN3(n6373), .IN4(n6374), .QN(
        s3_data_o[26]) );
  OA22X1 U29634 ( .IN1(n1715), .IN2(n20034), .IN3(n1610), .IN4(n20023), .Q(
        n6371) );
  OA22X1 U29635 ( .IN1(n1887), .IN2(n20067), .IN3(n1801), .IN4(n20058), .Q(
        n6372) );
  OA22X1 U29636 ( .IN1(n2059), .IN2(n20099), .IN3(n1973), .IN4(n20087), .Q(
        n6373) );
  NAND4X0 U29637 ( .IN1(n6367), .IN2(n6368), .IN3(n6369), .IN4(n6370), .QN(
        s3_data_o[27]) );
  OA22X1 U29638 ( .IN1(n1714), .IN2(n20034), .IN3(n1609), .IN4(n20026), .Q(
        n6367) );
  OA22X1 U29639 ( .IN1(n1886), .IN2(n20071), .IN3(n1800), .IN4(n20057), .Q(
        n6368) );
  OA22X1 U29640 ( .IN1(n2058), .IN2(n20103), .IN3(n1972), .IN4(n20088), .Q(
        n6369) );
  NAND4X0 U29641 ( .IN1(n6363), .IN2(n6364), .IN3(n6365), .IN4(n6366), .QN(
        s3_data_o[28]) );
  OA22X1 U29642 ( .IN1(n1713), .IN2(n20032), .IN3(n1608), .IN4(n20023), .Q(
        n6363) );
  OA22X1 U29643 ( .IN1(n1885), .IN2(n6287), .IN3(n1799), .IN4(n20058), .Q(
        n6364) );
  OA22X1 U29644 ( .IN1(n2057), .IN2(n20102), .IN3(n1971), .IN4(n20088), .Q(
        n6365) );
  NAND4X0 U29645 ( .IN1(n6359), .IN2(n6360), .IN3(n6361), .IN4(n6362), .QN(
        s3_data_o[29]) );
  OA22X1 U29646 ( .IN1(n1712), .IN2(n6289), .IN3(n1607), .IN4(n20025), .Q(
        n6359) );
  OA22X1 U29647 ( .IN1(n1884), .IN2(n6287), .IN3(n1798), .IN4(n20057), .Q(
        n6360) );
  OA22X1 U29648 ( .IN1(n2056), .IN2(n20099), .IN3(n1970), .IN4(n20088), .Q(
        n6361) );
  NAND4X0 U29649 ( .IN1(n6351), .IN2(n6352), .IN3(n6353), .IN4(n6354), .QN(
        s3_data_o[30]) );
  OA22X1 U29650 ( .IN1(n1711), .IN2(n6289), .IN3(n1606), .IN4(n20024), .Q(
        n6351) );
  OA22X1 U29651 ( .IN1(n1883), .IN2(n6287), .IN3(n1797), .IN4(n20059), .Q(
        n6352) );
  OA22X1 U29652 ( .IN1(n2055), .IN2(n20103), .IN3(n1969), .IN4(n20089), .Q(
        n6353) );
  NAND4X0 U29653 ( .IN1(n6347), .IN2(n6348), .IN3(n6349), .IN4(n6350), .QN(
        s3_data_o[31]) );
  OA22X1 U29654 ( .IN1(n1710), .IN2(n20034), .IN3(n1605), .IN4(n20024), .Q(
        n6347) );
  OA22X1 U29655 ( .IN1(n1882), .IN2(n20067), .IN3(n1796), .IN4(n20059), .Q(
        n6348) );
  OA22X1 U29656 ( .IN1(n2054), .IN2(n20100), .IN3(n1968), .IN4(n20089), .Q(
        n6349) );
  NAND4X0 U29657 ( .IN1(n6587), .IN2(n6588), .IN3(n6589), .IN4(n6590), .QN(
        s2_stb_o) );
  OA22X1 U29658 ( .IN1(n1795), .IN2(n6597), .IN3(n1709), .IN4(n6598), .Q(n6587) );
  OA22X1 U29659 ( .IN1(n1967), .IN2(n6595), .IN3(n1881), .IN4(n6596), .Q(n6588) );
  OA22X1 U29660 ( .IN1(n2139), .IN2(n6593), .IN3(n2053), .IN4(n6594), .Q(n6589) );
  NAND4X0 U29661 ( .IN1(n6575), .IN2(n6576), .IN3(n6577), .IN4(n6578), .QN(
        s2_we_o) );
  OA22X1 U29662 ( .IN1(n1794), .IN2(n19901), .IN3(n1708), .IN4(n19895), .Q(
        n6575) );
  OA22X1 U29663 ( .IN1(n1966), .IN2(n19934), .IN3(n1880), .IN4(n19911), .Q(
        n6576) );
  OA22X1 U29664 ( .IN1(n2138), .IN2(n19966), .IN3(n2052), .IN4(n19961), .Q(
        n6577) );
  NAND4X0 U29665 ( .IN1(n6611), .IN2(n6612), .IN3(n6613), .IN4(n6614), .QN(
        s2_sel_o[0]) );
  OA22X1 U29666 ( .IN1(n1793), .IN2(n6585), .IN3(n1707), .IN4(n19893), .Q(
        n6611) );
  OA22X1 U29667 ( .IN1(n1965), .IN2(n19941), .IN3(n1879), .IN4(n19928), .Q(
        n6612) );
  OA22X1 U29668 ( .IN1(n2137), .IN2(n6581), .IN3(n2051), .IN4(n19960), .Q(
        n6613) );
  NAND4X0 U29669 ( .IN1(n6607), .IN2(n6608), .IN3(n6609), .IN4(n6610), .QN(
        s2_sel_o[1]) );
  OA22X1 U29670 ( .IN1(n1792), .IN2(n6585), .IN3(n1706), .IN4(n19893), .Q(
        n6607) );
  OA22X1 U29671 ( .IN1(n1964), .IN2(n19941), .IN3(n1878), .IN4(n19928), .Q(
        n6608) );
  OA22X1 U29672 ( .IN1(n2136), .IN2(n6581), .IN3(n2050), .IN4(n19960), .Q(
        n6609) );
  NAND4X0 U29673 ( .IN1(n6603), .IN2(n6604), .IN3(n6605), .IN4(n6606), .QN(
        s2_sel_o[2]) );
  OA22X1 U29674 ( .IN1(n1791), .IN2(n6585), .IN3(n1705), .IN4(n19895), .Q(
        n6603) );
  OA22X1 U29675 ( .IN1(n1963), .IN2(n19941), .IN3(n1877), .IN4(n19912), .Q(
        n6604) );
  OA22X1 U29676 ( .IN1(n2135), .IN2(n6581), .IN3(n2049), .IN4(n19961), .Q(
        n6605) );
  NAND4X0 U29677 ( .IN1(n6599), .IN2(n6600), .IN3(n6601), .IN4(n6602), .QN(
        s2_sel_o[3]) );
  OA22X1 U29678 ( .IN1(n1790), .IN2(n6585), .IN3(n1704), .IN4(n19895), .Q(
        n6599) );
  OA22X1 U29679 ( .IN1(n1962), .IN2(n19941), .IN3(n1876), .IN4(n19913), .Q(
        n6600) );
  OA22X1 U29680 ( .IN1(n2134), .IN2(n6581), .IN3(n2048), .IN4(n19961), .Q(
        n6601) );
  NAND4X0 U29681 ( .IN1(n6867), .IN2(n6868), .IN3(n6869), .IN4(n6870), .QN(
        s2_addr_o[0]) );
  OA22X1 U29682 ( .IN1(n1789), .IN2(n19901), .IN3(n1703), .IN4(n19878), .Q(
        n6867) );
  OA22X1 U29683 ( .IN1(n1961), .IN2(n19934), .IN3(n1875), .IN4(n19911), .Q(
        n6868) );
  OA22X1 U29684 ( .IN1(n2133), .IN2(n19966), .IN3(n2047), .IN4(n19944), .Q(
        n6869) );
  NAND4X0 U29685 ( .IN1(n6823), .IN2(n6824), .IN3(n6825), .IN4(n6826), .QN(
        s2_addr_o[1]) );
  OA22X1 U29686 ( .IN1(n1788), .IN2(n19903), .IN3(n1702), .IN4(n19881), .Q(
        n6823) );
  OA22X1 U29687 ( .IN1(n1960), .IN2(n19936), .IN3(n1874), .IN4(n19914), .Q(
        n6824) );
  OA22X1 U29688 ( .IN1(n2132), .IN2(n19968), .IN3(n2046), .IN4(n19947), .Q(
        n6825) );
  NAND4X0 U29689 ( .IN1(n6779), .IN2(n6780), .IN3(n6781), .IN4(n6782), .QN(
        s2_addr_o[2]) );
  OA22X1 U29690 ( .IN1(n1787), .IN2(n19901), .IN3(n1701), .IN4(n19885), .Q(
        n6779) );
  OA22X1 U29691 ( .IN1(n1959), .IN2(n19934), .IN3(n1873), .IN4(n19918), .Q(
        n6780) );
  OA22X1 U29692 ( .IN1(n2131), .IN2(n19966), .IN3(n2045), .IN4(n19951), .Q(
        n6781) );
  NAND4X0 U29693 ( .IN1(n6767), .IN2(n6768), .IN3(n6769), .IN4(n6770), .QN(
        s2_addr_o[3]) );
  OA22X1 U29694 ( .IN1(n1786), .IN2(n6585), .IN3(n1699), .IN4(n19886), .Q(
        n6767) );
  OA22X1 U29695 ( .IN1(n1958), .IN2(n19941), .IN3(n1872), .IN4(n19919), .Q(
        n6768) );
  OA22X1 U29696 ( .IN1(n2130), .IN2(n6581), .IN3(n2044), .IN4(n19951), .Q(
        n6769) );
  NAND4X0 U29697 ( .IN1(n6763), .IN2(n6764), .IN3(n6765), .IN4(n6766), .QN(
        s2_addr_o[4]) );
  OA22X1 U29698 ( .IN1(n1785), .IN2(n19904), .IN3(n1697), .IN4(n19886), .Q(
        n6763) );
  OA22X1 U29699 ( .IN1(n1957), .IN2(n19937), .IN3(n1871), .IN4(n19919), .Q(
        n6764) );
  OA22X1 U29700 ( .IN1(n2129), .IN2(n19969), .IN3(n2043), .IN4(n19951), .Q(
        n6765) );
  NAND4X0 U29701 ( .IN1(n6759), .IN2(n6760), .IN3(n6761), .IN4(n6762), .QN(
        s2_addr_o[5]) );
  OA22X1 U29702 ( .IN1(n1784), .IN2(n6585), .IN3(n1696), .IN4(n19887), .Q(
        n6759) );
  OA22X1 U29703 ( .IN1(n1956), .IN2(n19941), .IN3(n1870), .IN4(n19920), .Q(
        n6760) );
  OA22X1 U29704 ( .IN1(n2128), .IN2(n6581), .IN3(n2042), .IN4(n19951), .Q(
        n6761) );
  NAND4X0 U29705 ( .IN1(n6755), .IN2(n6756), .IN3(n6757), .IN4(n6758), .QN(
        s2_addr_o[6]) );
  OA22X1 U29706 ( .IN1(n1783), .IN2(n19905), .IN3(n1679), .IN4(n19887), .Q(
        n6755) );
  OA22X1 U29707 ( .IN1(n1955), .IN2(n19938), .IN3(n1869), .IN4(n19920), .Q(
        n6756) );
  OA22X1 U29708 ( .IN1(n2127), .IN2(n19970), .IN3(n2041), .IN4(n19951), .Q(
        n6757) );
  NAND4X0 U29709 ( .IN1(n6751), .IN2(n6752), .IN3(n6753), .IN4(n6754), .QN(
        s2_addr_o[7]) );
  OA22X1 U29710 ( .IN1(n1782), .IN2(n19905), .IN3(n1678), .IN4(n19887), .Q(
        n6751) );
  OA22X1 U29711 ( .IN1(n1954), .IN2(n19938), .IN3(n1868), .IN4(n19920), .Q(
        n6752) );
  OA22X1 U29712 ( .IN1(n2126), .IN2(n19970), .IN3(n2040), .IN4(n19951), .Q(
        n6753) );
  NAND4X0 U29713 ( .IN1(n6747), .IN2(n6748), .IN3(n6749), .IN4(n6750), .QN(
        s2_addr_o[8]) );
  OA22X1 U29714 ( .IN1(n1781), .IN2(n19905), .IN3(n1677), .IN4(n19888), .Q(
        n6747) );
  OA22X1 U29715 ( .IN1(n1953), .IN2(n19938), .IN3(n1867), .IN4(n19921), .Q(
        n6748) );
  OA22X1 U29716 ( .IN1(n2125), .IN2(n19970), .IN3(n2039), .IN4(n19952), .Q(
        n6749) );
  NAND4X0 U29717 ( .IN1(n6743), .IN2(n6744), .IN3(n6745), .IN4(n6746), .QN(
        s2_addr_o[9]) );
  OA22X1 U29718 ( .IN1(n1780), .IN2(n19905), .IN3(n1676), .IN4(n19888), .Q(
        n6743) );
  OA22X1 U29719 ( .IN1(n1952), .IN2(n19938), .IN3(n1866), .IN4(n19921), .Q(
        n6744) );
  OA22X1 U29720 ( .IN1(n2124), .IN2(n19970), .IN3(n2038), .IN4(n19952), .Q(
        n6745) );
  NAND4X0 U29721 ( .IN1(n6863), .IN2(n6864), .IN3(n6865), .IN4(n6866), .QN(
        s2_addr_o[10]) );
  OA22X1 U29722 ( .IN1(n1779), .IN2(n19901), .IN3(n1675), .IN4(n19878), .Q(
        n6863) );
  OA22X1 U29723 ( .IN1(n1951), .IN2(n19934), .IN3(n1865), .IN4(n19911), .Q(
        n6864) );
  OA22X1 U29724 ( .IN1(n2123), .IN2(n19966), .IN3(n2037), .IN4(n19944), .Q(
        n6865) );
  NAND4X0 U29725 ( .IN1(n6859), .IN2(n6860), .IN3(n6861), .IN4(n6862), .QN(
        s2_addr_o[11]) );
  OA22X1 U29726 ( .IN1(n1778), .IN2(n19901), .IN3(n1674), .IN4(n19878), .Q(
        n6859) );
  OA22X1 U29727 ( .IN1(n1950), .IN2(n19934), .IN3(n1864), .IN4(n19911), .Q(
        n6860) );
  OA22X1 U29728 ( .IN1(n2122), .IN2(n19966), .IN3(n2036), .IN4(n19944), .Q(
        n6861) );
  NAND4X0 U29729 ( .IN1(n6855), .IN2(n6856), .IN3(n6857), .IN4(n6858), .QN(
        s2_addr_o[12]) );
  OA22X1 U29730 ( .IN1(n1777), .IN2(n19901), .IN3(n1673), .IN4(n19879), .Q(
        n6855) );
  OA22X1 U29731 ( .IN1(n1949), .IN2(n19934), .IN3(n1863), .IN4(n19912), .Q(
        n6856) );
  OA22X1 U29732 ( .IN1(n2121), .IN2(n19966), .IN3(n2035), .IN4(n19945), .Q(
        n6857) );
  NAND4X0 U29733 ( .IN1(n6851), .IN2(n6852), .IN3(n6853), .IN4(n6854), .QN(
        s2_addr_o[13]) );
  OA22X1 U29734 ( .IN1(n1776), .IN2(n19902), .IN3(n1672), .IN4(n19879), .Q(
        n6851) );
  OA22X1 U29735 ( .IN1(n1948), .IN2(n19935), .IN3(n1862), .IN4(n19912), .Q(
        n6852) );
  OA22X1 U29736 ( .IN1(n2120), .IN2(n19967), .IN3(n2034), .IN4(n19945), .Q(
        n6853) );
  NAND4X0 U29737 ( .IN1(n6847), .IN2(n6848), .IN3(n6849), .IN4(n6850), .QN(
        s2_addr_o[14]) );
  OA22X1 U29738 ( .IN1(n1775), .IN2(n19902), .IN3(n1671), .IN4(n19879), .Q(
        n6847) );
  OA22X1 U29739 ( .IN1(n1947), .IN2(n19935), .IN3(n1861), .IN4(n19912), .Q(
        n6848) );
  OA22X1 U29740 ( .IN1(n2119), .IN2(n19967), .IN3(n2033), .IN4(n19945), .Q(
        n6849) );
  NAND4X0 U29741 ( .IN1(n6843), .IN2(n6844), .IN3(n6845), .IN4(n6846), .QN(
        s2_addr_o[15]) );
  OA22X1 U29742 ( .IN1(n1774), .IN2(n19902), .IN3(n1670), .IN4(n19880), .Q(
        n6843) );
  OA22X1 U29743 ( .IN1(n1946), .IN2(n19935), .IN3(n1860), .IN4(n19913), .Q(
        n6844) );
  OA22X1 U29744 ( .IN1(n2118), .IN2(n19967), .IN3(n2032), .IN4(n19946), .Q(
        n6845) );
  NAND4X0 U29745 ( .IN1(n6839), .IN2(n6840), .IN3(n6841), .IN4(n6842), .QN(
        s2_addr_o[16]) );
  OA22X1 U29746 ( .IN1(n1773), .IN2(n19902), .IN3(n1669), .IN4(n19880), .Q(
        n6839) );
  OA22X1 U29747 ( .IN1(n1945), .IN2(n19935), .IN3(n1859), .IN4(n19913), .Q(
        n6840) );
  OA22X1 U29748 ( .IN1(n2117), .IN2(n19967), .IN3(n2031), .IN4(n19946), .Q(
        n6841) );
  NAND4X0 U29749 ( .IN1(n6835), .IN2(n6836), .IN3(n6837), .IN4(n6838), .QN(
        s2_addr_o[17]) );
  OA22X1 U29750 ( .IN1(n1772), .IN2(n19903), .IN3(n1668), .IN4(n19880), .Q(
        n6835) );
  OA22X1 U29751 ( .IN1(n1944), .IN2(n19936), .IN3(n1858), .IN4(n19913), .Q(
        n6836) );
  OA22X1 U29752 ( .IN1(n2116), .IN2(n19968), .IN3(n2030), .IN4(n19946), .Q(
        n6837) );
  NAND4X0 U29753 ( .IN1(n6831), .IN2(n6832), .IN3(n6833), .IN4(n6834), .QN(
        s2_addr_o[18]) );
  OA22X1 U29754 ( .IN1(n1771), .IN2(n19903), .IN3(n1667), .IN4(n19881), .Q(
        n6831) );
  OA22X1 U29755 ( .IN1(n1943), .IN2(n19936), .IN3(n1857), .IN4(n19914), .Q(
        n6832) );
  OA22X1 U29756 ( .IN1(n2115), .IN2(n19968), .IN3(n2029), .IN4(n19947), .Q(
        n6833) );
  NAND4X0 U29757 ( .IN1(n6827), .IN2(n6828), .IN3(n6829), .IN4(n6830), .QN(
        s2_addr_o[19]) );
  OA22X1 U29758 ( .IN1(n1770), .IN2(n19903), .IN3(n1666), .IN4(n19881), .Q(
        n6827) );
  OA22X1 U29759 ( .IN1(n1942), .IN2(n19936), .IN3(n1856), .IN4(n19914), .Q(
        n6828) );
  OA22X1 U29760 ( .IN1(n2114), .IN2(n19968), .IN3(n2028), .IN4(n19947), .Q(
        n6829) );
  NAND4X0 U29761 ( .IN1(n6819), .IN2(n6820), .IN3(n6821), .IN4(n6822), .QN(
        s2_addr_o[20]) );
  OA22X1 U29762 ( .IN1(n1769), .IN2(n19902), .IN3(n1665), .IN4(n19882), .Q(
        n6819) );
  OA22X1 U29763 ( .IN1(n1941), .IN2(n19935), .IN3(n1855), .IN4(n19915), .Q(
        n6820) );
  OA22X1 U29764 ( .IN1(n2113), .IN2(n19967), .IN3(n2027), .IN4(n19948), .Q(
        n6821) );
  NAND4X0 U29765 ( .IN1(n6815), .IN2(n6816), .IN3(n6817), .IN4(n6818), .QN(
        s2_addr_o[21]) );
  OA22X1 U29766 ( .IN1(n1768), .IN2(n19902), .IN3(n1664), .IN4(n19882), .Q(
        n6815) );
  OA22X1 U29767 ( .IN1(n1940), .IN2(n19935), .IN3(n1854), .IN4(n19915), .Q(
        n6816) );
  OA22X1 U29768 ( .IN1(n2112), .IN2(n19967), .IN3(n2026), .IN4(n19948), .Q(
        n6817) );
  NAND4X0 U29769 ( .IN1(n6811), .IN2(n6812), .IN3(n6813), .IN4(n6814), .QN(
        s2_addr_o[22]) );
  OA22X1 U29770 ( .IN1(n1767), .IN2(n19901), .IN3(n1663), .IN4(n19882), .Q(
        n6811) );
  OA22X1 U29771 ( .IN1(n1939), .IN2(n19934), .IN3(n1853), .IN4(n19915), .Q(
        n6812) );
  OA22X1 U29772 ( .IN1(n2111), .IN2(n19966), .IN3(n2025), .IN4(n19948), .Q(
        n6813) );
  NAND4X0 U29773 ( .IN1(n6807), .IN2(n6808), .IN3(n6809), .IN4(n6810), .QN(
        s2_addr_o[23]) );
  OA22X1 U29774 ( .IN1(n1766), .IN2(n19902), .IN3(n1662), .IN4(n19883), .Q(
        n6807) );
  OA22X1 U29775 ( .IN1(n1938), .IN2(n19935), .IN3(n1852), .IN4(n19916), .Q(
        n6808) );
  OA22X1 U29776 ( .IN1(n2110), .IN2(n19967), .IN3(n2024), .IN4(n19949), .Q(
        n6809) );
  NAND4X0 U29777 ( .IN1(n6803), .IN2(n6804), .IN3(n6805), .IN4(n6806), .QN(
        s2_addr_o[24]) );
  OA22X1 U29778 ( .IN1(n1765), .IN2(n19904), .IN3(n1661), .IN4(n19883), .Q(
        n6803) );
  OA22X1 U29779 ( .IN1(n1937), .IN2(n19937), .IN3(n1851), .IN4(n19916), .Q(
        n6804) );
  OA22X1 U29780 ( .IN1(n2109), .IN2(n19969), .IN3(n2023), .IN4(n19949), .Q(
        n6805) );
  NAND4X0 U29781 ( .IN1(n6799), .IN2(n6800), .IN3(n6801), .IN4(n6802), .QN(
        s2_addr_o[25]) );
  OA22X1 U29782 ( .IN1(n1764), .IN2(n19904), .IN3(n1660), .IN4(n19883), .Q(
        n6799) );
  OA22X1 U29783 ( .IN1(n1936), .IN2(n19937), .IN3(n1850), .IN4(n19916), .Q(
        n6800) );
  OA22X1 U29784 ( .IN1(n2108), .IN2(n19969), .IN3(n2022), .IN4(n19949), .Q(
        n6801) );
  NAND4X0 U29785 ( .IN1(n6795), .IN2(n6796), .IN3(n6797), .IN4(n6798), .QN(
        s2_addr_o[26]) );
  OA22X1 U29786 ( .IN1(n1763), .IN2(n19904), .IN3(n1659), .IN4(n19884), .Q(
        n6795) );
  OA22X1 U29787 ( .IN1(n1935), .IN2(n19937), .IN3(n1849), .IN4(n19917), .Q(
        n6796) );
  OA22X1 U29788 ( .IN1(n2107), .IN2(n19969), .IN3(n2021), .IN4(n19950), .Q(
        n6797) );
  NAND4X0 U29789 ( .IN1(n6791), .IN2(n6792), .IN3(n6793), .IN4(n6794), .QN(
        s2_addr_o[27]) );
  OA22X1 U29790 ( .IN1(n1762), .IN2(n19904), .IN3(n1658), .IN4(n19884), .Q(
        n6791) );
  OA22X1 U29791 ( .IN1(n1934), .IN2(n19937), .IN3(n1848), .IN4(n19917), .Q(
        n6792) );
  OA22X1 U29792 ( .IN1(n2106), .IN2(n19969), .IN3(n2020), .IN4(n19950), .Q(
        n6793) );
  NAND4X0 U29793 ( .IN1(n6787), .IN2(n6788), .IN3(n6789), .IN4(n6790), .QN(
        s2_addr_o[28]) );
  OA22X1 U29794 ( .IN1(n1761), .IN2(n19904), .IN3(n1657), .IN4(n19884), .Q(
        n6787) );
  OA22X1 U29795 ( .IN1(n1933), .IN2(n19937), .IN3(n1847), .IN4(n19917), .Q(
        n6788) );
  OA22X1 U29796 ( .IN1(n2105), .IN2(n19969), .IN3(n2019), .IN4(n19950), .Q(
        n6789) );
  NAND4X0 U29797 ( .IN1(n6783), .IN2(n6784), .IN3(n6785), .IN4(n6786), .QN(
        s2_addr_o[29]) );
  OA22X1 U29798 ( .IN1(n1760), .IN2(n19903), .IN3(n1656), .IN4(n19885), .Q(
        n6783) );
  OA22X1 U29799 ( .IN1(n1932), .IN2(n19936), .IN3(n1846), .IN4(n19918), .Q(
        n6784) );
  OA22X1 U29800 ( .IN1(n2104), .IN2(n19970), .IN3(n2018), .IN4(n19951), .Q(
        n6785) );
  NAND4X0 U29801 ( .IN1(n6775), .IN2(n6776), .IN3(n6777), .IN4(n6778), .QN(
        s2_addr_o[30]) );
  OA22X1 U29802 ( .IN1(n1759), .IN2(n19904), .IN3(n1655), .IN4(n19885), .Q(
        n6775) );
  OA22X1 U29803 ( .IN1(n1931), .IN2(n19937), .IN3(n1845), .IN4(n19918), .Q(
        n6776) );
  OA22X1 U29804 ( .IN1(n2103), .IN2(n19969), .IN3(n2017), .IN4(n19951), .Q(
        n6777) );
  NAND4X0 U29805 ( .IN1(n6771), .IN2(n6772), .IN3(n6773), .IN4(n6774), .QN(
        s2_addr_o[31]) );
  OA22X1 U29806 ( .IN1(n1758), .IN2(n19905), .IN3(n1650), .IN4(n19886), .Q(
        n6771) );
  OA22X1 U29807 ( .IN1(n1930), .IN2(n19938), .IN3(n1844), .IN4(n19919), .Q(
        n6772) );
  OA22X1 U29808 ( .IN1(n2102), .IN2(n19973), .IN3(n2016), .IN4(n19951), .Q(
        n6773) );
  NAND4X0 U29809 ( .IN1(n6739), .IN2(n6740), .IN3(n6741), .IN4(n6742), .QN(
        s2_data_o[0]) );
  OA22X1 U29810 ( .IN1(n1741), .IN2(n19906), .IN3(n1636), .IN4(n19888), .Q(
        n6739) );
  OA22X1 U29811 ( .IN1(n1913), .IN2(n19939), .IN3(n1827), .IN4(n19921), .Q(
        n6740) );
  OA22X1 U29812 ( .IN1(n2085), .IN2(n19972), .IN3(n1999), .IN4(n19952), .Q(
        n6741) );
  NAND4X0 U29813 ( .IN1(n6695), .IN2(n6696), .IN3(n6697), .IN4(n6698), .QN(
        s2_data_o[1]) );
  OA22X1 U29814 ( .IN1(n1740), .IN2(n19908), .IN3(n1635), .IN4(n19890), .Q(
        n6695) );
  OA22X1 U29815 ( .IN1(n1912), .IN2(n19934), .IN3(n1826), .IN4(n19925), .Q(
        n6696) );
  OA22X1 U29816 ( .IN1(n2084), .IN2(n19972), .IN3(n1998), .IN4(n19956), .Q(
        n6697) );
  NAND4X0 U29817 ( .IN1(n6651), .IN2(n6652), .IN3(n6653), .IN4(n6654), .QN(
        s2_data_o[2]) );
  OA22X1 U29818 ( .IN1(n1739), .IN2(n19908), .IN3(n1634), .IN4(n19893), .Q(
        n6651) );
  OA22X1 U29819 ( .IN1(n1911), .IN2(n6583), .IN3(n1825), .IN4(n19928), .Q(
        n6652) );
  OA22X1 U29820 ( .IN1(n2083), .IN2(n19971), .IN3(n1997), .IN4(n19959), .Q(
        n6653) );
  NAND4X0 U29821 ( .IN1(n6639), .IN2(n6640), .IN3(n6641), .IN4(n6642), .QN(
        s2_data_o[3]) );
  OA22X1 U29822 ( .IN1(n1738), .IN2(n19902), .IN3(n1633), .IN4(n19893), .Q(
        n6639) );
  OA22X1 U29823 ( .IN1(n1910), .IN2(n6583), .IN3(n1824), .IN4(n19928), .Q(
        n6640) );
  OA22X1 U29824 ( .IN1(n2082), .IN2(n19968), .IN3(n1996), .IN4(n19958), .Q(
        n6641) );
  NAND4X0 U29825 ( .IN1(n6635), .IN2(n6636), .IN3(n6637), .IN4(n6638), .QN(
        s2_data_o[4]) );
  OA22X1 U29826 ( .IN1(n1737), .IN2(n19907), .IN3(n1632), .IN4(n19893), .Q(
        n6635) );
  OA22X1 U29827 ( .IN1(n1909), .IN2(n19940), .IN3(n1823), .IN4(n19928), .Q(
        n6636) );
  OA22X1 U29828 ( .IN1(n2081), .IN2(n19971), .IN3(n1995), .IN4(n19958), .Q(
        n6637) );
  NAND4X0 U29829 ( .IN1(n6631), .IN2(n6632), .IN3(n6633), .IN4(n6634), .QN(
        s2_data_o[5]) );
  OA22X1 U29830 ( .IN1(n1736), .IN2(n19908), .IN3(n1631), .IN4(n19893), .Q(
        n6631) );
  OA22X1 U29831 ( .IN1(n1908), .IN2(n19935), .IN3(n1822), .IN4(n19928), .Q(
        n6632) );
  OA22X1 U29832 ( .IN1(n2080), .IN2(n19972), .IN3(n1994), .IN4(n19958), .Q(
        n6633) );
  NAND4X0 U29833 ( .IN1(n6627), .IN2(n6628), .IN3(n6629), .IN4(n6630), .QN(
        s2_data_o[6]) );
  OA22X1 U29834 ( .IN1(n1735), .IN2(n19907), .IN3(n1630), .IN4(n19894), .Q(
        n6627) );
  OA22X1 U29835 ( .IN1(n1907), .IN2(n19940), .IN3(n1821), .IN4(n19926), .Q(
        n6628) );
  OA22X1 U29836 ( .IN1(n2079), .IN2(n19973), .IN3(n1993), .IN4(n19959), .Q(
        n6629) );
  NAND4X0 U29837 ( .IN1(n6623), .IN2(n6624), .IN3(n6625), .IN4(n6626), .QN(
        s2_data_o[7]) );
  OA22X1 U29838 ( .IN1(n1734), .IN2(n19908), .IN3(n1629), .IN4(n19894), .Q(
        n6623) );
  OA22X1 U29839 ( .IN1(n1906), .IN2(n19939), .IN3(n1820), .IN4(n19926), .Q(
        n6624) );
  OA22X1 U29840 ( .IN1(n2078), .IN2(n19973), .IN3(n1992), .IN4(n19959), .Q(
        n6625) );
  NAND4X0 U29841 ( .IN1(n6619), .IN2(n6620), .IN3(n6621), .IN4(n6622), .QN(
        s2_data_o[8]) );
  OA22X1 U29842 ( .IN1(n1733), .IN2(n19905), .IN3(n1628), .IN4(n19894), .Q(
        n6619) );
  OA22X1 U29843 ( .IN1(n1905), .IN2(n19938), .IN3(n1819), .IN4(n19926), .Q(
        n6620) );
  OA22X1 U29844 ( .IN1(n2077), .IN2(n19973), .IN3(n1991), .IN4(n19959), .Q(
        n6621) );
  NAND4X0 U29845 ( .IN1(n6615), .IN2(n6616), .IN3(n6617), .IN4(n6618), .QN(
        s2_data_o[9]) );
  OA22X1 U29846 ( .IN1(n1732), .IN2(n19903), .IN3(n1627), .IN4(n19893), .Q(
        n6615) );
  OA22X1 U29847 ( .IN1(n1904), .IN2(n19936), .IN3(n1818), .IN4(n19926), .Q(
        n6616) );
  OA22X1 U29848 ( .IN1(n2076), .IN2(n19973), .IN3(n1990), .IN4(n19960), .Q(
        n6617) );
  NAND4X0 U29849 ( .IN1(n6735), .IN2(n6736), .IN3(n6737), .IN4(n6738), .QN(
        s2_data_o[10]) );
  OA22X1 U29850 ( .IN1(n1731), .IN2(n19906), .IN3(n1626), .IN4(n19889), .Q(
        n6735) );
  OA22X1 U29851 ( .IN1(n1903), .IN2(n19939), .IN3(n1817), .IN4(n19922), .Q(
        n6736) );
  OA22X1 U29852 ( .IN1(n2075), .IN2(n19968), .IN3(n1989), .IN4(n19953), .Q(
        n6737) );
  NAND4X0 U29853 ( .IN1(n6731), .IN2(n6732), .IN3(n6733), .IN4(n6734), .QN(
        s2_data_o[11]) );
  OA22X1 U29854 ( .IN1(n1730), .IN2(n19906), .IN3(n1625), .IN4(n19889), .Q(
        n6731) );
  OA22X1 U29855 ( .IN1(n1902), .IN2(n19939), .IN3(n1816), .IN4(n19922), .Q(
        n6732) );
  OA22X1 U29856 ( .IN1(n2074), .IN2(n19973), .IN3(n1988), .IN4(n19953), .Q(
        n6733) );
  NAND4X0 U29857 ( .IN1(n6727), .IN2(n6728), .IN3(n6729), .IN4(n6730), .QN(
        s2_data_o[12]) );
  OA22X1 U29858 ( .IN1(n1729), .IN2(n19906), .IN3(n1624), .IN4(n19889), .Q(
        n6727) );
  OA22X1 U29859 ( .IN1(n1901), .IN2(n19939), .IN3(n1815), .IN4(n19922), .Q(
        n6728) );
  OA22X1 U29860 ( .IN1(n2073), .IN2(n19970), .IN3(n1987), .IN4(n19953), .Q(
        n6729) );
  NAND4X0 U29861 ( .IN1(n6723), .IN2(n6724), .IN3(n6725), .IN4(n6726), .QN(
        s2_data_o[13]) );
  OA22X1 U29862 ( .IN1(n1728), .IN2(n19907), .IN3(n1623), .IN4(n19890), .Q(
        n6723) );
  OA22X1 U29863 ( .IN1(n1900), .IN2(n19940), .IN3(n1814), .IN4(n19923), .Q(
        n6724) );
  OA22X1 U29864 ( .IN1(n2072), .IN2(n19971), .IN3(n1986), .IN4(n19954), .Q(
        n6725) );
  NAND4X0 U29865 ( .IN1(n6719), .IN2(n6720), .IN3(n6721), .IN4(n6722), .QN(
        s2_data_o[14]) );
  OA22X1 U29866 ( .IN1(n1727), .IN2(n19907), .IN3(n1622), .IN4(n19890), .Q(
        n6719) );
  OA22X1 U29867 ( .IN1(n1899), .IN2(n19940), .IN3(n1813), .IN4(n19923), .Q(
        n6720) );
  OA22X1 U29868 ( .IN1(n2071), .IN2(n19971), .IN3(n1985), .IN4(n19954), .Q(
        n6721) );
  NAND4X0 U29869 ( .IN1(n6715), .IN2(n6716), .IN3(n6717), .IN4(n6718), .QN(
        s2_data_o[15]) );
  OA22X1 U29870 ( .IN1(n1726), .IN2(n19907), .IN3(n1621), .IN4(n19890), .Q(
        n6715) );
  OA22X1 U29871 ( .IN1(n1898), .IN2(n19940), .IN3(n1812), .IN4(n19923), .Q(
        n6716) );
  OA22X1 U29872 ( .IN1(n2070), .IN2(n19971), .IN3(n1984), .IN4(n19954), .Q(
        n6717) );
  NAND4X0 U29873 ( .IN1(n6711), .IN2(n6712), .IN3(n6713), .IN4(n6714), .QN(
        s2_data_o[16]) );
  OA22X1 U29874 ( .IN1(n1725), .IN2(n19907), .IN3(n1620), .IN4(n19891), .Q(
        n6711) );
  OA22X1 U29875 ( .IN1(n1897), .IN2(n19940), .IN3(n1811), .IN4(n19924), .Q(
        n6712) );
  OA22X1 U29876 ( .IN1(n2069), .IN2(n19971), .IN3(n1983), .IN4(n19955), .Q(
        n6713) );
  NAND4X0 U29877 ( .IN1(n6707), .IN2(n6708), .IN3(n6709), .IN4(n6710), .QN(
        s2_data_o[17]) );
  OA22X1 U29878 ( .IN1(n1724), .IN2(n19908), .IN3(n1619), .IN4(n19891), .Q(
        n6707) );
  OA22X1 U29879 ( .IN1(n1896), .IN2(n19941), .IN3(n1810), .IN4(n19924), .Q(
        n6708) );
  OA22X1 U29880 ( .IN1(n2068), .IN2(n19972), .IN3(n1982), .IN4(n19955), .Q(
        n6709) );
  NAND4X0 U29881 ( .IN1(n6703), .IN2(n6704), .IN3(n6705), .IN4(n6706), .QN(
        s2_data_o[18]) );
  OA22X1 U29882 ( .IN1(n1723), .IN2(n19908), .IN3(n1618), .IN4(n19891), .Q(
        n6703) );
  OA22X1 U29883 ( .IN1(n1895), .IN2(n6583), .IN3(n1809), .IN4(n19924), .Q(
        n6704) );
  OA22X1 U29884 ( .IN1(n2067), .IN2(n19972), .IN3(n1981), .IN4(n19955), .Q(
        n6705) );
  NAND4X0 U29885 ( .IN1(n6699), .IN2(n6700), .IN3(n6701), .IN4(n6702), .QN(
        s2_data_o[19]) );
  OA22X1 U29886 ( .IN1(n1722), .IN2(n19908), .IN3(n1617), .IN4(n19891), .Q(
        n6699) );
  OA22X1 U29887 ( .IN1(n1894), .IN2(n6583), .IN3(n1808), .IN4(n19925), .Q(
        n6700) );
  OA22X1 U29888 ( .IN1(n2066), .IN2(n19972), .IN3(n1980), .IN4(n19956), .Q(
        n6701) );
  NAND4X0 U29889 ( .IN1(n6691), .IN2(n6692), .IN3(n6693), .IN4(n6694), .QN(
        s2_data_o[20]) );
  OA22X1 U29890 ( .IN1(n1721), .IN2(n19906), .IN3(n1616), .IN4(n19890), .Q(
        n6691) );
  OA22X1 U29891 ( .IN1(n1893), .IN2(n19939), .IN3(n1807), .IN4(n19925), .Q(
        n6692) );
  OA22X1 U29892 ( .IN1(n2065), .IN2(n19972), .IN3(n1979), .IN4(n19956), .Q(
        n6693) );
  NAND4X0 U29893 ( .IN1(n6687), .IN2(n6688), .IN3(n6689), .IN4(n6690), .QN(
        s2_data_o[21]) );
  OA22X1 U29894 ( .IN1(n1720), .IN2(n19907), .IN3(n1615), .IN4(n19893), .Q(
        n6687) );
  OA22X1 U29895 ( .IN1(n1892), .IN2(n6583), .IN3(n1806), .IN4(n19926), .Q(
        n6688) );
  OA22X1 U29896 ( .IN1(n2064), .IN2(n19966), .IN3(n1978), .IN4(n19957), .Q(
        n6689) );
  NAND4X0 U29897 ( .IN1(n6683), .IN2(n6684), .IN3(n6685), .IN4(n6686), .QN(
        s2_data_o[22]) );
  OA22X1 U29898 ( .IN1(n1719), .IN2(n19907), .IN3(n1614), .IN4(n19877), .Q(
        n6683) );
  OA22X1 U29899 ( .IN1(n1891), .IN2(n19940), .IN3(n1805), .IN4(n19926), .Q(
        n6684) );
  OA22X1 U29900 ( .IN1(n2063), .IN2(n6581), .IN3(n1977), .IN4(n19957), .Q(
        n6685) );
  NAND4X0 U29901 ( .IN1(n6679), .IN2(n6680), .IN3(n6681), .IN4(n6682), .QN(
        s2_data_o[23]) );
  OA22X1 U29902 ( .IN1(n1718), .IN2(n19908), .IN3(n1613), .IN4(n19895), .Q(
        n6679) );
  OA22X1 U29903 ( .IN1(n1890), .IN2(n19940), .IN3(n1804), .IN4(n19926), .Q(
        n6680) );
  OA22X1 U29904 ( .IN1(n2062), .IN2(n6581), .IN3(n1976), .IN4(n19957), .Q(
        n6681) );
  NAND4X0 U29905 ( .IN1(n6675), .IN2(n6676), .IN3(n6677), .IN4(n6678), .QN(
        s2_data_o[24]) );
  OA22X1 U29906 ( .IN1(n1717), .IN2(n19906), .IN3(n1612), .IN4(n19892), .Q(
        n6675) );
  OA22X1 U29907 ( .IN1(n1889), .IN2(n19941), .IN3(n1803), .IN4(n19927), .Q(
        n6676) );
  OA22X1 U29908 ( .IN1(n2061), .IN2(n19973), .IN3(n1975), .IN4(n19958), .Q(
        n6677) );
  NAND4X0 U29909 ( .IN1(n6671), .IN2(n6672), .IN3(n6673), .IN4(n6674), .QN(
        s2_data_o[25]) );
  OA22X1 U29910 ( .IN1(n1716), .IN2(n19905), .IN3(n1611), .IN4(n19892), .Q(
        n6671) );
  OA22X1 U29911 ( .IN1(n1888), .IN2(n19938), .IN3(n1802), .IN4(n19927), .Q(
        n6672) );
  OA22X1 U29912 ( .IN1(n2060), .IN2(n19970), .IN3(n1974), .IN4(n19959), .Q(
        n6673) );
  NAND4X0 U29913 ( .IN1(n6667), .IN2(n6668), .IN3(n6669), .IN4(n6670), .QN(
        s2_data_o[26]) );
  OA22X1 U29914 ( .IN1(n1715), .IN2(n19903), .IN3(n1610), .IN4(n19892), .Q(
        n6667) );
  OA22X1 U29915 ( .IN1(n1887), .IN2(n19936), .IN3(n1801), .IN4(n19927), .Q(
        n6668) );
  OA22X1 U29916 ( .IN1(n2059), .IN2(n19968), .IN3(n1973), .IN4(n19961), .Q(
        n6669) );
  NAND4X0 U29917 ( .IN1(n6663), .IN2(n6664), .IN3(n6665), .IN4(n6666), .QN(
        s2_data_o[27]) );
  OA22X1 U29918 ( .IN1(n1714), .IN2(n19906), .IN3(n1609), .IN4(n19895), .Q(
        n6663) );
  OA22X1 U29919 ( .IN1(n1886), .IN2(n19939), .IN3(n1800), .IN4(n19926), .Q(
        n6664) );
  OA22X1 U29920 ( .IN1(n2058), .IN2(n19971), .IN3(n1972), .IN4(n19958), .Q(
        n6665) );
  NAND4X0 U29921 ( .IN1(n6659), .IN2(n6660), .IN3(n6661), .IN4(n6662), .QN(
        s2_data_o[28]) );
  OA22X1 U29922 ( .IN1(n1713), .IN2(n19901), .IN3(n1608), .IN4(n19892), .Q(
        n6659) );
  OA22X1 U29923 ( .IN1(n1885), .IN2(n6583), .IN3(n1799), .IN4(n19927), .Q(
        n6660) );
  OA22X1 U29924 ( .IN1(n2057), .IN2(n19972), .IN3(n1971), .IN4(n19945), .Q(
        n6661) );
  NAND4X0 U29925 ( .IN1(n6655), .IN2(n6656), .IN3(n6657), .IN4(n6658), .QN(
        s2_data_o[29]) );
  OA22X1 U29926 ( .IN1(n1712), .IN2(n6585), .IN3(n1607), .IN4(n19894), .Q(
        n6655) );
  OA22X1 U29927 ( .IN1(n1884), .IN2(n6583), .IN3(n1798), .IN4(n19926), .Q(
        n6656) );
  OA22X1 U29928 ( .IN1(n2056), .IN2(n19967), .IN3(n1970), .IN4(n19946), .Q(
        n6657) );
  NAND4X0 U29929 ( .IN1(n6647), .IN2(n6648), .IN3(n6649), .IN4(n6650), .QN(
        s2_data_o[30]) );
  OA22X1 U29930 ( .IN1(n1711), .IN2(n6585), .IN3(n1606), .IN4(n19893), .Q(
        n6647) );
  OA22X1 U29931 ( .IN1(n1883), .IN2(n6583), .IN3(n1797), .IN4(n19928), .Q(
        n6648) );
  OA22X1 U29932 ( .IN1(n2055), .IN2(n19968), .IN3(n1969), .IN4(n19961), .Q(
        n6649) );
  NAND4X0 U29933 ( .IN1(n6643), .IN2(n6644), .IN3(n6645), .IN4(n6646), .QN(
        s2_data_o[31]) );
  OA22X1 U29934 ( .IN1(n1710), .IN2(n19906), .IN3(n1605), .IN4(n19893), .Q(
        n6643) );
  OA22X1 U29935 ( .IN1(n1882), .IN2(n19939), .IN3(n1796), .IN4(n19928), .Q(
        n6644) );
  OA22X1 U29936 ( .IN1(n2054), .IN2(n19971), .IN3(n1968), .IN4(n19944), .Q(
        n6645) );
  NAND4X0 U29937 ( .IN1(n6883), .IN2(n6884), .IN3(n6885), .IN4(n6886), .QN(
        s1_stb_o) );
  OA22X1 U29938 ( .IN1(n1795), .IN2(n6893), .IN3(n1709), .IN4(n6894), .Q(n6883) );
  OA22X1 U29939 ( .IN1(n1967), .IN2(n6891), .IN3(n1881), .IN4(n6892), .Q(n6884) );
  OA22X1 U29940 ( .IN1(n2139), .IN2(n6889), .IN3(n2053), .IN4(n6890), .Q(n6885) );
  NAND4X0 U29941 ( .IN1(n6871), .IN2(n6872), .IN3(n6873), .IN4(n6874), .QN(
        s1_we_o) );
  OA22X1 U29942 ( .IN1(n1794), .IN2(n19769), .IN3(n1708), .IN4(n19763), .Q(
        n6871) );
  OA22X1 U29943 ( .IN1(n1966), .IN2(n19802), .IN3(n1880), .IN4(n19779), .Q(
        n6872) );
  OA22X1 U29944 ( .IN1(n2138), .IN2(n19835), .IN3(n2052), .IN4(n19828), .Q(
        n6873) );
  NAND4X0 U29945 ( .IN1(n6907), .IN2(n6908), .IN3(n6909), .IN4(n6910), .QN(
        s1_sel_o[0]) );
  OA22X1 U29946 ( .IN1(n1793), .IN2(n6881), .IN3(n1707), .IN4(n19761), .Q(
        n6907) );
  OA22X1 U29947 ( .IN1(n1965), .IN2(n19809), .IN3(n1879), .IN4(n19796), .Q(
        n6908) );
  OA22X1 U29948 ( .IN1(n2137), .IN2(n6877), .IN3(n2051), .IN4(n19829), .Q(
        n6909) );
  NAND4X0 U29949 ( .IN1(n6903), .IN2(n6904), .IN3(n6905), .IN4(n6906), .QN(
        s1_sel_o[1]) );
  OA22X1 U29950 ( .IN1(n1792), .IN2(n6881), .IN3(n1706), .IN4(n19761), .Q(
        n6903) );
  OA22X1 U29951 ( .IN1(n1964), .IN2(n19809), .IN3(n1878), .IN4(n19796), .Q(
        n6904) );
  OA22X1 U29952 ( .IN1(n2136), .IN2(n6877), .IN3(n2050), .IN4(n19829), .Q(
        n6905) );
  NAND4X0 U29953 ( .IN1(n6899), .IN2(n6900), .IN3(n6901), .IN4(n6902), .QN(
        s1_sel_o[2]) );
  OA22X1 U29954 ( .IN1(n1791), .IN2(n6881), .IN3(n1705), .IN4(n19763), .Q(
        n6899) );
  OA22X1 U29955 ( .IN1(n1963), .IN2(n19809), .IN3(n1877), .IN4(n19780), .Q(
        n6900) );
  OA22X1 U29956 ( .IN1(n2135), .IN2(n6877), .IN3(n2049), .IN4(n19813), .Q(
        n6901) );
  NAND4X0 U29957 ( .IN1(n6895), .IN2(n6896), .IN3(n6897), .IN4(n6898), .QN(
        s1_sel_o[3]) );
  OA22X1 U29958 ( .IN1(n1790), .IN2(n6881), .IN3(n1704), .IN4(n19763), .Q(
        n6895) );
  OA22X1 U29959 ( .IN1(n1962), .IN2(n19809), .IN3(n1876), .IN4(n19781), .Q(
        n6896) );
  OA22X1 U29960 ( .IN1(n2134), .IN2(n6877), .IN3(n2048), .IN4(n19811), .Q(
        n6897) );
  NAND4X0 U29961 ( .IN1(n7163), .IN2(n7164), .IN3(n7165), .IN4(n7166), .QN(
        s1_addr_o[0]) );
  OA22X1 U29962 ( .IN1(n1789), .IN2(n19769), .IN3(n1703), .IN4(n19746), .Q(
        n7163) );
  OA22X1 U29963 ( .IN1(n1961), .IN2(n19802), .IN3(n1875), .IN4(n19779), .Q(
        n7164) );
  OA22X1 U29964 ( .IN1(n2133), .IN2(n19835), .IN3(n2047), .IN4(n19825), .Q(
        n7165) );
  NAND4X0 U29965 ( .IN1(n7119), .IN2(n7120), .IN3(n7121), .IN4(n7122), .QN(
        s1_addr_o[1]) );
  OA22X1 U29966 ( .IN1(n1788), .IN2(n19771), .IN3(n1702), .IN4(n19749), .Q(
        n7119) );
  OA22X1 U29967 ( .IN1(n1960), .IN2(n19804), .IN3(n1874), .IN4(n19782), .Q(
        n7120) );
  OA22X1 U29968 ( .IN1(n2132), .IN2(n19837), .IN3(n2046), .IN4(n19813), .Q(
        n7121) );
  NAND4X0 U29969 ( .IN1(n7075), .IN2(n7076), .IN3(n7077), .IN4(n7078), .QN(
        s1_addr_o[2]) );
  OA22X1 U29970 ( .IN1(n1787), .IN2(n19769), .IN3(n1701), .IN4(n19753), .Q(
        n7075) );
  OA22X1 U29971 ( .IN1(n1959), .IN2(n19806), .IN3(n1873), .IN4(n19786), .Q(
        n7076) );
  OA22X1 U29972 ( .IN1(n2131), .IN2(n19839), .IN3(n2045), .IN4(n19817), .Q(
        n7077) );
  NAND4X0 U29973 ( .IN1(n7063), .IN2(n7064), .IN3(n7065), .IN4(n7066), .QN(
        s1_addr_o[3]) );
  OA22X1 U29974 ( .IN1(n1786), .IN2(n6881), .IN3(n1699), .IN4(n19754), .Q(
        n7063) );
  OA22X1 U29975 ( .IN1(n1958), .IN2(n19809), .IN3(n1872), .IN4(n19787), .Q(
        n7064) );
  OA22X1 U29976 ( .IN1(n2130), .IN2(n6877), .IN3(n2044), .IN4(n19818), .Q(
        n7065) );
  NAND4X0 U29977 ( .IN1(n7059), .IN2(n7060), .IN3(n7061), .IN4(n7062), .QN(
        s1_addr_o[4]) );
  OA22X1 U29978 ( .IN1(n1785), .IN2(n19772), .IN3(n1697), .IN4(n19754), .Q(
        n7059) );
  OA22X1 U29979 ( .IN1(n1957), .IN2(n19805), .IN3(n1871), .IN4(n19787), .Q(
        n7060) );
  OA22X1 U29980 ( .IN1(n2129), .IN2(n19838), .IN3(n2043), .IN4(n19818), .Q(
        n7061) );
  NAND4X0 U29981 ( .IN1(n7055), .IN2(n7056), .IN3(n7057), .IN4(n7058), .QN(
        s1_addr_o[5]) );
  OA22X1 U29982 ( .IN1(n1784), .IN2(n6881), .IN3(n1696), .IN4(n19755), .Q(
        n7055) );
  OA22X1 U29983 ( .IN1(n1956), .IN2(n19809), .IN3(n1870), .IN4(n19788), .Q(
        n7056) );
  OA22X1 U29984 ( .IN1(n2128), .IN2(n6877), .IN3(n2042), .IN4(n19819), .Q(
        n7057) );
  NAND4X0 U29985 ( .IN1(n7051), .IN2(n7052), .IN3(n7053), .IN4(n7054), .QN(
        s1_addr_o[6]) );
  OA22X1 U29986 ( .IN1(n1783), .IN2(n19773), .IN3(n1679), .IN4(n19755), .Q(
        n7051) );
  OA22X1 U29987 ( .IN1(n1955), .IN2(n19807), .IN3(n1869), .IN4(n19788), .Q(
        n7052) );
  OA22X1 U29988 ( .IN1(n2127), .IN2(n19840), .IN3(n2041), .IN4(n19819), .Q(
        n7053) );
  NAND4X0 U29989 ( .IN1(n7047), .IN2(n7048), .IN3(n7049), .IN4(n7050), .QN(
        s1_addr_o[7]) );
  OA22X1 U29990 ( .IN1(n1782), .IN2(n19773), .IN3(n1678), .IN4(n19755), .Q(
        n7047) );
  OA22X1 U29991 ( .IN1(n1954), .IN2(n19807), .IN3(n1868), .IN4(n19788), .Q(
        n7048) );
  OA22X1 U29992 ( .IN1(n2126), .IN2(n19840), .IN3(n2040), .IN4(n19819), .Q(
        n7049) );
  NAND4X0 U29993 ( .IN1(n7043), .IN2(n7044), .IN3(n7045), .IN4(n7046), .QN(
        s1_addr_o[8]) );
  OA22X1 U29994 ( .IN1(n1781), .IN2(n19773), .IN3(n1677), .IN4(n19756), .Q(
        n7043) );
  OA22X1 U29995 ( .IN1(n1953), .IN2(n19807), .IN3(n1867), .IN4(n19789), .Q(
        n7044) );
  OA22X1 U29996 ( .IN1(n2125), .IN2(n19840), .IN3(n2039), .IN4(n19820), .Q(
        n7045) );
  NAND4X0 U29997 ( .IN1(n7039), .IN2(n7040), .IN3(n7041), .IN4(n7042), .QN(
        s1_addr_o[9]) );
  OA22X1 U29998 ( .IN1(n1780), .IN2(n19773), .IN3(n1676), .IN4(n19756), .Q(
        n7039) );
  OA22X1 U29999 ( .IN1(n1952), .IN2(n19807), .IN3(n1866), .IN4(n19789), .Q(
        n7040) );
  OA22X1 U30000 ( .IN1(n2124), .IN2(n19840), .IN3(n2038), .IN4(n19820), .Q(
        n7041) );
  NAND4X0 U30001 ( .IN1(n7159), .IN2(n7160), .IN3(n7161), .IN4(n7162), .QN(
        s1_addr_o[10]) );
  OA22X1 U30002 ( .IN1(n1779), .IN2(n19769), .IN3(n1675), .IN4(n19746), .Q(
        n7159) );
  OA22X1 U30003 ( .IN1(n1951), .IN2(n19802), .IN3(n1865), .IN4(n19779), .Q(
        n7160) );
  OA22X1 U30004 ( .IN1(n2123), .IN2(n19835), .IN3(n2037), .IN4(n19828), .Q(
        n7161) );
  NAND4X0 U30005 ( .IN1(n7155), .IN2(n7156), .IN3(n7157), .IN4(n7158), .QN(
        s1_addr_o[11]) );
  OA22X1 U30006 ( .IN1(n1778), .IN2(n19769), .IN3(n1674), .IN4(n19746), .Q(
        n7155) );
  OA22X1 U30007 ( .IN1(n1950), .IN2(n19802), .IN3(n1864), .IN4(n19779), .Q(
        n7156) );
  OA22X1 U30008 ( .IN1(n2122), .IN2(n19835), .IN3(n2036), .IN4(n19823), .Q(
        n7157) );
  NAND4X0 U30009 ( .IN1(n7151), .IN2(n7152), .IN3(n7153), .IN4(n7154), .QN(
        s1_addr_o[12]) );
  OA22X1 U30010 ( .IN1(n1777), .IN2(n19769), .IN3(n1673), .IN4(n19747), .Q(
        n7151) );
  OA22X1 U30011 ( .IN1(n1949), .IN2(n19802), .IN3(n1863), .IN4(n19780), .Q(
        n7152) );
  OA22X1 U30012 ( .IN1(n2121), .IN2(n19835), .IN3(n2035), .IN4(n19812), .Q(
        n7153) );
  NAND4X0 U30013 ( .IN1(n7147), .IN2(n7148), .IN3(n7149), .IN4(n7150), .QN(
        s1_addr_o[13]) );
  OA22X1 U30014 ( .IN1(n1776), .IN2(n19770), .IN3(n1672), .IN4(n19747), .Q(
        n7147) );
  OA22X1 U30015 ( .IN1(n1948), .IN2(n19803), .IN3(n1862), .IN4(n19780), .Q(
        n7148) );
  OA22X1 U30016 ( .IN1(n2120), .IN2(n19836), .IN3(n2034), .IN4(n19812), .Q(
        n7149) );
  NAND4X0 U30017 ( .IN1(n7143), .IN2(n7144), .IN3(n7145), .IN4(n7146), .QN(
        s1_addr_o[14]) );
  OA22X1 U30018 ( .IN1(n1775), .IN2(n19770), .IN3(n1671), .IN4(n19747), .Q(
        n7143) );
  OA22X1 U30019 ( .IN1(n1947), .IN2(n19803), .IN3(n1861), .IN4(n19780), .Q(
        n7144) );
  OA22X1 U30020 ( .IN1(n2119), .IN2(n19836), .IN3(n2033), .IN4(n19812), .Q(
        n7145) );
  NAND4X0 U30021 ( .IN1(n7139), .IN2(n7140), .IN3(n7141), .IN4(n7142), .QN(
        s1_addr_o[15]) );
  OA22X1 U30022 ( .IN1(n1774), .IN2(n19770), .IN3(n1670), .IN4(n19748), .Q(
        n7139) );
  OA22X1 U30023 ( .IN1(n1946), .IN2(n19803), .IN3(n1860), .IN4(n19781), .Q(
        n7140) );
  OA22X1 U30024 ( .IN1(n2118), .IN2(n19836), .IN3(n2032), .IN4(n19823), .Q(
        n7141) );
  NAND4X0 U30025 ( .IN1(n7135), .IN2(n7136), .IN3(n7137), .IN4(n7138), .QN(
        s1_addr_o[16]) );
  OA22X1 U30026 ( .IN1(n1773), .IN2(n19770), .IN3(n1669), .IN4(n19748), .Q(
        n7135) );
  OA22X1 U30027 ( .IN1(n1945), .IN2(n19803), .IN3(n1859), .IN4(n19781), .Q(
        n7136) );
  OA22X1 U30028 ( .IN1(n2117), .IN2(n19836), .IN3(n2031), .IN4(n19812), .Q(
        n7137) );
  NAND4X0 U30029 ( .IN1(n7131), .IN2(n7132), .IN3(n7133), .IN4(n7134), .QN(
        s1_addr_o[17]) );
  OA22X1 U30030 ( .IN1(n1772), .IN2(n19771), .IN3(n1668), .IN4(n19748), .Q(
        n7131) );
  OA22X1 U30031 ( .IN1(n1944), .IN2(n19804), .IN3(n1858), .IN4(n19781), .Q(
        n7132) );
  OA22X1 U30032 ( .IN1(n2116), .IN2(n19837), .IN3(n2030), .IN4(n19824), .Q(
        n7133) );
  NAND4X0 U30033 ( .IN1(n7127), .IN2(n7128), .IN3(n7129), .IN4(n7130), .QN(
        s1_addr_o[18]) );
  OA22X1 U30034 ( .IN1(n1771), .IN2(n19771), .IN3(n1667), .IN4(n19749), .Q(
        n7127) );
  OA22X1 U30035 ( .IN1(n1943), .IN2(n19804), .IN3(n1857), .IN4(n19782), .Q(
        n7128) );
  OA22X1 U30036 ( .IN1(n2115), .IN2(n19837), .IN3(n2029), .IN4(n19813), .Q(
        n7129) );
  NAND4X0 U30037 ( .IN1(n7123), .IN2(n7124), .IN3(n7125), .IN4(n7126), .QN(
        s1_addr_o[19]) );
  OA22X1 U30038 ( .IN1(n1770), .IN2(n19771), .IN3(n1666), .IN4(n19749), .Q(
        n7123) );
  OA22X1 U30039 ( .IN1(n1942), .IN2(n19804), .IN3(n1856), .IN4(n19782), .Q(
        n7124) );
  OA22X1 U30040 ( .IN1(n2114), .IN2(n19837), .IN3(n2028), .IN4(n19813), .Q(
        n7125) );
  NAND4X0 U30041 ( .IN1(n7115), .IN2(n7116), .IN3(n7117), .IN4(n7118), .QN(
        s1_addr_o[20]) );
  OA22X1 U30042 ( .IN1(n1769), .IN2(n19770), .IN3(n1665), .IN4(n19750), .Q(
        n7115) );
  OA22X1 U30043 ( .IN1(n1941), .IN2(n19803), .IN3(n1855), .IN4(n19783), .Q(
        n7116) );
  OA22X1 U30044 ( .IN1(n2113), .IN2(n19836), .IN3(n2027), .IN4(n19814), .Q(
        n7117) );
  NAND4X0 U30045 ( .IN1(n7111), .IN2(n7112), .IN3(n7113), .IN4(n7114), .QN(
        s1_addr_o[21]) );
  OA22X1 U30046 ( .IN1(n1768), .IN2(n19770), .IN3(n1664), .IN4(n19750), .Q(
        n7111) );
  OA22X1 U30047 ( .IN1(n1940), .IN2(n19803), .IN3(n1854), .IN4(n19783), .Q(
        n7112) );
  OA22X1 U30048 ( .IN1(n2112), .IN2(n19836), .IN3(n2026), .IN4(n19814), .Q(
        n7113) );
  NAND4X0 U30049 ( .IN1(n7107), .IN2(n7108), .IN3(n7109), .IN4(n7110), .QN(
        s1_addr_o[22]) );
  OA22X1 U30050 ( .IN1(n1767), .IN2(n19769), .IN3(n1663), .IN4(n19750), .Q(
        n7107) );
  OA22X1 U30051 ( .IN1(n1939), .IN2(n19802), .IN3(n1853), .IN4(n19783), .Q(
        n7108) );
  OA22X1 U30052 ( .IN1(n2111), .IN2(n19835), .IN3(n2025), .IN4(n19814), .Q(
        n7109) );
  NAND4X0 U30053 ( .IN1(n7103), .IN2(n7104), .IN3(n7105), .IN4(n7106), .QN(
        s1_addr_o[23]) );
  OA22X1 U30054 ( .IN1(n1766), .IN2(n19770), .IN3(n1662), .IN4(n19751), .Q(
        n7103) );
  OA22X1 U30055 ( .IN1(n1938), .IN2(n19803), .IN3(n1852), .IN4(n19784), .Q(
        n7104) );
  OA22X1 U30056 ( .IN1(n2110), .IN2(n19836), .IN3(n2024), .IN4(n19815), .Q(
        n7105) );
  NAND4X0 U30057 ( .IN1(n7099), .IN2(n7100), .IN3(n7101), .IN4(n7102), .QN(
        s1_addr_o[24]) );
  OA22X1 U30058 ( .IN1(n1765), .IN2(n19772), .IN3(n1661), .IN4(n19751), .Q(
        n7099) );
  OA22X1 U30059 ( .IN1(n1937), .IN2(n19805), .IN3(n1851), .IN4(n19784), .Q(
        n7100) );
  OA22X1 U30060 ( .IN1(n2109), .IN2(n19838), .IN3(n2023), .IN4(n19815), .Q(
        n7101) );
  NAND4X0 U30061 ( .IN1(n7095), .IN2(n7096), .IN3(n7097), .IN4(n7098), .QN(
        s1_addr_o[25]) );
  OA22X1 U30062 ( .IN1(n1764), .IN2(n19772), .IN3(n1660), .IN4(n19751), .Q(
        n7095) );
  OA22X1 U30063 ( .IN1(n1936), .IN2(n19805), .IN3(n1850), .IN4(n19784), .Q(
        n7096) );
  OA22X1 U30064 ( .IN1(n2108), .IN2(n19838), .IN3(n2022), .IN4(n19815), .Q(
        n7097) );
  NAND4X0 U30065 ( .IN1(n7091), .IN2(n7092), .IN3(n7093), .IN4(n7094), .QN(
        s1_addr_o[26]) );
  OA22X1 U30066 ( .IN1(n1763), .IN2(n19772), .IN3(n1659), .IN4(n19752), .Q(
        n7091) );
  OA22X1 U30067 ( .IN1(n1935), .IN2(n19805), .IN3(n1849), .IN4(n19785), .Q(
        n7092) );
  OA22X1 U30068 ( .IN1(n2107), .IN2(n19838), .IN3(n2021), .IN4(n19816), .Q(
        n7093) );
  NAND4X0 U30069 ( .IN1(n7087), .IN2(n7088), .IN3(n7089), .IN4(n7090), .QN(
        s1_addr_o[27]) );
  OA22X1 U30070 ( .IN1(n1762), .IN2(n19772), .IN3(n1658), .IN4(n19752), .Q(
        n7087) );
  OA22X1 U30071 ( .IN1(n1934), .IN2(n19805), .IN3(n1848), .IN4(n19785), .Q(
        n7088) );
  OA22X1 U30072 ( .IN1(n2106), .IN2(n19838), .IN3(n2020), .IN4(n19816), .Q(
        n7089) );
  NAND4X0 U30073 ( .IN1(n7083), .IN2(n7084), .IN3(n7085), .IN4(n7086), .QN(
        s1_addr_o[28]) );
  OA22X1 U30074 ( .IN1(n1761), .IN2(n19773), .IN3(n1657), .IN4(n19752), .Q(
        n7083) );
  OA22X1 U30075 ( .IN1(n1933), .IN2(n19806), .IN3(n1847), .IN4(n19785), .Q(
        n7084) );
  OA22X1 U30076 ( .IN1(n2105), .IN2(n19839), .IN3(n2019), .IN4(n19816), .Q(
        n7085) );
  NAND4X0 U30077 ( .IN1(n7079), .IN2(n7080), .IN3(n7081), .IN4(n7082), .QN(
        s1_addr_o[29]) );
  OA22X1 U30078 ( .IN1(n1760), .IN2(n19772), .IN3(n1656), .IN4(n19753), .Q(
        n7079) );
  OA22X1 U30079 ( .IN1(n1932), .IN2(n19806), .IN3(n1846), .IN4(n19786), .Q(
        n7080) );
  OA22X1 U30080 ( .IN1(n2104), .IN2(n19839), .IN3(n2018), .IN4(n19817), .Q(
        n7081) );
  NAND4X0 U30081 ( .IN1(n7071), .IN2(n7072), .IN3(n7073), .IN4(n7074), .QN(
        s1_addr_o[30]) );
  OA22X1 U30082 ( .IN1(n1759), .IN2(n19772), .IN3(n1655), .IN4(n19753), .Q(
        n7071) );
  OA22X1 U30083 ( .IN1(n1931), .IN2(n19806), .IN3(n1845), .IN4(n19786), .Q(
        n7072) );
  OA22X1 U30084 ( .IN1(n2103), .IN2(n19839), .IN3(n2017), .IN4(n19817), .Q(
        n7073) );
  NAND4X0 U30085 ( .IN1(n7067), .IN2(n7068), .IN3(n7069), .IN4(n7070), .QN(
        s1_addr_o[31]) );
  OA22X1 U30086 ( .IN1(n1758), .IN2(n19773), .IN3(n1650), .IN4(n19754), .Q(
        n7067) );
  OA22X1 U30087 ( .IN1(n1930), .IN2(n19806), .IN3(n1844), .IN4(n19787), .Q(
        n7068) );
  OA22X1 U30088 ( .IN1(n2102), .IN2(n19839), .IN3(n2016), .IN4(n19818), .Q(
        n7069) );
  NAND4X0 U30089 ( .IN1(n7035), .IN2(n7036), .IN3(n7037), .IN4(n7038), .QN(
        s1_data_o[0]) );
  OA22X1 U30090 ( .IN1(n1741), .IN2(n19771), .IN3(n1636), .IN4(n19756), .Q(
        n7035) );
  OA22X1 U30091 ( .IN1(n1913), .IN2(n19804), .IN3(n1827), .IN4(n19789), .Q(
        n7036) );
  OA22X1 U30092 ( .IN1(n2085), .IN2(n19841), .IN3(n1999), .IN4(n19820), .Q(
        n7037) );
  NAND4X0 U30093 ( .IN1(n6991), .IN2(n6992), .IN3(n6993), .IN4(n6994), .QN(
        s1_data_o[1]) );
  OA22X1 U30094 ( .IN1(n1740), .IN2(n19775), .IN3(n1635), .IN4(n19758), .Q(
        n6991) );
  OA22X1 U30095 ( .IN1(n1912), .IN2(n19808), .IN3(n1826), .IN4(n19793), .Q(
        n6992) );
  OA22X1 U30096 ( .IN1(n2084), .IN2(n19837), .IN3(n1998), .IN4(n19821), .Q(
        n6993) );
  NAND4X0 U30097 ( .IN1(n6947), .IN2(n6948), .IN3(n6949), .IN4(n6950), .QN(
        s1_data_o[2]) );
  OA22X1 U30098 ( .IN1(n1739), .IN2(n19774), .IN3(n1634), .IN4(n19761), .Q(
        n6947) );
  OA22X1 U30099 ( .IN1(n1911), .IN2(n6879), .IN3(n1825), .IN4(n19796), .Q(
        n6948) );
  OA22X1 U30100 ( .IN1(n2083), .IN2(n19842), .IN3(n1997), .IN4(n19826), .Q(
        n6949) );
  NAND4X0 U30101 ( .IN1(n6935), .IN2(n6936), .IN3(n6937), .IN4(n6938), .QN(
        s1_data_o[3]) );
  OA22X1 U30102 ( .IN1(n1738), .IN2(n19771), .IN3(n1633), .IN4(n19761), .Q(
        n6935) );
  OA22X1 U30103 ( .IN1(n1910), .IN2(n6879), .IN3(n1824), .IN4(n19796), .Q(
        n6936) );
  OA22X1 U30104 ( .IN1(n2082), .IN2(n19842), .IN3(n1996), .IN4(n19827), .Q(
        n6937) );
  NAND4X0 U30105 ( .IN1(n6931), .IN2(n6932), .IN3(n6933), .IN4(n6934), .QN(
        s1_data_o[4]) );
  OA22X1 U30106 ( .IN1(n1737), .IN2(n19771), .IN3(n1632), .IN4(n19761), .Q(
        n6931) );
  OA22X1 U30107 ( .IN1(n1909), .IN2(n19805), .IN3(n1823), .IN4(n19796), .Q(
        n6932) );
  OA22X1 U30108 ( .IN1(n2081), .IN2(n19838), .IN3(n1995), .IN4(n19827), .Q(
        n6933) );
  NAND4X0 U30109 ( .IN1(n6927), .IN2(n6928), .IN3(n6929), .IN4(n6930), .QN(
        s1_data_o[5]) );
  OA22X1 U30110 ( .IN1(n1736), .IN2(n19774), .IN3(n1631), .IN4(n19761), .Q(
        n6927) );
  OA22X1 U30111 ( .IN1(n1908), .IN2(n6879), .IN3(n1822), .IN4(n19796), .Q(
        n6928) );
  OA22X1 U30112 ( .IN1(n2080), .IN2(n19840), .IN3(n1994), .IN4(n19827), .Q(
        n6929) );
  NAND4X0 U30113 ( .IN1(n6923), .IN2(n6924), .IN3(n6925), .IN4(n6926), .QN(
        s1_data_o[6]) );
  OA22X1 U30114 ( .IN1(n1735), .IN2(n19776), .IN3(n1630), .IN4(n19762), .Q(
        n6923) );
  OA22X1 U30115 ( .IN1(n1907), .IN2(n19808), .IN3(n1821), .IN4(n19794), .Q(
        n6924) );
  OA22X1 U30116 ( .IN1(n2079), .IN2(n19842), .IN3(n1993), .IN4(n19828), .Q(
        n6925) );
  NAND4X0 U30117 ( .IN1(n6919), .IN2(n6920), .IN3(n6921), .IN4(n6922), .QN(
        s1_data_o[7]) );
  OA22X1 U30118 ( .IN1(n1734), .IN2(n19776), .IN3(n1629), .IN4(n19762), .Q(
        n6919) );
  OA22X1 U30119 ( .IN1(n1906), .IN2(n19808), .IN3(n1820), .IN4(n19794), .Q(
        n6920) );
  OA22X1 U30120 ( .IN1(n2078), .IN2(n19842), .IN3(n1992), .IN4(n19828), .Q(
        n6921) );
  NAND4X0 U30121 ( .IN1(n6915), .IN2(n6916), .IN3(n6917), .IN4(n6918), .QN(
        s1_data_o[8]) );
  OA22X1 U30122 ( .IN1(n1733), .IN2(n19776), .IN3(n1628), .IN4(n19762), .Q(
        n6915) );
  OA22X1 U30123 ( .IN1(n1905), .IN2(n19808), .IN3(n1819), .IN4(n19794), .Q(
        n6916) );
  OA22X1 U30124 ( .IN1(n2077), .IN2(n19842), .IN3(n1991), .IN4(n19828), .Q(
        n6917) );
  NAND4X0 U30125 ( .IN1(n6911), .IN2(n6912), .IN3(n6913), .IN4(n6914), .QN(
        s1_data_o[9]) );
  OA22X1 U30126 ( .IN1(n1732), .IN2(n19776), .IN3(n1627), .IN4(n19761), .Q(
        n6911) );
  OA22X1 U30127 ( .IN1(n1904), .IN2(n19808), .IN3(n1818), .IN4(n19794), .Q(
        n6912) );
  OA22X1 U30128 ( .IN1(n2076), .IN2(n19842), .IN3(n1990), .IN4(n19829), .Q(
        n6913) );
  NAND4X0 U30129 ( .IN1(n7031), .IN2(n7032), .IN3(n7033), .IN4(n7034), .QN(
        s1_data_o[10]) );
  OA22X1 U30130 ( .IN1(n1731), .IN2(n19776), .IN3(n1626), .IN4(n19757), .Q(
        n7031) );
  OA22X1 U30131 ( .IN1(n1903), .IN2(n19802), .IN3(n1817), .IN4(n19790), .Q(
        n7032) );
  OA22X1 U30132 ( .IN1(n2075), .IN2(n19841), .IN3(n1989), .IN4(n19814), .Q(
        n7033) );
  NAND4X0 U30133 ( .IN1(n7027), .IN2(n7028), .IN3(n7029), .IN4(n7030), .QN(
        s1_data_o[11]) );
  OA22X1 U30134 ( .IN1(n1730), .IN2(n19774), .IN3(n1625), .IN4(n19757), .Q(
        n7027) );
  OA22X1 U30135 ( .IN1(n1902), .IN2(n19809), .IN3(n1816), .IN4(n19790), .Q(
        n7028) );
  OA22X1 U30136 ( .IN1(n2074), .IN2(n19841), .IN3(n1988), .IN4(n19820), .Q(
        n7029) );
  NAND4X0 U30137 ( .IN1(n7023), .IN2(n7024), .IN3(n7025), .IN4(n7026), .QN(
        s1_data_o[12]) );
  OA22X1 U30138 ( .IN1(n1729), .IN2(n19775), .IN3(n1624), .IN4(n19757), .Q(
        n7023) );
  OA22X1 U30139 ( .IN1(n1901), .IN2(n19805), .IN3(n1815), .IN4(n19790), .Q(
        n7024) );
  OA22X1 U30140 ( .IN1(n2073), .IN2(n19841), .IN3(n1987), .IN4(n19814), .Q(
        n7025) );
  NAND4X0 U30141 ( .IN1(n7019), .IN2(n7020), .IN3(n7021), .IN4(n7022), .QN(
        s1_data_o[13]) );
  OA22X1 U30142 ( .IN1(n1728), .IN2(n19774), .IN3(n1623), .IN4(n19758), .Q(
        n7019) );
  OA22X1 U30143 ( .IN1(n1900), .IN2(n19806), .IN3(n1814), .IN4(n19791), .Q(
        n7020) );
  OA22X1 U30144 ( .IN1(n2072), .IN2(n19839), .IN3(n1986), .IN4(n19821), .Q(
        n7021) );
  NAND4X0 U30145 ( .IN1(n7015), .IN2(n7016), .IN3(n7017), .IN4(n7018), .QN(
        s1_data_o[14]) );
  OA22X1 U30146 ( .IN1(n1727), .IN2(n19774), .IN3(n1622), .IN4(n19758), .Q(
        n7015) );
  OA22X1 U30147 ( .IN1(n1899), .IN2(n19805), .IN3(n1813), .IN4(n19791), .Q(
        n7016) );
  OA22X1 U30148 ( .IN1(n2071), .IN2(n19838), .IN3(n1985), .IN4(n19821), .Q(
        n7017) );
  NAND4X0 U30149 ( .IN1(n7011), .IN2(n7012), .IN3(n7013), .IN4(n7014), .QN(
        s1_data_o[15]) );
  OA22X1 U30150 ( .IN1(n1726), .IN2(n19774), .IN3(n1621), .IN4(n19758), .Q(
        n7011) );
  OA22X1 U30151 ( .IN1(n1898), .IN2(n19806), .IN3(n1812), .IN4(n19791), .Q(
        n7012) );
  OA22X1 U30152 ( .IN1(n2070), .IN2(n19839), .IN3(n1984), .IN4(n19821), .Q(
        n7013) );
  NAND4X0 U30153 ( .IN1(n7007), .IN2(n7008), .IN3(n7009), .IN4(n7010), .QN(
        s1_data_o[16]) );
  OA22X1 U30154 ( .IN1(n1725), .IN2(n19774), .IN3(n1620), .IN4(n19759), .Q(
        n7007) );
  OA22X1 U30155 ( .IN1(n1897), .IN2(n19802), .IN3(n1811), .IN4(n19792), .Q(
        n7008) );
  OA22X1 U30156 ( .IN1(n2069), .IN2(n19835), .IN3(n1983), .IN4(n19822), .Q(
        n7009) );
  NAND4X0 U30157 ( .IN1(n7003), .IN2(n7004), .IN3(n7005), .IN4(n7006), .QN(
        s1_data_o[17]) );
  OA22X1 U30158 ( .IN1(n1724), .IN2(n19775), .IN3(n1619), .IN4(n19759), .Q(
        n7003) );
  OA22X1 U30159 ( .IN1(n1896), .IN2(n19807), .IN3(n1810), .IN4(n19792), .Q(
        n7004) );
  OA22X1 U30160 ( .IN1(n2068), .IN2(n19841), .IN3(n1982), .IN4(n19822), .Q(
        n7005) );
  NAND4X0 U30161 ( .IN1(n6999), .IN2(n7000), .IN3(n7001), .IN4(n7002), .QN(
        s1_data_o[18]) );
  OA22X1 U30162 ( .IN1(n1723), .IN2(n19775), .IN3(n1618), .IN4(n19759), .Q(
        n6999) );
  OA22X1 U30163 ( .IN1(n1895), .IN2(n19804), .IN3(n1809), .IN4(n19792), .Q(
        n7000) );
  OA22X1 U30164 ( .IN1(n2067), .IN2(n19835), .IN3(n1981), .IN4(n19822), .Q(
        n7001) );
  NAND4X0 U30165 ( .IN1(n6995), .IN2(n6996), .IN3(n6997), .IN4(n6998), .QN(
        s1_data_o[19]) );
  OA22X1 U30166 ( .IN1(n1722), .IN2(n19775), .IN3(n1617), .IN4(n19759), .Q(
        n6995) );
  OA22X1 U30167 ( .IN1(n1894), .IN2(n19808), .IN3(n1808), .IN4(n19793), .Q(
        n6996) );
  OA22X1 U30168 ( .IN1(n2066), .IN2(n19838), .IN3(n1980), .IN4(n19822), .Q(
        n6997) );
  NAND4X0 U30169 ( .IN1(n6987), .IN2(n6988), .IN3(n6989), .IN4(n6990), .QN(
        s1_data_o[20]) );
  OA22X1 U30170 ( .IN1(n1721), .IN2(n19776), .IN3(n1616), .IN4(n19758), .Q(
        n6987) );
  OA22X1 U30171 ( .IN1(n1893), .IN2(n19808), .IN3(n1807), .IN4(n19793), .Q(
        n6988) );
  OA22X1 U30172 ( .IN1(n2065), .IN2(n19842), .IN3(n1979), .IN4(n19821), .Q(
        n6989) );
  NAND4X0 U30173 ( .IN1(n6983), .IN2(n6984), .IN3(n6985), .IN4(n6986), .QN(
        s1_data_o[21]) );
  OA22X1 U30174 ( .IN1(n1720), .IN2(n19770), .IN3(n1615), .IN4(n19761), .Q(
        n6983) );
  OA22X1 U30175 ( .IN1(n1892), .IN2(n19807), .IN3(n1806), .IN4(n19794), .Q(
        n6984) );
  OA22X1 U30176 ( .IN1(n2064), .IN2(n19840), .IN3(n1978), .IN4(n19823), .Q(
        n6985) );
  NAND4X0 U30177 ( .IN1(n6979), .IN2(n6980), .IN3(n6981), .IN4(n6982), .QN(
        s1_data_o[22]) );
  OA22X1 U30178 ( .IN1(n1719), .IN2(n19774), .IN3(n1614), .IN4(n19745), .Q(
        n6979) );
  OA22X1 U30179 ( .IN1(n1891), .IN2(n19804), .IN3(n1805), .IN4(n19794), .Q(
        n6980) );
  OA22X1 U30180 ( .IN1(n2063), .IN2(n19837), .IN3(n1977), .IN4(n19823), .Q(
        n6981) );
  NAND4X0 U30181 ( .IN1(n6975), .IN2(n6976), .IN3(n6977), .IN4(n6978), .QN(
        s1_data_o[23]) );
  OA22X1 U30182 ( .IN1(n1718), .IN2(n19775), .IN3(n1613), .IN4(n19763), .Q(
        n6975) );
  OA22X1 U30183 ( .IN1(n1890), .IN2(n19803), .IN3(n1804), .IN4(n19794), .Q(
        n6976) );
  OA22X1 U30184 ( .IN1(n2062), .IN2(n19841), .IN3(n1976), .IN4(n19823), .Q(
        n6977) );
  NAND4X0 U30185 ( .IN1(n6971), .IN2(n6972), .IN3(n6973), .IN4(n6974), .QN(
        s1_data_o[24]) );
  OA22X1 U30186 ( .IN1(n1717), .IN2(n19776), .IN3(n1612), .IN4(n19760), .Q(
        n6971) );
  OA22X1 U30187 ( .IN1(n1889), .IN2(n19808), .IN3(n1803), .IN4(n19795), .Q(
        n6972) );
  OA22X1 U30188 ( .IN1(n2061), .IN2(n19842), .IN3(n1975), .IN4(n19824), .Q(
        n6973) );
  NAND4X0 U30189 ( .IN1(n6967), .IN2(n6968), .IN3(n6969), .IN4(n6970), .QN(
        s1_data_o[25]) );
  OA22X1 U30190 ( .IN1(n1716), .IN2(n19773), .IN3(n1611), .IN4(n19760), .Q(
        n6967) );
  OA22X1 U30191 ( .IN1(n1888), .IN2(n19807), .IN3(n1802), .IN4(n19795), .Q(
        n6968) );
  OA22X1 U30192 ( .IN1(n2060), .IN2(n19840), .IN3(n1974), .IN4(n19824), .Q(
        n6969) );
  NAND4X0 U30193 ( .IN1(n6963), .IN2(n6964), .IN3(n6965), .IN4(n6966), .QN(
        s1_data_o[26]) );
  OA22X1 U30194 ( .IN1(n1715), .IN2(n19771), .IN3(n1610), .IN4(n19760), .Q(
        n6963) );
  OA22X1 U30195 ( .IN1(n1887), .IN2(n19804), .IN3(n1801), .IN4(n19795), .Q(
        n6964) );
  OA22X1 U30196 ( .IN1(n2059), .IN2(n19837), .IN3(n1973), .IN4(n19824), .Q(
        n6965) );
  NAND4X0 U30197 ( .IN1(n6959), .IN2(n6960), .IN3(n6961), .IN4(n6962), .QN(
        s1_data_o[27]) );
  OA22X1 U30198 ( .IN1(n1714), .IN2(n19776), .IN3(n1609), .IN4(n19763), .Q(
        n6959) );
  OA22X1 U30199 ( .IN1(n1886), .IN2(n19807), .IN3(n1800), .IN4(n19794), .Q(
        n6960) );
  OA22X1 U30200 ( .IN1(n2058), .IN2(n19841), .IN3(n1972), .IN4(n19825), .Q(
        n6961) );
  NAND4X0 U30201 ( .IN1(n6955), .IN2(n6956), .IN3(n6957), .IN4(n6958), .QN(
        s1_data_o[28]) );
  OA22X1 U30202 ( .IN1(n1713), .IN2(n19775), .IN3(n1608), .IN4(n19760), .Q(
        n6955) );
  OA22X1 U30203 ( .IN1(n1885), .IN2(n6879), .IN3(n1799), .IN4(n19795), .Q(
        n6956) );
  OA22X1 U30204 ( .IN1(n2057), .IN2(n19840), .IN3(n1971), .IN4(n19825), .Q(
        n6957) );
  NAND4X0 U30205 ( .IN1(n6951), .IN2(n6952), .IN3(n6953), .IN4(n6954), .QN(
        s1_data_o[29]) );
  OA22X1 U30206 ( .IN1(n1712), .IN2(n19769), .IN3(n1607), .IN4(n19762), .Q(
        n6951) );
  OA22X1 U30207 ( .IN1(n1884), .IN2(n6879), .IN3(n1798), .IN4(n19794), .Q(
        n6952) );
  OA22X1 U30208 ( .IN1(n2056), .IN2(n19837), .IN3(n1970), .IN4(n19825), .Q(
        n6953) );
  NAND4X0 U30209 ( .IN1(n6943), .IN2(n6944), .IN3(n6945), .IN4(n6946), .QN(
        s1_data_o[30]) );
  OA22X1 U30210 ( .IN1(n1711), .IN2(n6881), .IN3(n1606), .IN4(n19761), .Q(
        n6943) );
  OA22X1 U30211 ( .IN1(n1883), .IN2(n6879), .IN3(n1797), .IN4(n19796), .Q(
        n6944) );
  OA22X1 U30212 ( .IN1(n2055), .IN2(n19841), .IN3(n1969), .IN4(n19826), .Q(
        n6945) );
  NAND4X0 U30213 ( .IN1(n6939), .IN2(n6940), .IN3(n6941), .IN4(n6942), .QN(
        s1_data_o[31]) );
  OA22X1 U30214 ( .IN1(n1710), .IN2(n19775), .IN3(n1605), .IN4(n19761), .Q(
        n6939) );
  OA22X1 U30215 ( .IN1(n1882), .IN2(n19809), .IN3(n1796), .IN4(n19796), .Q(
        n6940) );
  OA22X1 U30216 ( .IN1(n2054), .IN2(n19836), .IN3(n1968), .IN4(n19826), .Q(
        n6941) );
  NAND4X0 U30217 ( .IN1(n8843), .IN2(n8844), .IN3(n8845), .IN4(n8846), .QN(
        s0_stb_o) );
  OA22X1 U30218 ( .IN1(n1795), .IN2(n8853), .IN3(n1709), .IN4(n8854), .Q(n8843) );
  OA22X1 U30219 ( .IN1(n1967), .IN2(n8851), .IN3(n1881), .IN4(n8852), .Q(n8844) );
  OA22X1 U30220 ( .IN1(n2139), .IN2(n8849), .IN3(n2053), .IN4(n8850), .Q(n8845) );
  NAND4X0 U30221 ( .IN1(n8831), .IN2(n8832), .IN3(n8833), .IN4(n8834), .QN(
        s0_we_o) );
  OA22X1 U30222 ( .IN1(n1794), .IN2(n18845), .IN3(n1708), .IN4(n18839), .Q(
        n8831) );
  OA22X1 U30223 ( .IN1(n1966), .IN2(n18878), .IN3(n1880), .IN4(n18855), .Q(
        n8832) );
  OA22X1 U30224 ( .IN1(n2138), .IN2(n18911), .IN3(n2052), .IN4(n18904), .Q(
        n8833) );
  NAND4X0 U30225 ( .IN1(n8867), .IN2(n8868), .IN3(n8869), .IN4(n8870), .QN(
        s0_sel_o[0]) );
  OA22X1 U30226 ( .IN1(n1793), .IN2(n8841), .IN3(n1707), .IN4(n18837), .Q(
        n8867) );
  OA22X1 U30227 ( .IN1(n1965), .IN2(n18885), .IN3(n1879), .IN4(n18872), .Q(
        n8868) );
  OA22X1 U30228 ( .IN1(n2137), .IN2(n8837), .IN3(n2051), .IN4(n18905), .Q(
        n8869) );
  NAND4X0 U30229 ( .IN1(n8863), .IN2(n8864), .IN3(n8865), .IN4(n8866), .QN(
        s0_sel_o[1]) );
  OA22X1 U30230 ( .IN1(n1792), .IN2(n8841), .IN3(n1706), .IN4(n18837), .Q(
        n8863) );
  OA22X1 U30231 ( .IN1(n1964), .IN2(n18885), .IN3(n1878), .IN4(n18872), .Q(
        n8864) );
  OA22X1 U30232 ( .IN1(n2136), .IN2(n8837), .IN3(n2050), .IN4(n18905), .Q(
        n8865) );
  NAND4X0 U30233 ( .IN1(n8859), .IN2(n8860), .IN3(n8861), .IN4(n8862), .QN(
        s0_sel_o[2]) );
  OA22X1 U30234 ( .IN1(n1791), .IN2(n8841), .IN3(n1705), .IN4(n18839), .Q(
        n8859) );
  OA22X1 U30235 ( .IN1(n1963), .IN2(n18885), .IN3(n1877), .IN4(n18856), .Q(
        n8860) );
  OA22X1 U30236 ( .IN1(n2135), .IN2(n8837), .IN3(n2049), .IN4(n18889), .Q(
        n8861) );
  NAND4X0 U30237 ( .IN1(n8855), .IN2(n8856), .IN3(n8857), .IN4(n8858), .QN(
        s0_sel_o[3]) );
  OA22X1 U30238 ( .IN1(n1790), .IN2(n8841), .IN3(n1704), .IN4(n18839), .Q(
        n8855) );
  OA22X1 U30239 ( .IN1(n1962), .IN2(n18885), .IN3(n1876), .IN4(n18857), .Q(
        n8856) );
  OA22X1 U30240 ( .IN1(n2134), .IN2(n8837), .IN3(n2048), .IN4(n18887), .Q(
        n8857) );
  NAND4X0 U30241 ( .IN1(n9123), .IN2(n9124), .IN3(n9125), .IN4(n9126), .QN(
        s0_addr_o[0]) );
  OA22X1 U30242 ( .IN1(n1789), .IN2(n18845), .IN3(n1703), .IN4(n18822), .Q(
        n9123) );
  OA22X1 U30243 ( .IN1(n1961), .IN2(n18878), .IN3(n1875), .IN4(n18855), .Q(
        n9124) );
  OA22X1 U30244 ( .IN1(n2133), .IN2(n18911), .IN3(n2047), .IN4(n18901), .Q(
        n9125) );
  NAND4X0 U30245 ( .IN1(n9079), .IN2(n9080), .IN3(n9081), .IN4(n9082), .QN(
        s0_addr_o[1]) );
  OA22X1 U30246 ( .IN1(n1788), .IN2(n18847), .IN3(n1702), .IN4(n18825), .Q(
        n9079) );
  OA22X1 U30247 ( .IN1(n1960), .IN2(n18880), .IN3(n1874), .IN4(n18858), .Q(
        n9080) );
  OA22X1 U30248 ( .IN1(n2132), .IN2(n18913), .IN3(n2046), .IN4(n18889), .Q(
        n9081) );
  NAND4X0 U30249 ( .IN1(n9035), .IN2(n9036), .IN3(n9037), .IN4(n9038), .QN(
        s0_addr_o[2]) );
  OA22X1 U30250 ( .IN1(n1787), .IN2(n18845), .IN3(n1701), .IN4(n18829), .Q(
        n9035) );
  OA22X1 U30251 ( .IN1(n1959), .IN2(n18882), .IN3(n1873), .IN4(n18862), .Q(
        n9036) );
  OA22X1 U30252 ( .IN1(n2131), .IN2(n18915), .IN3(n2045), .IN4(n18893), .Q(
        n9037) );
  NAND4X0 U30253 ( .IN1(n9023), .IN2(n9024), .IN3(n9025), .IN4(n9026), .QN(
        s0_addr_o[3]) );
  OA22X1 U30254 ( .IN1(n1786), .IN2(n8841), .IN3(n1699), .IN4(n18830), .Q(
        n9023) );
  OA22X1 U30255 ( .IN1(n1958), .IN2(n18885), .IN3(n1872), .IN4(n18863), .Q(
        n9024) );
  OA22X1 U30256 ( .IN1(n2130), .IN2(n8837), .IN3(n2044), .IN4(n18894), .Q(
        n9025) );
  NAND4X0 U30257 ( .IN1(n9019), .IN2(n9020), .IN3(n9021), .IN4(n9022), .QN(
        s0_addr_o[4]) );
  OA22X1 U30258 ( .IN1(n1785), .IN2(n18848), .IN3(n1697), .IN4(n18830), .Q(
        n9019) );
  OA22X1 U30259 ( .IN1(n1957), .IN2(n18881), .IN3(n1871), .IN4(n18863), .Q(
        n9020) );
  OA22X1 U30260 ( .IN1(n2129), .IN2(n18914), .IN3(n2043), .IN4(n18894), .Q(
        n9021) );
  NAND4X0 U30261 ( .IN1(n9015), .IN2(n9016), .IN3(n9017), .IN4(n9018), .QN(
        s0_addr_o[5]) );
  OA22X1 U30262 ( .IN1(n1784), .IN2(n8841), .IN3(n1696), .IN4(n18831), .Q(
        n9015) );
  OA22X1 U30263 ( .IN1(n1956), .IN2(n18885), .IN3(n1870), .IN4(n18864), .Q(
        n9016) );
  OA22X1 U30264 ( .IN1(n2128), .IN2(n8837), .IN3(n2042), .IN4(n18895), .Q(
        n9017) );
  NAND4X0 U30265 ( .IN1(n9011), .IN2(n9012), .IN3(n9013), .IN4(n9014), .QN(
        s0_addr_o[6]) );
  OA22X1 U30266 ( .IN1(n1783), .IN2(n18849), .IN3(n1679), .IN4(n18831), .Q(
        n9011) );
  OA22X1 U30267 ( .IN1(n1955), .IN2(n18883), .IN3(n1869), .IN4(n18864), .Q(
        n9012) );
  OA22X1 U30268 ( .IN1(n2127), .IN2(n18916), .IN3(n2041), .IN4(n18895), .Q(
        n9013) );
  NAND4X0 U30269 ( .IN1(n9007), .IN2(n9008), .IN3(n9009), .IN4(n9010), .QN(
        s0_addr_o[7]) );
  OA22X1 U30270 ( .IN1(n1782), .IN2(n18849), .IN3(n1678), .IN4(n18831), .Q(
        n9007) );
  OA22X1 U30271 ( .IN1(n1954), .IN2(n18883), .IN3(n1868), .IN4(n18864), .Q(
        n9008) );
  OA22X1 U30272 ( .IN1(n2126), .IN2(n18916), .IN3(n2040), .IN4(n18895), .Q(
        n9009) );
  NAND4X0 U30273 ( .IN1(n9003), .IN2(n9004), .IN3(n9005), .IN4(n9006), .QN(
        s0_addr_o[8]) );
  OA22X1 U30274 ( .IN1(n1781), .IN2(n18849), .IN3(n1677), .IN4(n18832), .Q(
        n9003) );
  OA22X1 U30275 ( .IN1(n1953), .IN2(n18883), .IN3(n1867), .IN4(n18865), .Q(
        n9004) );
  OA22X1 U30276 ( .IN1(n2125), .IN2(n18916), .IN3(n2039), .IN4(n18896), .Q(
        n9005) );
  NAND4X0 U30277 ( .IN1(n8999), .IN2(n9000), .IN3(n9001), .IN4(n9002), .QN(
        s0_addr_o[9]) );
  OA22X1 U30278 ( .IN1(n1780), .IN2(n18849), .IN3(n1676), .IN4(n18832), .Q(
        n8999) );
  OA22X1 U30279 ( .IN1(n1952), .IN2(n18883), .IN3(n1866), .IN4(n18865), .Q(
        n9000) );
  OA22X1 U30280 ( .IN1(n2124), .IN2(n18916), .IN3(n2038), .IN4(n18896), .Q(
        n9001) );
  NAND4X0 U30281 ( .IN1(n9119), .IN2(n9120), .IN3(n9121), .IN4(n9122), .QN(
        s0_addr_o[10]) );
  OA22X1 U30282 ( .IN1(n1779), .IN2(n18845), .IN3(n1675), .IN4(n18822), .Q(
        n9119) );
  OA22X1 U30283 ( .IN1(n1951), .IN2(n18878), .IN3(n1865), .IN4(n18855), .Q(
        n9120) );
  OA22X1 U30284 ( .IN1(n2123), .IN2(n18911), .IN3(n2037), .IN4(n18904), .Q(
        n9121) );
  NAND4X0 U30285 ( .IN1(n9115), .IN2(n9116), .IN3(n9117), .IN4(n9118), .QN(
        s0_addr_o[11]) );
  OA22X1 U30286 ( .IN1(n1778), .IN2(n18845), .IN3(n1674), .IN4(n18822), .Q(
        n9115) );
  OA22X1 U30287 ( .IN1(n1950), .IN2(n18878), .IN3(n1864), .IN4(n18855), .Q(
        n9116) );
  OA22X1 U30288 ( .IN1(n2122), .IN2(n18911), .IN3(n2036), .IN4(n18899), .Q(
        n9117) );
  NAND4X0 U30289 ( .IN1(n9111), .IN2(n9112), .IN3(n9113), .IN4(n9114), .QN(
        s0_addr_o[12]) );
  OA22X1 U30290 ( .IN1(n1777), .IN2(n18845), .IN3(n1673), .IN4(n18823), .Q(
        n9111) );
  OA22X1 U30291 ( .IN1(n1949), .IN2(n18878), .IN3(n1863), .IN4(n18856), .Q(
        n9112) );
  OA22X1 U30292 ( .IN1(n2121), .IN2(n18911), .IN3(n2035), .IN4(n18888), .Q(
        n9113) );
  NAND4X0 U30293 ( .IN1(n9107), .IN2(n9108), .IN3(n9109), .IN4(n9110), .QN(
        s0_addr_o[13]) );
  OA22X1 U30294 ( .IN1(n1776), .IN2(n18846), .IN3(n1672), .IN4(n18823), .Q(
        n9107) );
  OA22X1 U30295 ( .IN1(n1948), .IN2(n18879), .IN3(n1862), .IN4(n18856), .Q(
        n9108) );
  OA22X1 U30296 ( .IN1(n2120), .IN2(n18912), .IN3(n2034), .IN4(n18888), .Q(
        n9109) );
  NAND4X0 U30297 ( .IN1(n9103), .IN2(n9104), .IN3(n9105), .IN4(n9106), .QN(
        s0_addr_o[14]) );
  OA22X1 U30298 ( .IN1(n1775), .IN2(n18846), .IN3(n1671), .IN4(n18823), .Q(
        n9103) );
  OA22X1 U30299 ( .IN1(n1947), .IN2(n18879), .IN3(n1861), .IN4(n18856), .Q(
        n9104) );
  OA22X1 U30300 ( .IN1(n2119), .IN2(n18912), .IN3(n2033), .IN4(n18888), .Q(
        n9105) );
  NAND4X0 U30301 ( .IN1(n9099), .IN2(n9100), .IN3(n9101), .IN4(n9102), .QN(
        s0_addr_o[15]) );
  OA22X1 U30302 ( .IN1(n1774), .IN2(n18846), .IN3(n1670), .IN4(n18824), .Q(
        n9099) );
  OA22X1 U30303 ( .IN1(n1946), .IN2(n18879), .IN3(n1860), .IN4(n18857), .Q(
        n9100) );
  OA22X1 U30304 ( .IN1(n2118), .IN2(n18912), .IN3(n2032), .IN4(n18899), .Q(
        n9101) );
  NAND4X0 U30305 ( .IN1(n9095), .IN2(n9096), .IN3(n9097), .IN4(n9098), .QN(
        s0_addr_o[16]) );
  OA22X1 U30306 ( .IN1(n1773), .IN2(n18846), .IN3(n1669), .IN4(n18824), .Q(
        n9095) );
  OA22X1 U30307 ( .IN1(n1945), .IN2(n18879), .IN3(n1859), .IN4(n18857), .Q(
        n9096) );
  OA22X1 U30308 ( .IN1(n2117), .IN2(n18912), .IN3(n2031), .IN4(n18888), .Q(
        n9097) );
  NAND4X0 U30309 ( .IN1(n9091), .IN2(n9092), .IN3(n9093), .IN4(n9094), .QN(
        s0_addr_o[17]) );
  OA22X1 U30310 ( .IN1(n1772), .IN2(n18847), .IN3(n1668), .IN4(n18824), .Q(
        n9091) );
  OA22X1 U30311 ( .IN1(n1944), .IN2(n18880), .IN3(n1858), .IN4(n18857), .Q(
        n9092) );
  OA22X1 U30312 ( .IN1(n2116), .IN2(n18913), .IN3(n2030), .IN4(n18900), .Q(
        n9093) );
  NAND4X0 U30313 ( .IN1(n9087), .IN2(n9088), .IN3(n9089), .IN4(n9090), .QN(
        s0_addr_o[18]) );
  OA22X1 U30314 ( .IN1(n1771), .IN2(n18847), .IN3(n1667), .IN4(n18825), .Q(
        n9087) );
  OA22X1 U30315 ( .IN1(n1943), .IN2(n18880), .IN3(n1857), .IN4(n18858), .Q(
        n9088) );
  OA22X1 U30316 ( .IN1(n2115), .IN2(n18913), .IN3(n2029), .IN4(n18889), .Q(
        n9089) );
  NAND4X0 U30317 ( .IN1(n9083), .IN2(n9084), .IN3(n9085), .IN4(n9086), .QN(
        s0_addr_o[19]) );
  OA22X1 U30318 ( .IN1(n1770), .IN2(n18847), .IN3(n1666), .IN4(n18825), .Q(
        n9083) );
  OA22X1 U30319 ( .IN1(n1942), .IN2(n18880), .IN3(n1856), .IN4(n18858), .Q(
        n9084) );
  OA22X1 U30320 ( .IN1(n2114), .IN2(n18913), .IN3(n2028), .IN4(n18889), .Q(
        n9085) );
  NAND4X0 U30321 ( .IN1(n9075), .IN2(n9076), .IN3(n9077), .IN4(n9078), .QN(
        s0_addr_o[20]) );
  OA22X1 U30322 ( .IN1(n1769), .IN2(n18846), .IN3(n1665), .IN4(n18826), .Q(
        n9075) );
  OA22X1 U30323 ( .IN1(n1941), .IN2(n18879), .IN3(n1855), .IN4(n18859), .Q(
        n9076) );
  OA22X1 U30324 ( .IN1(n2113), .IN2(n18912), .IN3(n2027), .IN4(n18890), .Q(
        n9077) );
  NAND4X0 U30325 ( .IN1(n9071), .IN2(n9072), .IN3(n9073), .IN4(n9074), .QN(
        s0_addr_o[21]) );
  OA22X1 U30326 ( .IN1(n1768), .IN2(n18846), .IN3(n1664), .IN4(n18826), .Q(
        n9071) );
  OA22X1 U30327 ( .IN1(n1940), .IN2(n18879), .IN3(n1854), .IN4(n18859), .Q(
        n9072) );
  OA22X1 U30328 ( .IN1(n2112), .IN2(n18912), .IN3(n2026), .IN4(n18890), .Q(
        n9073) );
  NAND4X0 U30329 ( .IN1(n9067), .IN2(n9068), .IN3(n9069), .IN4(n9070), .QN(
        s0_addr_o[22]) );
  OA22X1 U30330 ( .IN1(n1767), .IN2(n18845), .IN3(n1663), .IN4(n18826), .Q(
        n9067) );
  OA22X1 U30331 ( .IN1(n1939), .IN2(n18878), .IN3(n1853), .IN4(n18859), .Q(
        n9068) );
  OA22X1 U30332 ( .IN1(n2111), .IN2(n18911), .IN3(n2025), .IN4(n18890), .Q(
        n9069) );
  NAND4X0 U30333 ( .IN1(n9063), .IN2(n9064), .IN3(n9065), .IN4(n9066), .QN(
        s0_addr_o[23]) );
  OA22X1 U30334 ( .IN1(n1766), .IN2(n18846), .IN3(n1662), .IN4(n18827), .Q(
        n9063) );
  OA22X1 U30335 ( .IN1(n1938), .IN2(n18879), .IN3(n1852), .IN4(n18860), .Q(
        n9064) );
  OA22X1 U30336 ( .IN1(n2110), .IN2(n18912), .IN3(n2024), .IN4(n18891), .Q(
        n9065) );
  NAND4X0 U30337 ( .IN1(n9059), .IN2(n9060), .IN3(n9061), .IN4(n9062), .QN(
        s0_addr_o[24]) );
  OA22X1 U30338 ( .IN1(n1765), .IN2(n18848), .IN3(n1661), .IN4(n18827), .Q(
        n9059) );
  OA22X1 U30339 ( .IN1(n1937), .IN2(n18881), .IN3(n1851), .IN4(n18860), .Q(
        n9060) );
  OA22X1 U30340 ( .IN1(n2109), .IN2(n18914), .IN3(n2023), .IN4(n18891), .Q(
        n9061) );
  NAND4X0 U30341 ( .IN1(n9055), .IN2(n9056), .IN3(n9057), .IN4(n9058), .QN(
        s0_addr_o[25]) );
  OA22X1 U30342 ( .IN1(n1764), .IN2(n18848), .IN3(n1660), .IN4(n18827), .Q(
        n9055) );
  OA22X1 U30343 ( .IN1(n1936), .IN2(n18881), .IN3(n1850), .IN4(n18860), .Q(
        n9056) );
  OA22X1 U30344 ( .IN1(n2108), .IN2(n18914), .IN3(n2022), .IN4(n18891), .Q(
        n9057) );
  NAND4X0 U30345 ( .IN1(n9051), .IN2(n9052), .IN3(n9053), .IN4(n9054), .QN(
        s0_addr_o[26]) );
  OA22X1 U30346 ( .IN1(n1763), .IN2(n18848), .IN3(n1659), .IN4(n18828), .Q(
        n9051) );
  OA22X1 U30347 ( .IN1(n1935), .IN2(n18881), .IN3(n1849), .IN4(n18861), .Q(
        n9052) );
  OA22X1 U30348 ( .IN1(n2107), .IN2(n18914), .IN3(n2021), .IN4(n18892), .Q(
        n9053) );
  NAND4X0 U30349 ( .IN1(n9047), .IN2(n9048), .IN3(n9049), .IN4(n9050), .QN(
        s0_addr_o[27]) );
  OA22X1 U30350 ( .IN1(n1762), .IN2(n18848), .IN3(n1658), .IN4(n18828), .Q(
        n9047) );
  OA22X1 U30351 ( .IN1(n1934), .IN2(n18881), .IN3(n1848), .IN4(n18861), .Q(
        n9048) );
  OA22X1 U30352 ( .IN1(n2106), .IN2(n18914), .IN3(n2020), .IN4(n18892), .Q(
        n9049) );
  NAND4X0 U30353 ( .IN1(n9043), .IN2(n9044), .IN3(n9045), .IN4(n9046), .QN(
        s0_addr_o[28]) );
  OA22X1 U30354 ( .IN1(n1761), .IN2(n18848), .IN3(n1657), .IN4(n18828), .Q(
        n9043) );
  OA22X1 U30355 ( .IN1(n1933), .IN2(n18882), .IN3(n1847), .IN4(n18861), .Q(
        n9044) );
  OA22X1 U30356 ( .IN1(n2105), .IN2(n18915), .IN3(n2019), .IN4(n18892), .Q(
        n9045) );
  NAND4X0 U30357 ( .IN1(n9039), .IN2(n9040), .IN3(n9041), .IN4(n9042), .QN(
        s0_addr_o[29]) );
  OA22X1 U30358 ( .IN1(n1760), .IN2(n18849), .IN3(n1656), .IN4(n18829), .Q(
        n9039) );
  OA22X1 U30359 ( .IN1(n1932), .IN2(n18882), .IN3(n1846), .IN4(n18862), .Q(
        n9040) );
  OA22X1 U30360 ( .IN1(n2104), .IN2(n18915), .IN3(n2018), .IN4(n18893), .Q(
        n9041) );
  NAND4X0 U30361 ( .IN1(n9031), .IN2(n9032), .IN3(n9033), .IN4(n9034), .QN(
        s0_addr_o[30]) );
  OA22X1 U30362 ( .IN1(n1759), .IN2(n18848), .IN3(n1655), .IN4(n18829), .Q(
        n9031) );
  OA22X1 U30363 ( .IN1(n1931), .IN2(n18882), .IN3(n1845), .IN4(n18862), .Q(
        n9032) );
  OA22X1 U30364 ( .IN1(n2103), .IN2(n18915), .IN3(n2017), .IN4(n18893), .Q(
        n9033) );
  NAND4X0 U30365 ( .IN1(n9027), .IN2(n9028), .IN3(n9029), .IN4(n9030), .QN(
        s0_addr_o[31]) );
  OA22X1 U30366 ( .IN1(n1758), .IN2(n18852), .IN3(n1650), .IN4(n18830), .Q(
        n9027) );
  OA22X1 U30367 ( .IN1(n1930), .IN2(n18882), .IN3(n1844), .IN4(n18863), .Q(
        n9028) );
  OA22X1 U30368 ( .IN1(n2102), .IN2(n18915), .IN3(n2016), .IN4(n18894), .Q(
        n9029) );
  NAND4X0 U30369 ( .IN1(n8995), .IN2(n8996), .IN3(n8997), .IN4(n8998), .QN(
        s0_data_o[0]) );
  OA22X1 U30370 ( .IN1(n1741), .IN2(n18850), .IN3(n1636), .IN4(n18832), .Q(
        n8995) );
  OA22X1 U30371 ( .IN1(n1913), .IN2(n18880), .IN3(n1827), .IN4(n18865), .Q(
        n8996) );
  OA22X1 U30372 ( .IN1(n2085), .IN2(n18917), .IN3(n1999), .IN4(n18896), .Q(
        n8997) );
  NAND4X0 U30373 ( .IN1(n8951), .IN2(n8952), .IN3(n8953), .IN4(n8954), .QN(
        s0_data_o[1]) );
  OA22X1 U30374 ( .IN1(n1740), .IN2(n18851), .IN3(n1635), .IN4(n18834), .Q(
        n8951) );
  OA22X1 U30375 ( .IN1(n1912), .IN2(n18884), .IN3(n1826), .IN4(n18869), .Q(
        n8952) );
  OA22X1 U30376 ( .IN1(n2084), .IN2(n18913), .IN3(n1998), .IN4(n18897), .Q(
        n8953) );
  NAND4X0 U30377 ( .IN1(n8907), .IN2(n8908), .IN3(n8909), .IN4(n8910), .QN(
        s0_data_o[2]) );
  OA22X1 U30378 ( .IN1(n1739), .IN2(n18851), .IN3(n1634), .IN4(n18837), .Q(
        n8907) );
  OA22X1 U30379 ( .IN1(n1911), .IN2(n8839), .IN3(n1825), .IN4(n18872), .Q(
        n8908) );
  OA22X1 U30380 ( .IN1(n2083), .IN2(n18918), .IN3(n1997), .IN4(n18902), .Q(
        n8909) );
  NAND4X0 U30381 ( .IN1(n8895), .IN2(n8896), .IN3(n8897), .IN4(n8898), .QN(
        s0_data_o[3]) );
  OA22X1 U30382 ( .IN1(n1738), .IN2(n18846), .IN3(n1633), .IN4(n18837), .Q(
        n8895) );
  OA22X1 U30383 ( .IN1(n1910), .IN2(n8839), .IN3(n1824), .IN4(n18872), .Q(
        n8896) );
  OA22X1 U30384 ( .IN1(n2082), .IN2(n18918), .IN3(n1996), .IN4(n18903), .Q(
        n8897) );
  NAND4X0 U30385 ( .IN1(n8891), .IN2(n8892), .IN3(n8893), .IN4(n8894), .QN(
        s0_data_o[4]) );
  OA22X1 U30386 ( .IN1(n1737), .IN2(n18850), .IN3(n1632), .IN4(n18837), .Q(
        n8891) );
  OA22X1 U30387 ( .IN1(n1909), .IN2(n18881), .IN3(n1823), .IN4(n18872), .Q(
        n8892) );
  OA22X1 U30388 ( .IN1(n2081), .IN2(n18914), .IN3(n1995), .IN4(n18903), .Q(
        n8893) );
  NAND4X0 U30389 ( .IN1(n8887), .IN2(n8888), .IN3(n8889), .IN4(n8890), .QN(
        s0_data_o[5]) );
  OA22X1 U30390 ( .IN1(n1736), .IN2(n18851), .IN3(n1631), .IN4(n18837), .Q(
        n8887) );
  OA22X1 U30391 ( .IN1(n1908), .IN2(n8839), .IN3(n1822), .IN4(n18872), .Q(
        n8888) );
  OA22X1 U30392 ( .IN1(n2080), .IN2(n18916), .IN3(n1994), .IN4(n18903), .Q(
        n8889) );
  NAND4X0 U30393 ( .IN1(n8883), .IN2(n8884), .IN3(n8885), .IN4(n8886), .QN(
        s0_data_o[6]) );
  OA22X1 U30394 ( .IN1(n1735), .IN2(n18852), .IN3(n1630), .IN4(n18838), .Q(
        n8883) );
  OA22X1 U30395 ( .IN1(n1907), .IN2(n18884), .IN3(n1821), .IN4(n18870), .Q(
        n8884) );
  OA22X1 U30396 ( .IN1(n2079), .IN2(n18918), .IN3(n1993), .IN4(n18904), .Q(
        n8885) );
  NAND4X0 U30397 ( .IN1(n8879), .IN2(n8880), .IN3(n8881), .IN4(n8882), .QN(
        s0_data_o[7]) );
  OA22X1 U30398 ( .IN1(n1734), .IN2(n18852), .IN3(n1629), .IN4(n18838), .Q(
        n8879) );
  OA22X1 U30399 ( .IN1(n1906), .IN2(n18884), .IN3(n1820), .IN4(n18870), .Q(
        n8880) );
  OA22X1 U30400 ( .IN1(n2078), .IN2(n18918), .IN3(n1992), .IN4(n18904), .Q(
        n8881) );
  NAND4X0 U30401 ( .IN1(n8875), .IN2(n8876), .IN3(n8877), .IN4(n8878), .QN(
        s0_data_o[8]) );
  OA22X1 U30402 ( .IN1(n1733), .IN2(n18852), .IN3(n1628), .IN4(n18838), .Q(
        n8875) );
  OA22X1 U30403 ( .IN1(n1905), .IN2(n18884), .IN3(n1819), .IN4(n18870), .Q(
        n8876) );
  OA22X1 U30404 ( .IN1(n2077), .IN2(n18918), .IN3(n1991), .IN4(n18904), .Q(
        n8877) );
  NAND4X0 U30405 ( .IN1(n8871), .IN2(n8872), .IN3(n8873), .IN4(n8874), .QN(
        s0_data_o[9]) );
  OA22X1 U30406 ( .IN1(n1732), .IN2(n18852), .IN3(n1627), .IN4(n18837), .Q(
        n8871) );
  OA22X1 U30407 ( .IN1(n1904), .IN2(n18884), .IN3(n1818), .IN4(n18870), .Q(
        n8872) );
  OA22X1 U30408 ( .IN1(n2076), .IN2(n18918), .IN3(n1990), .IN4(n18905), .Q(
        n8873) );
  NAND4X0 U30409 ( .IN1(n8991), .IN2(n8992), .IN3(n8993), .IN4(n8994), .QN(
        s0_data_o[10]) );
  OA22X1 U30410 ( .IN1(n1731), .IN2(n18851), .IN3(n1626), .IN4(n18833), .Q(
        n8991) );
  OA22X1 U30411 ( .IN1(n1903), .IN2(n18878), .IN3(n1817), .IN4(n18866), .Q(
        n8992) );
  OA22X1 U30412 ( .IN1(n2075), .IN2(n18917), .IN3(n1989), .IN4(n18890), .Q(
        n8993) );
  NAND4X0 U30413 ( .IN1(n8987), .IN2(n8988), .IN3(n8989), .IN4(n8990), .QN(
        s0_data_o[11]) );
  OA22X1 U30414 ( .IN1(n1730), .IN2(n18852), .IN3(n1625), .IN4(n18833), .Q(
        n8987) );
  OA22X1 U30415 ( .IN1(n1902), .IN2(n18885), .IN3(n1816), .IN4(n18866), .Q(
        n8988) );
  OA22X1 U30416 ( .IN1(n2074), .IN2(n18917), .IN3(n1988), .IN4(n18896), .Q(
        n8989) );
  NAND4X0 U30417 ( .IN1(n8983), .IN2(n8984), .IN3(n8985), .IN4(n8986), .QN(
        s0_data_o[12]) );
  OA22X1 U30418 ( .IN1(n1729), .IN2(n18849), .IN3(n1624), .IN4(n18833), .Q(
        n8983) );
  OA22X1 U30419 ( .IN1(n1901), .IN2(n18881), .IN3(n1815), .IN4(n18866), .Q(
        n8984) );
  OA22X1 U30420 ( .IN1(n2073), .IN2(n18917), .IN3(n1987), .IN4(n18890), .Q(
        n8985) );
  NAND4X0 U30421 ( .IN1(n8979), .IN2(n8980), .IN3(n8981), .IN4(n8982), .QN(
        s0_data_o[13]) );
  OA22X1 U30422 ( .IN1(n1728), .IN2(n18850), .IN3(n1623), .IN4(n18834), .Q(
        n8979) );
  OA22X1 U30423 ( .IN1(n1900), .IN2(n18882), .IN3(n1814), .IN4(n18867), .Q(
        n8980) );
  OA22X1 U30424 ( .IN1(n2072), .IN2(n18915), .IN3(n1986), .IN4(n18897), .Q(
        n8981) );
  NAND4X0 U30425 ( .IN1(n8975), .IN2(n8976), .IN3(n8977), .IN4(n8978), .QN(
        s0_data_o[14]) );
  OA22X1 U30426 ( .IN1(n1727), .IN2(n18850), .IN3(n1622), .IN4(n18834), .Q(
        n8975) );
  OA22X1 U30427 ( .IN1(n1899), .IN2(n18881), .IN3(n1813), .IN4(n18867), .Q(
        n8976) );
  OA22X1 U30428 ( .IN1(n2071), .IN2(n18914), .IN3(n1985), .IN4(n18897), .Q(
        n8977) );
  NAND4X0 U30429 ( .IN1(n8971), .IN2(n8972), .IN3(n8973), .IN4(n8974), .QN(
        s0_data_o[15]) );
  OA22X1 U30430 ( .IN1(n1726), .IN2(n18850), .IN3(n1621), .IN4(n18834), .Q(
        n8971) );
  OA22X1 U30431 ( .IN1(n1898), .IN2(n18882), .IN3(n1812), .IN4(n18867), .Q(
        n8972) );
  OA22X1 U30432 ( .IN1(n2070), .IN2(n18915), .IN3(n1984), .IN4(n18897), .Q(
        n8973) );
  NAND4X0 U30433 ( .IN1(n8967), .IN2(n8968), .IN3(n8969), .IN4(n8970), .QN(
        s0_data_o[16]) );
  OA22X1 U30434 ( .IN1(n1725), .IN2(n18850), .IN3(n1620), .IN4(n18835), .Q(
        n8967) );
  OA22X1 U30435 ( .IN1(n1897), .IN2(n18878), .IN3(n1811), .IN4(n18868), .Q(
        n8968) );
  OA22X1 U30436 ( .IN1(n2069), .IN2(n18911), .IN3(n1983), .IN4(n18898), .Q(
        n8969) );
  NAND4X0 U30437 ( .IN1(n8963), .IN2(n8964), .IN3(n8965), .IN4(n8966), .QN(
        s0_data_o[17]) );
  OA22X1 U30438 ( .IN1(n1724), .IN2(n18851), .IN3(n1619), .IN4(n18835), .Q(
        n8963) );
  OA22X1 U30439 ( .IN1(n1896), .IN2(n18883), .IN3(n1810), .IN4(n18868), .Q(
        n8964) );
  OA22X1 U30440 ( .IN1(n2068), .IN2(n18917), .IN3(n1982), .IN4(n18898), .Q(
        n8965) );
  NAND4X0 U30441 ( .IN1(n8959), .IN2(n8960), .IN3(n8961), .IN4(n8962), .QN(
        s0_data_o[18]) );
  OA22X1 U30442 ( .IN1(n1723), .IN2(n18851), .IN3(n1618), .IN4(n18835), .Q(
        n8959) );
  OA22X1 U30443 ( .IN1(n1895), .IN2(n18880), .IN3(n1809), .IN4(n18868), .Q(
        n8960) );
  OA22X1 U30444 ( .IN1(n2067), .IN2(n18911), .IN3(n1981), .IN4(n18898), .Q(
        n8961) );
  NAND4X0 U30445 ( .IN1(n8955), .IN2(n8956), .IN3(n8957), .IN4(n8958), .QN(
        s0_data_o[19]) );
  OA22X1 U30446 ( .IN1(n1722), .IN2(n18851), .IN3(n1617), .IN4(n18835), .Q(
        n8955) );
  OA22X1 U30447 ( .IN1(n1894), .IN2(n18884), .IN3(n1808), .IN4(n18869), .Q(
        n8956) );
  OA22X1 U30448 ( .IN1(n2066), .IN2(n18914), .IN3(n1980), .IN4(n18898), .Q(
        n8957) );
  NAND4X0 U30449 ( .IN1(n8947), .IN2(n8948), .IN3(n8949), .IN4(n8950), .QN(
        s0_data_o[20]) );
  OA22X1 U30450 ( .IN1(n1721), .IN2(n18847), .IN3(n1616), .IN4(n18834), .Q(
        n8947) );
  OA22X1 U30451 ( .IN1(n1893), .IN2(n18884), .IN3(n1807), .IN4(n18869), .Q(
        n8948) );
  OA22X1 U30452 ( .IN1(n2065), .IN2(n18918), .IN3(n1979), .IN4(n18897), .Q(
        n8949) );
  NAND4X0 U30453 ( .IN1(n8943), .IN2(n8944), .IN3(n8945), .IN4(n8946), .QN(
        s0_data_o[21]) );
  OA22X1 U30454 ( .IN1(n1720), .IN2(n18850), .IN3(n1615), .IN4(n18837), .Q(
        n8943) );
  OA22X1 U30455 ( .IN1(n1892), .IN2(n18883), .IN3(n1806), .IN4(n18870), .Q(
        n8944) );
  OA22X1 U30456 ( .IN1(n2064), .IN2(n18916), .IN3(n1978), .IN4(n18899), .Q(
        n8945) );
  NAND4X0 U30457 ( .IN1(n8939), .IN2(n8940), .IN3(n8941), .IN4(n8942), .QN(
        s0_data_o[22]) );
  OA22X1 U30458 ( .IN1(n1719), .IN2(n18850), .IN3(n1614), .IN4(n18821), .Q(
        n8939) );
  OA22X1 U30459 ( .IN1(n1891), .IN2(n18880), .IN3(n1805), .IN4(n18870), .Q(
        n8940) );
  OA22X1 U30460 ( .IN1(n2063), .IN2(n18913), .IN3(n1977), .IN4(n18899), .Q(
        n8941) );
  NAND4X0 U30461 ( .IN1(n8935), .IN2(n8936), .IN3(n8937), .IN4(n8938), .QN(
        s0_data_o[23]) );
  OA22X1 U30462 ( .IN1(n1718), .IN2(n18851), .IN3(n1613), .IN4(n18839), .Q(
        n8935) );
  OA22X1 U30463 ( .IN1(n1890), .IN2(n18879), .IN3(n1804), .IN4(n18870), .Q(
        n8936) );
  OA22X1 U30464 ( .IN1(n2062), .IN2(n18917), .IN3(n1976), .IN4(n18899), .Q(
        n8937) );
  NAND4X0 U30465 ( .IN1(n8931), .IN2(n8932), .IN3(n8933), .IN4(n8934), .QN(
        s0_data_o[24]) );
  OA22X1 U30466 ( .IN1(n1717), .IN2(n18852), .IN3(n1612), .IN4(n18836), .Q(
        n8931) );
  OA22X1 U30467 ( .IN1(n1889), .IN2(n18884), .IN3(n1803), .IN4(n18871), .Q(
        n8932) );
  OA22X1 U30468 ( .IN1(n2061), .IN2(n18918), .IN3(n1975), .IN4(n18900), .Q(
        n8933) );
  NAND4X0 U30469 ( .IN1(n8927), .IN2(n8928), .IN3(n8929), .IN4(n8930), .QN(
        s0_data_o[25]) );
  OA22X1 U30470 ( .IN1(n1716), .IN2(n18849), .IN3(n1611), .IN4(n18836), .Q(
        n8927) );
  OA22X1 U30471 ( .IN1(n1888), .IN2(n18883), .IN3(n1802), .IN4(n18871), .Q(
        n8928) );
  OA22X1 U30472 ( .IN1(n2060), .IN2(n18916), .IN3(n1974), .IN4(n18900), .Q(
        n8929) );
  NAND4X0 U30473 ( .IN1(n8923), .IN2(n8924), .IN3(n8925), .IN4(n8926), .QN(
        s0_data_o[26]) );
  OA22X1 U30474 ( .IN1(n1715), .IN2(n18847), .IN3(n1610), .IN4(n18836), .Q(
        n8923) );
  OA22X1 U30475 ( .IN1(n1887), .IN2(n18880), .IN3(n1801), .IN4(n18871), .Q(
        n8924) );
  OA22X1 U30476 ( .IN1(n2059), .IN2(n18913), .IN3(n1973), .IN4(n18900), .Q(
        n8925) );
  NAND4X0 U30477 ( .IN1(n8919), .IN2(n8920), .IN3(n8921), .IN4(n8922), .QN(
        s0_data_o[27]) );
  OA22X1 U30478 ( .IN1(n1714), .IN2(n18847), .IN3(n1609), .IN4(n18839), .Q(
        n8919) );
  OA22X1 U30479 ( .IN1(n1886), .IN2(n18883), .IN3(n1800), .IN4(n18870), .Q(
        n8920) );
  OA22X1 U30480 ( .IN1(n2058), .IN2(n18917), .IN3(n1972), .IN4(n18901), .Q(
        n8921) );
  NAND4X0 U30481 ( .IN1(n8915), .IN2(n8916), .IN3(n8917), .IN4(n8918), .QN(
        s0_data_o[28]) );
  OA22X1 U30482 ( .IN1(n1713), .IN2(n18845), .IN3(n1608), .IN4(n18836), .Q(
        n8915) );
  OA22X1 U30483 ( .IN1(n1885), .IN2(n8839), .IN3(n1799), .IN4(n18871), .Q(
        n8916) );
  OA22X1 U30484 ( .IN1(n2057), .IN2(n18916), .IN3(n1971), .IN4(n18901), .Q(
        n8917) );
  NAND4X0 U30485 ( .IN1(n8911), .IN2(n8912), .IN3(n8913), .IN4(n8914), .QN(
        s0_data_o[29]) );
  OA22X1 U30486 ( .IN1(n1712), .IN2(n8841), .IN3(n1607), .IN4(n18838), .Q(
        n8911) );
  OA22X1 U30487 ( .IN1(n1884), .IN2(n8839), .IN3(n1798), .IN4(n18870), .Q(
        n8912) );
  OA22X1 U30488 ( .IN1(n2056), .IN2(n18913), .IN3(n1970), .IN4(n18901), .Q(
        n8913) );
  NAND4X0 U30489 ( .IN1(n8903), .IN2(n8904), .IN3(n8905), .IN4(n8906), .QN(
        s0_data_o[30]) );
  OA22X1 U30490 ( .IN1(n1711), .IN2(n8841), .IN3(n1606), .IN4(n18837), .Q(
        n8903) );
  OA22X1 U30491 ( .IN1(n1883), .IN2(n8839), .IN3(n1797), .IN4(n18872), .Q(
        n8904) );
  OA22X1 U30492 ( .IN1(n2055), .IN2(n18917), .IN3(n1969), .IN4(n18902), .Q(
        n8905) );
  NAND4X0 U30493 ( .IN1(n8899), .IN2(n8900), .IN3(n8901), .IN4(n8902), .QN(
        s0_data_o[31]) );
  OA22X1 U30494 ( .IN1(n1710), .IN2(n18847), .IN3(n1605), .IN4(n18837), .Q(
        n8899) );
  OA22X1 U30495 ( .IN1(n1882), .IN2(n18885), .IN3(n1796), .IN4(n18872), .Q(
        n8900) );
  OA22X1 U30496 ( .IN1(n2054), .IN2(n18912), .IN3(n1968), .IN4(n18902), .Q(
        n8901) );
  NAND3X0 U30497 ( .IN1(n14825), .IN2(n14824), .IN3(n3845), .QN(n5101) );
  NAND3X0 U30498 ( .IN1(n14823), .IN2(n14824), .IN3(n14825), .QN(n5099) );
  NAND3X0 U30499 ( .IN1(n14825), .IN2(n14823), .IN3(n3851), .QN(n5103) );
  NAND3X0 U30500 ( .IN1(n14820), .IN2(n14819), .IN3(n3800), .QN(n5397) );
  NAND3X0 U30501 ( .IN1(n14818), .IN2(n14819), .IN3(n14820), .QN(n5395) );
  NAND3X0 U30502 ( .IN1(n14820), .IN2(n14818), .IN3(n3806), .QN(n5399) );
  NAND3X0 U30503 ( .IN1(n14858), .IN2(n14857), .IN3(n4160), .QN(n7357) );
  NAND3X0 U30504 ( .IN1(n14856), .IN2(n14857), .IN3(n14858), .QN(n7355) );
  NAND3X0 U30505 ( .IN1(n14858), .IN2(n14856), .IN3(n4166), .QN(n7359) );
  NAND3X0 U30506 ( .IN1(n14843), .IN2(n14842), .IN3(n3755), .QN(n5693) );
  NAND3X0 U30507 ( .IN1(n14841), .IN2(n14842), .IN3(n14843), .QN(n5691) );
  NAND3X0 U30508 ( .IN1(n14843), .IN2(n14841), .IN3(n3761), .QN(n5695) );
  NAND3X0 U30509 ( .IN1(n14839), .IN2(n14838), .IN3(n3710), .QN(n5989) );
  NAND3X0 U30510 ( .IN1(n14837), .IN2(n14838), .IN3(n14839), .QN(n5987) );
  NAND3X0 U30511 ( .IN1(n14839), .IN2(n14837), .IN3(n3716), .QN(n5991) );
  NAND3X0 U30512 ( .IN1(n14855), .IN2(n14854), .IN3(n4115), .QN(n7653) );
  NAND3X0 U30513 ( .IN1(n14853), .IN2(n14854), .IN3(n14855), .QN(n7651) );
  NAND3X0 U30514 ( .IN1(n14855), .IN2(n14853), .IN3(n4121), .QN(n7655) );
  NAND3X0 U30515 ( .IN1(n14868), .IN2(n14867), .IN3(n4070), .QN(n7949) );
  NAND3X0 U30516 ( .IN1(n14866), .IN2(n14867), .IN3(n14868), .QN(n7947) );
  NAND3X0 U30517 ( .IN1(n14868), .IN2(n14866), .IN3(n4076), .QN(n7951) );
  NAND3X0 U30518 ( .IN1(n14846), .IN2(n14845), .IN3(n3665), .QN(n6285) );
  NAND3X0 U30519 ( .IN1(n14844), .IN2(n14845), .IN3(n14846), .QN(n6283) );
  NAND3X0 U30520 ( .IN1(n14846), .IN2(n14844), .IN3(n3671), .QN(n6287) );
  NAND3X0 U30521 ( .IN1(n14850), .IN2(n14849), .IN3(n3620), .QN(n6581) );
  NAND3X0 U30522 ( .IN1(n14848), .IN2(n14849), .IN3(n14850), .QN(n6579) );
  NAND3X0 U30523 ( .IN1(n14850), .IN2(n14848), .IN3(n3626), .QN(n6583) );
  NAND3X0 U30524 ( .IN1(n14865), .IN2(n14864), .IN3(n4025), .QN(n8245) );
  NAND3X0 U30525 ( .IN1(n14863), .IN2(n14864), .IN3(n14865), .QN(n8243) );
  NAND3X0 U30526 ( .IN1(n14865), .IN2(n14863), .IN3(n4031), .QN(n8247) );
  NAND3X0 U30527 ( .IN1(n14871), .IN2(n14870), .IN3(n3980), .QN(n8541) );
  NAND3X0 U30528 ( .IN1(n14869), .IN2(n14870), .IN3(n14871), .QN(n8539) );
  NAND3X0 U30529 ( .IN1(n14871), .IN2(n14869), .IN3(n3986), .QN(n8543) );
  NAND3X0 U30530 ( .IN1(n14861), .IN2(n14860), .IN3(n3575), .QN(n6877) );
  NAND3X0 U30531 ( .IN1(n14859), .IN2(n14860), .IN3(n14861), .QN(n6875) );
  NAND3X0 U30532 ( .IN1(n14861), .IN2(n14859), .IN3(n3581), .QN(n6879) );
  NAND3X0 U30533 ( .IN1(n14874), .IN2(n14873), .IN3(n3530), .QN(n8837) );
  NAND3X0 U30534 ( .IN1(n14872), .IN2(n14873), .IN3(n14874), .QN(n8835) );
  NAND3X0 U30535 ( .IN1(n14874), .IN2(n14872), .IN3(n3536), .QN(n8839) );
  NAND3X0 U30536 ( .IN1(n14829), .IN2(n14828), .IN3(n3935), .QN(n4509) );
  NAND3X0 U30537 ( .IN1(n14827), .IN2(n14828), .IN3(n3940), .QN(n4508) );
  NAND3X0 U30538 ( .IN1(n14827), .IN2(n14828), .IN3(n14829), .QN(n4507) );
  NAND3X0 U30539 ( .IN1(n14829), .IN2(n14827), .IN3(n3941), .QN(n4511) );
  NAND3X0 U30540 ( .IN1(n14834), .IN2(n14833), .IN3(n3890), .QN(n4805) );
  NAND3X0 U30541 ( .IN1(n14832), .IN2(n14833), .IN3(n14834), .QN(n4803) );
  NAND3X0 U30542 ( .IN1(n14834), .IN2(n14832), .IN3(n3896), .QN(n4807) );
  NAND3X0 U30543 ( .IN1(n3845), .IN2(n14825), .IN3(n3851), .QN(n5105) );
  NAND3X0 U30544 ( .IN1(n3800), .IN2(n14820), .IN3(n3806), .QN(n5401) );
  NAND3X0 U30545 ( .IN1(n4160), .IN2(n14858), .IN3(n4166), .QN(n7361) );
  NAND3X0 U30546 ( .IN1(n3755), .IN2(n14843), .IN3(n3761), .QN(n5697) );
  NAND3X0 U30547 ( .IN1(n3710), .IN2(n14839), .IN3(n3716), .QN(n5993) );
  NAND3X0 U30548 ( .IN1(n4115), .IN2(n14855), .IN3(n4121), .QN(n7657) );
  NAND3X0 U30549 ( .IN1(n4070), .IN2(n14868), .IN3(n4076), .QN(n7953) );
  NAND3X0 U30550 ( .IN1(n3665), .IN2(n14846), .IN3(n3671), .QN(n6289) );
  NAND3X0 U30551 ( .IN1(n3620), .IN2(n14850), .IN3(n3626), .QN(n6585) );
  NAND3X0 U30552 ( .IN1(n4025), .IN2(n14865), .IN3(n4031), .QN(n8249) );
  NAND3X0 U30553 ( .IN1(n3980), .IN2(n14871), .IN3(n3986), .QN(n8545) );
  NAND3X0 U30554 ( .IN1(n3575), .IN2(n14861), .IN3(n3581), .QN(n6881) );
  NAND3X0 U30555 ( .IN1(n3530), .IN2(n14874), .IN3(n3536), .QN(n8841) );
  NAND3X0 U30556 ( .IN1(n3940), .IN2(n14828), .IN3(n3935), .QN(n4510) );
  NAND3X0 U30557 ( .IN1(n3940), .IN2(n14827), .IN3(n3941), .QN(n4512) );
  NAND3X0 U30558 ( .IN1(n3935), .IN2(n14829), .IN3(n3941), .QN(n4513) );
  NAND3X0 U30559 ( .IN1(n3890), .IN2(n14834), .IN3(n3896), .QN(n4809) );
  INVX0 U30560 ( .IN(n21089), .QN(n21086) );
  INVX0 U30561 ( .IN(n21088), .QN(n21087) );
  INVX0 U30562 ( .IN(n21089), .QN(n21085) );
  NAND2X0 U30563 ( .IN1(n14847), .IN2(n14835), .QN(n14523) );
  NAND2X0 U30564 ( .IN1(n14821), .IN2(n14830), .QN(n14533) );
  NAND2X0 U30565 ( .IN1(n15176), .IN2(n15174), .QN(n14900) );
  NAND2X0 U30566 ( .IN1(n15177), .IN2(n15174), .QN(n14905) );
  NAND2X0 U30567 ( .IN1(n15169), .IN2(n15172), .QN(n14915) );
  NAND2X0 U30568 ( .IN1(n15482), .IN2(n15479), .QN(n15210) );
  NAND2X0 U30569 ( .IN1(n15474), .IN2(n15477), .QN(n15220) );
  NAND2X0 U30570 ( .IN1(n15786), .IN2(n15784), .QN(n15510) );
  NAND2X0 U30571 ( .IN1(n15787), .IN2(n15784), .QN(n15515) );
  NAND2X0 U30572 ( .IN1(n15779), .IN2(n15782), .QN(n15525) );
  NAND2X0 U30573 ( .IN1(n16092), .IN2(n16089), .QN(n15820) );
  NAND2X0 U30574 ( .IN1(n16084), .IN2(n16087), .QN(n15830) );
  NAND2X0 U30575 ( .IN1(n16396), .IN2(n16394), .QN(n16120) );
  NAND2X0 U30576 ( .IN1(n16397), .IN2(n16394), .QN(n16125) );
  NAND2X0 U30577 ( .IN1(n16389), .IN2(n16392), .QN(n16135) );
  NAND2X0 U30578 ( .IN1(n16702), .IN2(n16699), .QN(n16430) );
  NAND2X0 U30579 ( .IN1(n16694), .IN2(n16697), .QN(n16440) );
  NAND2X0 U30580 ( .IN1(n17041), .IN2(n17032), .QN(n16730) );
  NAND2X0 U30581 ( .IN1(n17056), .IN2(n17032), .QN(n16735) );
  NAND2X0 U30582 ( .IN1(n17006), .IN2(n17023), .QN(n16745) );
  NAND2X0 U30583 ( .IN1(n15177), .IN2(n15171), .QN(n14912) );
  NAND2X0 U30584 ( .IN1(n15787), .IN2(n15781), .QN(n15522) );
  NAND2X0 U30585 ( .IN1(n16397), .IN2(n16391), .QN(n16132) );
  NAND2X0 U30586 ( .IN1(n17056), .IN2(n17015), .QN(n16742) );
  NAND2X0 U30587 ( .IN1(n15169), .IN2(n15170), .QN(n14910) );
  NAND2X0 U30588 ( .IN1(n15779), .IN2(n15780), .QN(n15520) );
  NAND2X0 U30589 ( .IN1(n16389), .IN2(n16390), .QN(n16130) );
  NAND2X0 U30590 ( .IN1(n17006), .IN2(n17007), .QN(n16740) );
  NOR2X0 U30591 ( .IN1(n13627), .IN2(n21001), .QN(n13632) );
  NOR2X0 U30592 ( .IN1(n13318), .IN2(n21000), .QN(n13323) );
  NOR2X0 U30593 ( .IN1(n11152), .IN2(n20990), .QN(n11157) );
  NOR2X0 U30594 ( .IN1(n13009), .IN2(n20996), .QN(n13014) );
  NOR2X0 U30595 ( .IN1(n12700), .IN2(n20998), .QN(n12705) );
  NOR2X0 U30596 ( .IN1(n10843), .IN2(n20992), .QN(n10848) );
  NOR2X0 U30597 ( .IN1(n10533), .IN2(n20991), .QN(n10538) );
  NOR2X0 U30598 ( .IN1(n12391), .IN2(n20997), .QN(n12396) );
  NOR2X0 U30599 ( .IN1(n12082), .IN2(n20993), .QN(n12087) );
  NOR2X0 U30600 ( .IN1(n10224), .IN2(n20987), .QN(n10229) );
  NOR2X0 U30601 ( .IN1(n9914), .IN2(n20989), .QN(n9919) );
  NOR2X0 U30602 ( .IN1(n11772), .IN2(n20995), .QN(n11777) );
  NOR2X0 U30603 ( .IN1(n11462), .IN2(n20994), .QN(n11467) );
  NOR2X0 U30604 ( .IN1(n9604), .IN2(n20988), .QN(n9609) );
  NOR2X0 U30605 ( .IN1(n9293), .IN2(n20986), .QN(n9298) );
  NOR2X0 U30606 ( .IN1(n14270), .IN2(n20999), .QN(n14275) );
  NAND4X0 U30607 ( .IN1(n14265), .IN2(n14266), .IN3(n14267), .IN4(n14268), 
        .QN(n21105) );
  OA22X1 U30608 ( .IN1(n1741), .IN2(n19641), .IN3(n1636), .IN4(n19622), .Q(
        n14265) );
  OA22X1 U30609 ( .IN1(n1913), .IN2(n19673), .IN3(n1827), .IN4(n19655), .Q(
        n14266) );
  OA22X1 U30610 ( .IN1(n2085), .IN2(n19706), .IN3(n1999), .IN4(n19688), .Q(
        n14267) );
  NAND4X0 U30611 ( .IN1(n14261), .IN2(n14262), .IN3(n14263), .IN4(n14264), 
        .QN(n21104) );
  OA22X1 U30612 ( .IN1(n1740), .IN2(n19640), .IN3(n1635), .IN4(n19631), .Q(
        n14261) );
  OA22X1 U30613 ( .IN1(n1912), .IN2(n19673), .IN3(n1826), .IN4(n19655), .Q(
        n14262) );
  OA22X1 U30614 ( .IN1(n2084), .IN2(n19706), .IN3(n1998), .IN4(n19688), .Q(
        n14263) );
  NAND4X0 U30615 ( .IN1(n14257), .IN2(n14258), .IN3(n14259), .IN4(n14260), 
        .QN(n21103) );
  OA22X1 U30616 ( .IN1(n1739), .IN2(n19643), .IN3(n1634), .IN4(n19623), .Q(
        n14257) );
  OA22X1 U30617 ( .IN1(n1911), .IN2(n19675), .IN3(n1825), .IN4(n19655), .Q(
        n14258) );
  OA22X1 U30618 ( .IN1(n2083), .IN2(n19708), .IN3(n1997), .IN4(n19688), .Q(
        n14259) );
  NAND4X0 U30619 ( .IN1(n14253), .IN2(n14254), .IN3(n14255), .IN4(n14256), 
        .QN(n21102) );
  OA22X1 U30620 ( .IN1(n1738), .IN2(n19639), .IN3(n1633), .IN4(n19631), .Q(
        n14253) );
  OA22X1 U30621 ( .IN1(n1910), .IN2(n19672), .IN3(n1824), .IN4(n19657), .Q(
        n14254) );
  OA22X1 U30622 ( .IN1(n2082), .IN2(n19705), .IN3(n1996), .IN4(n19690), .Q(
        n14255) );
  NAND4X0 U30623 ( .IN1(n14249), .IN2(n14250), .IN3(n14251), .IN4(n14252), 
        .QN(n21101) );
  OA22X1 U30624 ( .IN1(n1737), .IN2(n19639), .IN3(n1632), .IN4(n19625), .Q(
        n14249) );
  OA22X1 U30625 ( .IN1(n1909), .IN2(n19672), .IN3(n1823), .IN4(n19663), .Q(
        n14250) );
  OA22X1 U30626 ( .IN1(n2081), .IN2(n19705), .IN3(n1995), .IN4(n19696), .Q(
        n14251) );
  NAND4X0 U30627 ( .IN1(n14245), .IN2(n14246), .IN3(n14247), .IN4(n14248), 
        .QN(n21100) );
  OA22X1 U30628 ( .IN1(n1736), .IN2(n19639), .IN3(n1631), .IN4(n19623), .Q(
        n14245) );
  OA22X1 U30629 ( .IN1(n1908), .IN2(n19672), .IN3(n1822), .IN4(n19659), .Q(
        n14246) );
  OA22X1 U30630 ( .IN1(n2080), .IN2(n19705), .IN3(n1994), .IN4(n19692), .Q(
        n14247) );
  NAND4X0 U30631 ( .IN1(n14241), .IN2(n14242), .IN3(n14243), .IN4(n14244), 
        .QN(n21099) );
  OA22X1 U30632 ( .IN1(n1735), .IN2(n19639), .IN3(n1630), .IN4(n19622), .Q(
        n14241) );
  OA22X1 U30633 ( .IN1(n1907), .IN2(n19672), .IN3(n1821), .IN4(n19656), .Q(
        n14242) );
  OA22X1 U30634 ( .IN1(n2079), .IN2(n19705), .IN3(n1993), .IN4(n19689), .Q(
        n14243) );
  NAND4X0 U30635 ( .IN1(n14237), .IN2(n14238), .IN3(n14239), .IN4(n14240), 
        .QN(n21098) );
  OA22X1 U30636 ( .IN1(n1734), .IN2(n19640), .IN3(n1629), .IN4(n19622), .Q(
        n14237) );
  OA22X1 U30637 ( .IN1(n1906), .IN2(n19673), .IN3(n1820), .IN4(n19656), .Q(
        n14238) );
  OA22X1 U30638 ( .IN1(n2078), .IN2(n19706), .IN3(n1992), .IN4(n19689), .Q(
        n14239) );
  NAND4X0 U30639 ( .IN1(n14233), .IN2(n14234), .IN3(n14235), .IN4(n14236), 
        .QN(n21097) );
  OA22X1 U30640 ( .IN1(n1733), .IN2(n19642), .IN3(n1628), .IN4(n19622), .Q(
        n14233) );
  OA22X1 U30641 ( .IN1(n1905), .IN2(n19673), .IN3(n1819), .IN4(n19656), .Q(
        n14234) );
  OA22X1 U30642 ( .IN1(n2077), .IN2(n19706), .IN3(n1991), .IN4(n19689), .Q(
        n14235) );
  NAND4X0 U30643 ( .IN1(n14229), .IN2(n14230), .IN3(n14231), .IN4(n14232), 
        .QN(n21096) );
  OA22X1 U30644 ( .IN1(n1732), .IN2(n19641), .IN3(n1627), .IN4(n19625), .Q(
        n14229) );
  OA22X1 U30645 ( .IN1(n1904), .IN2(n19673), .IN3(n1818), .IN4(n19655), .Q(
        n14230) );
  OA22X1 U30646 ( .IN1(n2076), .IN2(n19706), .IN3(n1990), .IN4(n19688), .Q(
        n14231) );
  NAND4X0 U30647 ( .IN1(n14225), .IN2(n14226), .IN3(n14227), .IN4(n14228), 
        .QN(n21095) );
  OA22X1 U30648 ( .IN1(n1731), .IN2(n19643), .IN3(n1626), .IN4(n19624), .Q(
        n14225) );
  OA22X1 U30649 ( .IN1(n1903), .IN2(n19673), .IN3(n1817), .IN4(n19655), .Q(
        n14226) );
  OA22X1 U30650 ( .IN1(n2075), .IN2(n19706), .IN3(n1989), .IN4(n19688), .Q(
        n14227) );
  NAND4X0 U30651 ( .IN1(n14221), .IN2(n14222), .IN3(n14223), .IN4(n14224), 
        .QN(n21094) );
  OA22X1 U30652 ( .IN1(n1730), .IN2(n19640), .IN3(n1625), .IN4(n19627), .Q(
        n14221) );
  OA22X1 U30653 ( .IN1(n1902), .IN2(n19673), .IN3(n1816), .IN4(n19656), .Q(
        n14222) );
  OA22X1 U30654 ( .IN1(n2074), .IN2(n19706), .IN3(n1988), .IN4(n19689), .Q(
        n14223) );
  NAND4X0 U30655 ( .IN1(n14217), .IN2(n14218), .IN3(n14219), .IN4(n14220), 
        .QN(n21093) );
  OA22X1 U30656 ( .IN1(n1729), .IN2(n19642), .IN3(n1624), .IN4(n19623), .Q(
        n14217) );
  OA22X1 U30657 ( .IN1(n1901), .IN2(n19673), .IN3(n1815), .IN4(n19657), .Q(
        n14218) );
  OA22X1 U30658 ( .IN1(n2073), .IN2(n19706), .IN3(n1987), .IN4(n19690), .Q(
        n14219) );
  NAND4X0 U30659 ( .IN1(n14213), .IN2(n14214), .IN3(n14215), .IN4(n14216), 
        .QN(n21092) );
  OA22X1 U30660 ( .IN1(n1728), .IN2(n19641), .IN3(n1623), .IN4(n19623), .Q(
        n14213) );
  OA22X1 U30661 ( .IN1(n1900), .IN2(n19672), .IN3(n1814), .IN4(n19657), .Q(
        n14214) );
  OA22X1 U30662 ( .IN1(n2072), .IN2(n19705), .IN3(n1986), .IN4(n19690), .Q(
        n14215) );
  NAND4X0 U30663 ( .IN1(n14209), .IN2(n14210), .IN3(n14211), .IN4(n14212), 
        .QN(n21091) );
  OA22X1 U30664 ( .IN1(n1727), .IN2(n19643), .IN3(n1622), .IN4(n19623), .Q(
        n14209) );
  OA22X1 U30665 ( .IN1(n1899), .IN2(n19673), .IN3(n1813), .IN4(n19657), .Q(
        n14210) );
  OA22X1 U30666 ( .IN1(n2071), .IN2(n19706), .IN3(n1985), .IN4(n19690), .Q(
        n14211) );
  NAND4X0 U30667 ( .IN1(n14304), .IN2(n14305), .IN3(n14306), .IN4(n14307), 
        .QN(n21090) );
  OA22X1 U30668 ( .IN1(n1726), .IN2(n19642), .IN3(n1621), .IN4(n19621), .Q(
        n14304) );
  OA22X1 U30669 ( .IN1(n1898), .IN2(n19674), .IN3(n1812), .IN4(n19654), .Q(
        n14305) );
  OA22X1 U30670 ( .IN1(n2070), .IN2(n19707), .IN3(n1984), .IN4(n19687), .Q(
        n14306) );
  NAND3X0 U30671 ( .IN1(n3805), .IN2(n14819), .IN3(n3800), .QN(n5398) );
  NAND3X0 U30672 ( .IN1(n4165), .IN2(n14857), .IN3(n4160), .QN(n7358) );
  NAND3X0 U30673 ( .IN1(n3670), .IN2(n14845), .IN3(n3665), .QN(n6286) );
  NAND3X0 U30674 ( .IN1(n3625), .IN2(n14849), .IN3(n3620), .QN(n6582) );
  OA22X1 U30675 ( .IN1(n2257), .IN2(n19739), .IN3(n2171), .IN4(n19721), .Q(
        n14268) );
  OA22X1 U30676 ( .IN1(n2256), .IN2(n19740), .IN3(n2170), .IN4(n19721), .Q(
        n14264) );
  OA22X1 U30677 ( .IN1(n2255), .IN2(n19739), .IN3(n2169), .IN4(n19721), .Q(
        n14260) );
  OA22X1 U30678 ( .IN1(n2254), .IN2(n19738), .IN3(n2168), .IN4(n19723), .Q(
        n14256) );
  OA22X1 U30679 ( .IN1(n2253), .IN2(n19738), .IN3(n2167), .IN4(n19725), .Q(
        n14252) );
  OA22X1 U30680 ( .IN1(n2252), .IN2(n19738), .IN3(n2166), .IN4(n19726), .Q(
        n14248) );
  OA22X1 U30681 ( .IN1(n2251), .IN2(n19738), .IN3(n2165), .IN4(n19722), .Q(
        n14244) );
  OA22X1 U30682 ( .IN1(n2250), .IN2(n19739), .IN3(n2164), .IN4(n19722), .Q(
        n14240) );
  OA22X1 U30683 ( .IN1(n2249), .IN2(n19739), .IN3(n2163), .IN4(n19722), .Q(
        n14236) );
  OA22X1 U30684 ( .IN1(n2248), .IN2(n19739), .IN3(n2162), .IN4(n19721), .Q(
        n14232) );
  OA22X1 U30685 ( .IN1(n2247), .IN2(n19739), .IN3(n2161), .IN4(n19721), .Q(
        n14228) );
  OA22X1 U30686 ( .IN1(n2246), .IN2(n19740), .IN3(n2160), .IN4(n19722), .Q(
        n14224) );
  OA22X1 U30687 ( .IN1(n2245), .IN2(n19740), .IN3(n2159), .IN4(n19723), .Q(
        n14220) );
  OA22X1 U30688 ( .IN1(n2244), .IN2(n19740), .IN3(n2158), .IN4(n19723), .Q(
        n14216) );
  OA22X1 U30689 ( .IN1(n2243), .IN2(n19740), .IN3(n2157), .IN4(n19723), .Q(
        n14212) );
  OA22X1 U30690 ( .IN1(n2242), .IN2(n19740), .IN3(n2156), .IN4(n19720), .Q(
        n14307) );
  OA22X1 U30691 ( .IN1(n2310), .IN2(n19741), .IN3(n2224), .IN4(n19724), .Q(
        n9131) );
  OA22X1 U30692 ( .IN1(n2309), .IN2(n19743), .IN3(n2223), .IN4(n19730), .Q(
        n7190) );
  OA22X1 U30693 ( .IN1(n2308), .IN2(n19743), .IN3(n2222), .IN4(n19730), .Q(
        n7186) );
  OA22X1 U30694 ( .IN1(n2307), .IN2(n19743), .IN3(n2221), .IN4(n19730), .Q(
        n7182) );
  OA22X1 U30695 ( .IN1(n2306), .IN2(n19738), .IN3(n2220), .IN4(n19730), .Q(
        n7170) );
  OA22X1 U30696 ( .IN1(n2305), .IN2(n19741), .IN3(n2219), .IN4(n19724), .Q(
        n7350) );
  OA22X1 U30697 ( .IN1(n2304), .IN2(n19742), .IN3(n2218), .IN4(n19722), .Q(
        n7306) );
  OA22X1 U30698 ( .IN1(n2299), .IN2(n19742), .IN3(n2213), .IN4(n19728), .Q(
        n7270) );
  OA22X1 U30699 ( .IN1(n2298), .IN2(n19740), .IN3(n2212), .IN4(n19728), .Q(
        n7266) );
  OA22X1 U30700 ( .IN1(n2297), .IN2(n19741), .IN3(n2211), .IN4(n19728), .Q(
        n7262) );
  OA22X1 U30701 ( .IN1(n2296), .IN2(n19738), .IN3(n2210), .IN4(n19729), .Q(
        n7258) );
  OA22X1 U30702 ( .IN1(n2295), .IN2(n19741), .IN3(n2209), .IN4(n19724), .Q(
        n7346) );
  OA22X1 U30703 ( .IN1(n2294), .IN2(n19741), .IN3(n2208), .IN4(n19725), .Q(
        n7342) );
  OA22X1 U30704 ( .IN1(n2293), .IN2(n19739), .IN3(n2207), .IN4(n19725), .Q(
        n7338) );
  OA22X1 U30705 ( .IN1(n2292), .IN2(n19740), .IN3(n2206), .IN4(n19725), .Q(
        n7334) );
  OA22X1 U30706 ( .IN1(n2291), .IN2(n19742), .IN3(n2205), .IN4(n19726), .Q(
        n7330) );
  OA22X1 U30707 ( .IN1(n2290), .IN2(n19741), .IN3(n2204), .IN4(n19726), .Q(
        n7326) );
  OA22X1 U30708 ( .IN1(n2289), .IN2(n19742), .IN3(n2203), .IN4(n19726), .Q(
        n7322) );
  OA22X1 U30709 ( .IN1(n2288), .IN2(n19742), .IN3(n2202), .IN4(n19727), .Q(
        n7318) );
  OA22X1 U30710 ( .IN1(n2287), .IN2(n19742), .IN3(n2201), .IN4(n19727), .Q(
        n7314) );
  OA22X1 U30711 ( .IN1(n2286), .IN2(n19742), .IN3(n2200), .IN4(n19727), .Q(
        n7310) );
  OA22X1 U30712 ( .IN1(n2285), .IN2(n19739), .IN3(n2199), .IN4(n19722), .Q(
        n7302) );
  OA22X1 U30713 ( .IN1(n2284), .IN2(n19738), .IN3(n2198), .IN4(n19722), .Q(
        n7298) );
  OA22X1 U30714 ( .IN1(n2283), .IN2(n19741), .IN3(n2197), .IN4(n19721), .Q(
        n7294) );
  OA22X1 U30715 ( .IN1(n2282), .IN2(n19741), .IN3(n2196), .IN4(n19721), .Q(
        n7290) );
  OA22X1 U30716 ( .IN1(n2241), .IN2(n19741), .IN3(n2155), .IN4(n19729), .Q(
        n7254) );
  OA22X1 U30717 ( .IN1(n2240), .IN2(n19739), .IN3(n2154), .IN4(n19729), .Q(
        n7250) );
  OA22X1 U30718 ( .IN1(n2239), .IN2(n19743), .IN3(n2153), .IN4(n19723), .Q(
        n7246) );
  OA22X1 U30719 ( .IN1(n2238), .IN2(n19740), .IN3(n2152), .IN4(n19728), .Q(
        n7242) );
  OA22X1 U30720 ( .IN1(n2237), .IN2(n19739), .IN3(n2151), .IN4(n19729), .Q(
        n7238) );
  OA22X1 U30721 ( .IN1(n2236), .IN2(n19740), .IN3(n2150), .IN4(n19725), .Q(
        n7234) );
  OA22X1 U30722 ( .IN1(n2235), .IN2(n19741), .IN3(n2149), .IN4(n19726), .Q(
        n7230) );
  OA22X1 U30723 ( .IN1(n2234), .IN2(n19738), .IN3(n2148), .IN4(n19727), .Q(
        n7226) );
  OA22X1 U30724 ( .IN1(n2233), .IN2(n19743), .IN3(n2147), .IN4(n19727), .Q(
        n7222) );
  OA22X1 U30725 ( .IN1(n2232), .IN2(n19738), .IN3(n2146), .IN4(n19728), .Q(
        n7218) );
  OA22X1 U30726 ( .IN1(n2231), .IN2(n19743), .IN3(n2145), .IN4(n19729), .Q(
        n7214) );
  OA22X1 U30727 ( .IN1(n2230), .IN2(n19743), .IN3(n2144), .IN4(n19722), .Q(
        n7210) );
  OA22X1 U30728 ( .IN1(n2229), .IN2(n19743), .IN3(n2143), .IN4(n19730), .Q(
        n7206) );
  OA22X1 U30729 ( .IN1(n2228), .IN2(n19743), .IN3(n2142), .IN4(n19722), .Q(
        n7202) );
  OA22X1 U30730 ( .IN1(n2227), .IN2(n19743), .IN3(n2141), .IN4(n19730), .Q(
        n7198) );
  OA22X1 U30731 ( .IN1(n2226), .IN2(n19738), .IN3(n2140), .IN4(n19722), .Q(
        n7194) );
  OA22X1 U30732 ( .IN1(n2310), .IN2(n19604), .IN3(n2224), .IN4(n19598), .Q(
        n7354) );
  OA22X1 U30733 ( .IN1(n2309), .IN2(n19611), .IN3(n2223), .IN4(n19597), .Q(
        n7390) );
  OA22X1 U30734 ( .IN1(n2308), .IN2(n19611), .IN3(n2222), .IN4(n19597), .Q(
        n7386) );
  OA22X1 U30735 ( .IN1(n2307), .IN2(n19611), .IN3(n2221), .IN4(n19598), .Q(
        n7382) );
  OA22X1 U30736 ( .IN1(n2306), .IN2(n19611), .IN3(n2220), .IN4(n19598), .Q(
        n7378) );
  OA22X1 U30737 ( .IN1(n2305), .IN2(n19604), .IN3(n2219), .IN4(n19581), .Q(
        n7646) );
  OA22X1 U30738 ( .IN1(n2304), .IN2(n19606), .IN3(n2218), .IN4(n19584), .Q(
        n7602) );
  OA22X1 U30739 ( .IN1(n2303), .IN2(n19609), .IN3(n2217), .IN4(n19588), .Q(
        n7558) );
  OA22X1 U30740 ( .IN1(n2302), .IN2(n19605), .IN3(n2216), .IN4(n19585), .Q(
        n7546) );
  OA22X1 U30741 ( .IN1(n2301), .IN2(n19609), .IN3(n2215), .IN4(n19589), .Q(
        n7542) );
  OA22X1 U30742 ( .IN1(n2300), .IN2(n19610), .IN3(n2214), .IN4(n19590), .Q(
        n7538) );
  OA22X1 U30743 ( .IN1(n2299), .IN2(n19608), .IN3(n2213), .IN4(n19591), .Q(
        n7534) );
  OA22X1 U30744 ( .IN1(n2298), .IN2(n19608), .IN3(n2212), .IN4(n19593), .Q(
        n7530) );
  OA22X1 U30745 ( .IN1(n2297), .IN2(n19608), .IN3(n2211), .IN4(n19589), .Q(
        n7526) );
  OA22X1 U30746 ( .IN1(n2296), .IN2(n19608), .IN3(n2210), .IN4(n19589), .Q(
        n7522) );
  OA22X1 U30747 ( .IN1(n2295), .IN2(n19604), .IN3(n2209), .IN4(n19581), .Q(
        n7642) );
  OA22X1 U30748 ( .IN1(n2294), .IN2(n19604), .IN3(n2208), .IN4(n19581), .Q(
        n7638) );
  OA22X1 U30749 ( .IN1(n2293), .IN2(n19604), .IN3(n2207), .IN4(n19582), .Q(
        n7634) );
  OA22X1 U30750 ( .IN1(n2292), .IN2(n19605), .IN3(n2206), .IN4(n19582), .Q(
        n7630) );
  OA22X1 U30751 ( .IN1(n2291), .IN2(n19605), .IN3(n2205), .IN4(n19582), .Q(
        n7626) );
  OA22X1 U30752 ( .IN1(n2290), .IN2(n19605), .IN3(n2204), .IN4(n19583), .Q(
        n7622) );
  OA22X1 U30753 ( .IN1(n2289), .IN2(n19605), .IN3(n2203), .IN4(n19583), .Q(
        n7618) );
  OA22X1 U30754 ( .IN1(n2288), .IN2(n19606), .IN3(n2202), .IN4(n19583), .Q(
        n7614) );
  OA22X1 U30755 ( .IN1(n2287), .IN2(n19606), .IN3(n2201), .IN4(n19584), .Q(
        n7610) );
  OA22X1 U30756 ( .IN1(n2286), .IN2(n19606), .IN3(n2200), .IN4(n19584), .Q(
        n7606) );
  OA22X1 U30757 ( .IN1(n2285), .IN2(n19605), .IN3(n2199), .IN4(n19585), .Q(
        n7598) );
  OA22X1 U30758 ( .IN1(n2284), .IN2(n19605), .IN3(n2198), .IN4(n19585), .Q(
        n7594) );
  OA22X1 U30759 ( .IN1(n2283), .IN2(n19604), .IN3(n2197), .IN4(n19585), .Q(
        n7590) );
  OA22X1 U30760 ( .IN1(n2282), .IN2(n19605), .IN3(n2196), .IN4(n19586), .Q(
        n7586) );
  OA22X1 U30761 ( .IN1(n2281), .IN2(n19607), .IN3(n2195), .IN4(n19586), .Q(
        n7582) );
  OA22X1 U30762 ( .IN1(n2280), .IN2(n19607), .IN3(n2194), .IN4(n19586), .Q(
        n7578) );
  OA22X1 U30763 ( .IN1(n2279), .IN2(n19607), .IN3(n2193), .IN4(n19587), .Q(
        n7574) );
  OA22X1 U30764 ( .IN1(n2278), .IN2(n19607), .IN3(n2192), .IN4(n19587), .Q(
        n7570) );
  OA22X1 U30765 ( .IN1(n2257), .IN2(n19609), .IN3(n2171), .IN4(n19589), .Q(
        n7518) );
  OA22X1 U30766 ( .IN1(n2256), .IN2(n19607), .IN3(n2170), .IN4(n19591), .Q(
        n7474) );
  OA22X1 U30767 ( .IN1(n2255), .IN2(n19610), .IN3(n2169), .IN4(n19581), .Q(
        n7430) );
  OA22X1 U30768 ( .IN1(n2254), .IN2(n19609), .IN3(n2168), .IN4(n19595), .Q(
        n7418) );
  OA22X1 U30769 ( .IN1(n2253), .IN2(n19611), .IN3(n2167), .IN4(n19595), .Q(
        n7414) );
  OA22X1 U30770 ( .IN1(n2252), .IN2(n19606), .IN3(n2166), .IN4(n19595), .Q(
        n7410) );
  OA22X1 U30771 ( .IN1(n2251), .IN2(n19610), .IN3(n2165), .IN4(n19596), .Q(
        n7406) );
  OA22X1 U30772 ( .IN1(n2250), .IN2(n19610), .IN3(n2164), .IN4(n19596), .Q(
        n7402) );
  OA22X1 U30773 ( .IN1(n2249), .IN2(n19610), .IN3(n2163), .IN4(n19596), .Q(
        n7398) );
  OA22X1 U30774 ( .IN1(n2248), .IN2(n19610), .IN3(n2162), .IN4(n19597), .Q(
        n7394) );
  OA22X1 U30775 ( .IN1(n2247), .IN2(n19609), .IN3(n2161), .IN4(n19590), .Q(
        n7514) );
  OA22X1 U30776 ( .IN1(n2246), .IN2(n19609), .IN3(n2160), .IN4(n19590), .Q(
        n7510) );
  OA22X1 U30777 ( .IN1(n2245), .IN2(n19609), .IN3(n2159), .IN4(n19590), .Q(
        n7506) );
  OA22X1 U30778 ( .IN1(n2244), .IN2(n19606), .IN3(n2158), .IN4(n19591), .Q(
        n7502) );
  OA22X1 U30779 ( .IN1(n2243), .IN2(n19605), .IN3(n2157), .IN4(n19591), .Q(
        n7498) );
  OA22X1 U30780 ( .IN1(n2242), .IN2(n19610), .IN3(n2156), .IN4(n19591), .Q(
        n7494) );
  OA22X1 U30781 ( .IN1(n2241), .IN2(n19607), .IN3(n2155), .IN4(n19594), .Q(
        n7490) );
  OA22X1 U30782 ( .IN1(n2240), .IN2(n19611), .IN3(n2154), .IN4(n19595), .Q(
        n7486) );
  OA22X1 U30783 ( .IN1(n2239), .IN2(n19609), .IN3(n2153), .IN4(n19597), .Q(
        n7482) );
  OA22X1 U30784 ( .IN1(n2238), .IN2(n19604), .IN3(n2152), .IN4(n19592), .Q(
        n7478) );
  OA22X1 U30785 ( .IN1(n2237), .IN2(n19604), .IN3(n2151), .IN4(n19585), .Q(
        n7470) );
  OA22X1 U30786 ( .IN1(n2236), .IN2(n19606), .IN3(n2150), .IN4(n19592), .Q(
        n7466) );
  OA22X1 U30787 ( .IN1(n2235), .IN2(n19608), .IN3(n2149), .IN4(n19592), .Q(
        n7462) );
  OA22X1 U30788 ( .IN1(n2234), .IN2(n19606), .IN3(n2148), .IN4(n19592), .Q(
        n7458) );
  OA22X1 U30789 ( .IN1(n2233), .IN2(n19607), .IN3(n2147), .IN4(n19593), .Q(
        n7454) );
  OA22X1 U30790 ( .IN1(n2232), .IN2(n19611), .IN3(n2146), .IN4(n19593), .Q(
        n7450) );
  OA22X1 U30791 ( .IN1(n2231), .IN2(n19610), .IN3(n2145), .IN4(n19593), .Q(
        n7446) );
  OA22X1 U30792 ( .IN1(n2230), .IN2(n19607), .IN3(n2144), .IN4(n19594), .Q(
        n7442) );
  OA22X1 U30793 ( .IN1(n2229), .IN2(n19607), .IN3(n2143), .IN4(n19594), .Q(
        n7438) );
  OA22X1 U30794 ( .IN1(n2228), .IN2(n19611), .IN3(n2142), .IN4(n19594), .Q(
        n7434) );
  OA22X1 U30795 ( .IN1(n2227), .IN2(n19610), .IN3(n2141), .IN4(n19582), .Q(
        n7426) );
  OA22X1 U30796 ( .IN1(n2226), .IN2(n19608), .IN3(n2140), .IN4(n19583), .Q(
        n7422) );
  OA22X1 U30797 ( .IN1(n2310), .IN2(n19472), .IN3(n2224), .IN4(n19466), .Q(
        n7650) );
  OA22X1 U30798 ( .IN1(n2309), .IN2(n19479), .IN3(n2223), .IN4(n19465), .Q(
        n7686) );
  OA22X1 U30799 ( .IN1(n2308), .IN2(n19479), .IN3(n2222), .IN4(n19465), .Q(
        n7682) );
  OA22X1 U30800 ( .IN1(n2307), .IN2(n19479), .IN3(n2221), .IN4(n19466), .Q(
        n7678) );
  OA22X1 U30801 ( .IN1(n2306), .IN2(n19479), .IN3(n2220), .IN4(n19466), .Q(
        n7674) );
  OA22X1 U30802 ( .IN1(n2305), .IN2(n19472), .IN3(n2219), .IN4(n19449), .Q(
        n7942) );
  OA22X1 U30803 ( .IN1(n2304), .IN2(n19474), .IN3(n2218), .IN4(n19452), .Q(
        n7898) );
  OA22X1 U30804 ( .IN1(n2303), .IN2(n19477), .IN3(n2217), .IN4(n19455), .Q(
        n7854) );
  OA22X1 U30805 ( .IN1(n2302), .IN2(n19474), .IN3(n2216), .IN4(n19455), .Q(
        n7842) );
  OA22X1 U30806 ( .IN1(n2301), .IN2(n19477), .IN3(n2215), .IN4(n19455), .Q(
        n7838) );
  OA22X1 U30807 ( .IN1(n2300), .IN2(n19476), .IN3(n2214), .IN4(n19455), .Q(
        n7834) );
  OA22X1 U30808 ( .IN1(n2299), .IN2(n19476), .IN3(n2213), .IN4(n19455), .Q(
        n7830) );
  OA22X1 U30809 ( .IN1(n2298), .IN2(n19476), .IN3(n2212), .IN4(n19455), .Q(
        n7826) );
  OA22X1 U30810 ( .IN1(n2297), .IN2(n19476), .IN3(n2211), .IN4(n19456), .Q(
        n7822) );
  OA22X1 U30811 ( .IN1(n2296), .IN2(n19476), .IN3(n2210), .IN4(n19456), .Q(
        n7818) );
  OA22X1 U30812 ( .IN1(n2295), .IN2(n19472), .IN3(n2209), .IN4(n19449), .Q(
        n7938) );
  OA22X1 U30813 ( .IN1(n2294), .IN2(n19472), .IN3(n2208), .IN4(n19449), .Q(
        n7934) );
  OA22X1 U30814 ( .IN1(n2293), .IN2(n19472), .IN3(n2207), .IN4(n19450), .Q(
        n7930) );
  OA22X1 U30815 ( .IN1(n2292), .IN2(n19473), .IN3(n2206), .IN4(n19450), .Q(
        n7926) );
  OA22X1 U30816 ( .IN1(n2291), .IN2(n19473), .IN3(n2205), .IN4(n19450), .Q(
        n7922) );
  OA22X1 U30817 ( .IN1(n2290), .IN2(n19473), .IN3(n2204), .IN4(n19451), .Q(
        n7918) );
  OA22X1 U30818 ( .IN1(n2289), .IN2(n19473), .IN3(n2203), .IN4(n19451), .Q(
        n7914) );
  OA22X1 U30819 ( .IN1(n2288), .IN2(n19474), .IN3(n2202), .IN4(n19451), .Q(
        n7910) );
  OA22X1 U30820 ( .IN1(n2287), .IN2(n19474), .IN3(n2201), .IN4(n19452), .Q(
        n7906) );
  OA22X1 U30821 ( .IN1(n2286), .IN2(n19474), .IN3(n2200), .IN4(n19452), .Q(
        n7902) );
  OA22X1 U30822 ( .IN1(n2285), .IN2(n19473), .IN3(n2199), .IN4(n19453), .Q(
        n7894) );
  OA22X1 U30823 ( .IN1(n2284), .IN2(n19473), .IN3(n2198), .IN4(n19453), .Q(
        n7890) );
  OA22X1 U30824 ( .IN1(n2283), .IN2(n19472), .IN3(n2197), .IN4(n19453), .Q(
        n7886) );
  OA22X1 U30825 ( .IN1(n2282), .IN2(n19473), .IN3(n2196), .IN4(n19454), .Q(
        n7882) );
  OA22X1 U30826 ( .IN1(n2281), .IN2(n19475), .IN3(n2195), .IN4(n19454), .Q(
        n7878) );
  OA22X1 U30827 ( .IN1(n2280), .IN2(n19475), .IN3(n2194), .IN4(n19454), .Q(
        n7874) );
  OA22X1 U30828 ( .IN1(n2279), .IN2(n19475), .IN3(n2193), .IN4(n19454), .Q(
        n7870) );
  OA22X1 U30829 ( .IN1(n2278), .IN2(n19475), .IN3(n2192), .IN4(n19454), .Q(
        n7866) );
  OA22X1 U30830 ( .IN1(n2257), .IN2(n19477), .IN3(n2171), .IN4(n19456), .Q(
        n7814) );
  OA22X1 U30831 ( .IN1(n2256), .IN2(n19474), .IN3(n2170), .IN4(n19460), .Q(
        n7770) );
  OA22X1 U30832 ( .IN1(n2255), .IN2(n19478), .IN3(n2169), .IN4(n19464), .Q(
        n7726) );
  OA22X1 U30833 ( .IN1(n2254), .IN2(n19477), .IN3(n2168), .IN4(n19464), .Q(
        n7714) );
  OA22X1 U30834 ( .IN1(n2253), .IN2(n19479), .IN3(n2167), .IN4(n19464), .Q(
        n7710) );
  OA22X1 U30835 ( .IN1(n2252), .IN2(n19474), .IN3(n2166), .IN4(n19464), .Q(
        n7706) );
  OA22X1 U30836 ( .IN1(n2251), .IN2(n19478), .IN3(n2165), .IN4(n19466), .Q(
        n7702) );
  OA22X1 U30837 ( .IN1(n2250), .IN2(n19478), .IN3(n2164), .IN4(n19466), .Q(
        n7698) );
  OA22X1 U30838 ( .IN1(n2249), .IN2(n19478), .IN3(n2163), .IN4(n19466), .Q(
        n7694) );
  OA22X1 U30839 ( .IN1(n2248), .IN2(n19478), .IN3(n2162), .IN4(n19465), .Q(
        n7690) );
  OA22X1 U30840 ( .IN1(n2247), .IN2(n19477), .IN3(n2161), .IN4(n19457), .Q(
        n7810) );
  OA22X1 U30841 ( .IN1(n2246), .IN2(n19477), .IN3(n2160), .IN4(n19457), .Q(
        n7806) );
  OA22X1 U30842 ( .IN1(n2245), .IN2(n19477), .IN3(n2159), .IN4(n19457), .Q(
        n7802) );
  OA22X1 U30843 ( .IN1(n2244), .IN2(n19475), .IN3(n2158), .IN4(n19458), .Q(
        n7798) );
  OA22X1 U30844 ( .IN1(n2243), .IN2(n19479), .IN3(n2157), .IN4(n19458), .Q(
        n7794) );
  OA22X1 U30845 ( .IN1(n2242), .IN2(n19477), .IN3(n2156), .IN4(n19458), .Q(
        n7790) );
  OA22X1 U30846 ( .IN1(n2241), .IN2(n19472), .IN3(n2155), .IN4(n19459), .Q(
        n7786) );
  OA22X1 U30847 ( .IN1(n2240), .IN2(n19478), .IN3(n2154), .IN4(n19459), .Q(
        n7782) );
  OA22X1 U30848 ( .IN1(n2239), .IN2(n19475), .IN3(n2153), .IN4(n19459), .Q(
        n7778) );
  OA22X1 U30849 ( .IN1(n2238), .IN2(n19479), .IN3(n2152), .IN4(n19460), .Q(
        n7774) );
  OA22X1 U30850 ( .IN1(n2237), .IN2(n19472), .IN3(n2151), .IN4(n19460), .Q(
        n7766) );
  OA22X1 U30851 ( .IN1(n2236), .IN2(n19476), .IN3(n2150), .IN4(n19461), .Q(
        n7762) );
  OA22X1 U30852 ( .IN1(n2235), .IN2(n19476), .IN3(n2149), .IN4(n19461), .Q(
        n7758) );
  OA22X1 U30853 ( .IN1(n2234), .IN2(n19474), .IN3(n2148), .IN4(n19461), .Q(
        n7754) );
  OA22X1 U30854 ( .IN1(n2233), .IN2(n19475), .IN3(n2147), .IN4(n19462), .Q(
        n7750) );
  OA22X1 U30855 ( .IN1(n2232), .IN2(n19479), .IN3(n2146), .IN4(n19462), .Q(
        n7746) );
  OA22X1 U30856 ( .IN1(n2231), .IN2(n19478), .IN3(n2145), .IN4(n19462), .Q(
        n7742) );
  OA22X1 U30857 ( .IN1(n2230), .IN2(n19475), .IN3(n2144), .IN4(n19463), .Q(
        n7738) );
  OA22X1 U30858 ( .IN1(n2229), .IN2(n19475), .IN3(n2143), .IN4(n19463), .Q(
        n7734) );
  OA22X1 U30859 ( .IN1(n2228), .IN2(n19479), .IN3(n2142), .IN4(n19463), .Q(
        n7730) );
  OA22X1 U30860 ( .IN1(n2227), .IN2(n19478), .IN3(n2141), .IN4(n19465), .Q(
        n7722) );
  OA22X1 U30861 ( .IN1(n2226), .IN2(n19478), .IN3(n2140), .IN4(n19455), .Q(
        n7718) );
  OA22X1 U30862 ( .IN1(n2310), .IN2(n19340), .IN3(n2224), .IN4(n19334), .Q(
        n7946) );
  OA22X1 U30863 ( .IN1(n2309), .IN2(n19347), .IN3(n2223), .IN4(n19333), .Q(
        n7982) );
  OA22X1 U30864 ( .IN1(n2308), .IN2(n19347), .IN3(n2222), .IN4(n19333), .Q(
        n7978) );
  OA22X1 U30865 ( .IN1(n2307), .IN2(n19347), .IN3(n2221), .IN4(n19334), .Q(
        n7974) );
  OA22X1 U30866 ( .IN1(n2306), .IN2(n19347), .IN3(n2220), .IN4(n19334), .Q(
        n7970) );
  OA22X1 U30867 ( .IN1(n2305), .IN2(n19340), .IN3(n2219), .IN4(n19317), .Q(
        n8238) );
  OA22X1 U30868 ( .IN1(n2304), .IN2(n19342), .IN3(n2218), .IN4(n19320), .Q(
        n8194) );
  OA22X1 U30869 ( .IN1(n2303), .IN2(n19345), .IN3(n2217), .IN4(n19323), .Q(
        n8150) );
  OA22X1 U30870 ( .IN1(n2302), .IN2(n19342), .IN3(n2216), .IN4(n19323), .Q(
        n8138) );
  OA22X1 U30871 ( .IN1(n2301), .IN2(n19345), .IN3(n2215), .IN4(n19323), .Q(
        n8134) );
  OA22X1 U30872 ( .IN1(n2300), .IN2(n19344), .IN3(n2214), .IN4(n19323), .Q(
        n8130) );
  OA22X1 U30873 ( .IN1(n2299), .IN2(n19344), .IN3(n2213), .IN4(n19323), .Q(
        n8126) );
  OA22X1 U30874 ( .IN1(n2298), .IN2(n19344), .IN3(n2212), .IN4(n19323), .Q(
        n8122) );
  OA22X1 U30875 ( .IN1(n2297), .IN2(n19344), .IN3(n2211), .IN4(n19324), .Q(
        n8118) );
  OA22X1 U30876 ( .IN1(n2296), .IN2(n19344), .IN3(n2210), .IN4(n19324), .Q(
        n8114) );
  OA22X1 U30877 ( .IN1(n2295), .IN2(n19340), .IN3(n2209), .IN4(n19317), .Q(
        n8234) );
  OA22X1 U30878 ( .IN1(n2294), .IN2(n19340), .IN3(n2208), .IN4(n19317), .Q(
        n8230) );
  OA22X1 U30879 ( .IN1(n2293), .IN2(n19340), .IN3(n2207), .IN4(n19318), .Q(
        n8226) );
  OA22X1 U30880 ( .IN1(n2292), .IN2(n19341), .IN3(n2206), .IN4(n19318), .Q(
        n8222) );
  OA22X1 U30881 ( .IN1(n2291), .IN2(n19341), .IN3(n2205), .IN4(n19318), .Q(
        n8218) );
  OA22X1 U30882 ( .IN1(n2290), .IN2(n19341), .IN3(n2204), .IN4(n19319), .Q(
        n8214) );
  OA22X1 U30883 ( .IN1(n2289), .IN2(n19341), .IN3(n2203), .IN4(n19319), .Q(
        n8210) );
  OA22X1 U30884 ( .IN1(n2288), .IN2(n19342), .IN3(n2202), .IN4(n19319), .Q(
        n8206) );
  OA22X1 U30885 ( .IN1(n2287), .IN2(n19342), .IN3(n2201), .IN4(n19320), .Q(
        n8202) );
  OA22X1 U30886 ( .IN1(n2286), .IN2(n19342), .IN3(n2200), .IN4(n19320), .Q(
        n8198) );
  OA22X1 U30887 ( .IN1(n2285), .IN2(n19341), .IN3(n2199), .IN4(n19321), .Q(
        n8190) );
  OA22X1 U30888 ( .IN1(n2284), .IN2(n19341), .IN3(n2198), .IN4(n19321), .Q(
        n8186) );
  OA22X1 U30889 ( .IN1(n2283), .IN2(n19340), .IN3(n2197), .IN4(n19321), .Q(
        n8182) );
  OA22X1 U30890 ( .IN1(n2282), .IN2(n19341), .IN3(n2196), .IN4(n19322), .Q(
        n8178) );
  OA22X1 U30891 ( .IN1(n2281), .IN2(n19343), .IN3(n2195), .IN4(n19322), .Q(
        n8174) );
  OA22X1 U30892 ( .IN1(n2280), .IN2(n19343), .IN3(n2194), .IN4(n19322), .Q(
        n8170) );
  OA22X1 U30893 ( .IN1(n2279), .IN2(n19343), .IN3(n2193), .IN4(n19322), .Q(
        n8166) );
  OA22X1 U30894 ( .IN1(n2278), .IN2(n19343), .IN3(n2192), .IN4(n19322), .Q(
        n8162) );
  OA22X1 U30895 ( .IN1(n2257), .IN2(n19345), .IN3(n2171), .IN4(n19324), .Q(
        n8110) );
  OA22X1 U30896 ( .IN1(n2256), .IN2(n19342), .IN3(n2170), .IN4(n19328), .Q(
        n8066) );
  OA22X1 U30897 ( .IN1(n2255), .IN2(n19346), .IN3(n2169), .IN4(n19332), .Q(
        n8022) );
  OA22X1 U30898 ( .IN1(n2254), .IN2(n19345), .IN3(n2168), .IN4(n19332), .Q(
        n8010) );
  OA22X1 U30899 ( .IN1(n2253), .IN2(n19347), .IN3(n2167), .IN4(n19332), .Q(
        n8006) );
  OA22X1 U30900 ( .IN1(n2252), .IN2(n19342), .IN3(n2166), .IN4(n19332), .Q(
        n8002) );
  OA22X1 U30901 ( .IN1(n2251), .IN2(n19346), .IN3(n2165), .IN4(n19334), .Q(
        n7998) );
  OA22X1 U30902 ( .IN1(n2250), .IN2(n19346), .IN3(n2164), .IN4(n19334), .Q(
        n7994) );
  OA22X1 U30903 ( .IN1(n2249), .IN2(n19346), .IN3(n2163), .IN4(n19334), .Q(
        n7990) );
  OA22X1 U30904 ( .IN1(n2248), .IN2(n19346), .IN3(n2162), .IN4(n19333), .Q(
        n7986) );
  OA22X1 U30905 ( .IN1(n2247), .IN2(n19345), .IN3(n2161), .IN4(n19325), .Q(
        n8106) );
  OA22X1 U30906 ( .IN1(n2246), .IN2(n19345), .IN3(n2160), .IN4(n19325), .Q(
        n8102) );
  OA22X1 U30907 ( .IN1(n2245), .IN2(n19345), .IN3(n2159), .IN4(n19325), .Q(
        n8098) );
  OA22X1 U30908 ( .IN1(n2244), .IN2(n19343), .IN3(n2158), .IN4(n19326), .Q(
        n8094) );
  OA22X1 U30909 ( .IN1(n2243), .IN2(n19347), .IN3(n2157), .IN4(n19326), .Q(
        n8090) );
  OA22X1 U30910 ( .IN1(n2242), .IN2(n19345), .IN3(n2156), .IN4(n19326), .Q(
        n8086) );
  OA22X1 U30911 ( .IN1(n2241), .IN2(n19340), .IN3(n2155), .IN4(n19327), .Q(
        n8082) );
  OA22X1 U30912 ( .IN1(n2240), .IN2(n19346), .IN3(n2154), .IN4(n19327), .Q(
        n8078) );
  OA22X1 U30913 ( .IN1(n2239), .IN2(n19343), .IN3(n2153), .IN4(n19327), .Q(
        n8074) );
  OA22X1 U30914 ( .IN1(n2238), .IN2(n19347), .IN3(n2152), .IN4(n19328), .Q(
        n8070) );
  OA22X1 U30915 ( .IN1(n2237), .IN2(n19340), .IN3(n2151), .IN4(n19328), .Q(
        n8062) );
  OA22X1 U30916 ( .IN1(n2236), .IN2(n19344), .IN3(n2150), .IN4(n19329), .Q(
        n8058) );
  OA22X1 U30917 ( .IN1(n2235), .IN2(n19344), .IN3(n2149), .IN4(n19329), .Q(
        n8054) );
  OA22X1 U30918 ( .IN1(n2234), .IN2(n19342), .IN3(n2148), .IN4(n19329), .Q(
        n8050) );
  OA22X1 U30919 ( .IN1(n2233), .IN2(n19343), .IN3(n2147), .IN4(n19330), .Q(
        n8046) );
  OA22X1 U30920 ( .IN1(n2232), .IN2(n19347), .IN3(n2146), .IN4(n19330), .Q(
        n8042) );
  OA22X1 U30921 ( .IN1(n2231), .IN2(n19346), .IN3(n2145), .IN4(n19330), .Q(
        n8038) );
  OA22X1 U30922 ( .IN1(n2230), .IN2(n19343), .IN3(n2144), .IN4(n19331), .Q(
        n8034) );
  OA22X1 U30923 ( .IN1(n2229), .IN2(n19343), .IN3(n2143), .IN4(n19331), .Q(
        n8030) );
  OA22X1 U30924 ( .IN1(n2228), .IN2(n19347), .IN3(n2142), .IN4(n19331), .Q(
        n8026) );
  OA22X1 U30925 ( .IN1(n2227), .IN2(n19346), .IN3(n2141), .IN4(n19333), .Q(
        n8018) );
  OA22X1 U30926 ( .IN1(n2226), .IN2(n19346), .IN3(n2140), .IN4(n19323), .Q(
        n8014) );
  OA22X1 U30927 ( .IN1(n2310), .IN2(n19208), .IN3(n2224), .IN4(n19202), .Q(
        n8242) );
  OA22X1 U30928 ( .IN1(n2309), .IN2(n19215), .IN3(n2223), .IN4(n19201), .Q(
        n8278) );
  OA22X1 U30929 ( .IN1(n2308), .IN2(n19215), .IN3(n2222), .IN4(n19201), .Q(
        n8274) );
  OA22X1 U30930 ( .IN1(n2307), .IN2(n19215), .IN3(n2221), .IN4(n19202), .Q(
        n8270) );
  OA22X1 U30931 ( .IN1(n2306), .IN2(n19215), .IN3(n2220), .IN4(n19202), .Q(
        n8266) );
  OA22X1 U30932 ( .IN1(n2305), .IN2(n19208), .IN3(n2219), .IN4(n19185), .Q(
        n8534) );
  OA22X1 U30933 ( .IN1(n2304), .IN2(n19210), .IN3(n2218), .IN4(n19188), .Q(
        n8490) );
  OA22X1 U30934 ( .IN1(n2303), .IN2(n19213), .IN3(n2217), .IN4(n19191), .Q(
        n8446) );
  OA22X1 U30935 ( .IN1(n2302), .IN2(n19210), .IN3(n2216), .IN4(n19191), .Q(
        n8434) );
  OA22X1 U30936 ( .IN1(n2301), .IN2(n19213), .IN3(n2215), .IN4(n19191), .Q(
        n8430) );
  OA22X1 U30937 ( .IN1(n2300), .IN2(n19212), .IN3(n2214), .IN4(n19191), .Q(
        n8426) );
  OA22X1 U30938 ( .IN1(n2299), .IN2(n19212), .IN3(n2213), .IN4(n19191), .Q(
        n8422) );
  OA22X1 U30939 ( .IN1(n2298), .IN2(n19212), .IN3(n2212), .IN4(n19191), .Q(
        n8418) );
  OA22X1 U30940 ( .IN1(n2297), .IN2(n19212), .IN3(n2211), .IN4(n19192), .Q(
        n8414) );
  OA22X1 U30941 ( .IN1(n2296), .IN2(n19212), .IN3(n2210), .IN4(n19192), .Q(
        n8410) );
  OA22X1 U30942 ( .IN1(n2295), .IN2(n19208), .IN3(n2209), .IN4(n19185), .Q(
        n8530) );
  OA22X1 U30943 ( .IN1(n2294), .IN2(n19208), .IN3(n2208), .IN4(n19185), .Q(
        n8526) );
  OA22X1 U30944 ( .IN1(n2293), .IN2(n19208), .IN3(n2207), .IN4(n19186), .Q(
        n8522) );
  OA22X1 U30945 ( .IN1(n2292), .IN2(n19209), .IN3(n2206), .IN4(n19186), .Q(
        n8518) );
  OA22X1 U30946 ( .IN1(n2291), .IN2(n19209), .IN3(n2205), .IN4(n19186), .Q(
        n8514) );
  OA22X1 U30947 ( .IN1(n2290), .IN2(n19209), .IN3(n2204), .IN4(n19187), .Q(
        n8510) );
  OA22X1 U30948 ( .IN1(n2289), .IN2(n19209), .IN3(n2203), .IN4(n19187), .Q(
        n8506) );
  OA22X1 U30949 ( .IN1(n2288), .IN2(n19210), .IN3(n2202), .IN4(n19187), .Q(
        n8502) );
  OA22X1 U30950 ( .IN1(n2287), .IN2(n19210), .IN3(n2201), .IN4(n19188), .Q(
        n8498) );
  OA22X1 U30951 ( .IN1(n2286), .IN2(n19210), .IN3(n2200), .IN4(n19188), .Q(
        n8494) );
  OA22X1 U30952 ( .IN1(n2285), .IN2(n19209), .IN3(n2199), .IN4(n19189), .Q(
        n8486) );
  OA22X1 U30953 ( .IN1(n2284), .IN2(n19209), .IN3(n2198), .IN4(n19189), .Q(
        n8482) );
  OA22X1 U30954 ( .IN1(n2283), .IN2(n19208), .IN3(n2197), .IN4(n19189), .Q(
        n8478) );
  OA22X1 U30955 ( .IN1(n2282), .IN2(n19209), .IN3(n2196), .IN4(n19190), .Q(
        n8474) );
  OA22X1 U30956 ( .IN1(n2281), .IN2(n19211), .IN3(n2195), .IN4(n19190), .Q(
        n8470) );
  OA22X1 U30957 ( .IN1(n2280), .IN2(n19211), .IN3(n2194), .IN4(n19190), .Q(
        n8466) );
  OA22X1 U30958 ( .IN1(n2279), .IN2(n19211), .IN3(n2193), .IN4(n19190), .Q(
        n8462) );
  OA22X1 U30959 ( .IN1(n2278), .IN2(n19211), .IN3(n2192), .IN4(n19190), .Q(
        n8458) );
  OA22X1 U30960 ( .IN1(n2257), .IN2(n19213), .IN3(n2171), .IN4(n19192), .Q(
        n8406) );
  OA22X1 U30961 ( .IN1(n2256), .IN2(n19210), .IN3(n2170), .IN4(n19196), .Q(
        n8362) );
  OA22X1 U30962 ( .IN1(n2255), .IN2(n19214), .IN3(n2169), .IN4(n19200), .Q(
        n8318) );
  OA22X1 U30963 ( .IN1(n2254), .IN2(n19213), .IN3(n2168), .IN4(n19200), .Q(
        n8306) );
  OA22X1 U30964 ( .IN1(n2253), .IN2(n19215), .IN3(n2167), .IN4(n19200), .Q(
        n8302) );
  OA22X1 U30965 ( .IN1(n2252), .IN2(n19210), .IN3(n2166), .IN4(n19200), .Q(
        n8298) );
  OA22X1 U30966 ( .IN1(n2251), .IN2(n19214), .IN3(n2165), .IN4(n19202), .Q(
        n8294) );
  OA22X1 U30967 ( .IN1(n2250), .IN2(n19214), .IN3(n2164), .IN4(n19202), .Q(
        n8290) );
  OA22X1 U30968 ( .IN1(n2249), .IN2(n19214), .IN3(n2163), .IN4(n19202), .Q(
        n8286) );
  OA22X1 U30969 ( .IN1(n2248), .IN2(n19214), .IN3(n2162), .IN4(n19201), .Q(
        n8282) );
  OA22X1 U30970 ( .IN1(n2247), .IN2(n19213), .IN3(n2161), .IN4(n19193), .Q(
        n8402) );
  OA22X1 U30971 ( .IN1(n2246), .IN2(n19213), .IN3(n2160), .IN4(n19193), .Q(
        n8398) );
  OA22X1 U30972 ( .IN1(n2245), .IN2(n19213), .IN3(n2159), .IN4(n19193), .Q(
        n8394) );
  OA22X1 U30973 ( .IN1(n2244), .IN2(n19211), .IN3(n2158), .IN4(n19194), .Q(
        n8390) );
  OA22X1 U30974 ( .IN1(n2243), .IN2(n19215), .IN3(n2157), .IN4(n19194), .Q(
        n8386) );
  OA22X1 U30975 ( .IN1(n2242), .IN2(n19213), .IN3(n2156), .IN4(n19194), .Q(
        n8382) );
  OA22X1 U30976 ( .IN1(n2241), .IN2(n19208), .IN3(n2155), .IN4(n19195), .Q(
        n8378) );
  OA22X1 U30977 ( .IN1(n2240), .IN2(n19214), .IN3(n2154), .IN4(n19195), .Q(
        n8374) );
  OA22X1 U30978 ( .IN1(n2239), .IN2(n19211), .IN3(n2153), .IN4(n19195), .Q(
        n8370) );
  OA22X1 U30979 ( .IN1(n2238), .IN2(n19215), .IN3(n2152), .IN4(n19196), .Q(
        n8366) );
  OA22X1 U30980 ( .IN1(n2237), .IN2(n19208), .IN3(n2151), .IN4(n19196), .Q(
        n8358) );
  OA22X1 U30981 ( .IN1(n2236), .IN2(n19212), .IN3(n2150), .IN4(n19197), .Q(
        n8354) );
  OA22X1 U30982 ( .IN1(n2235), .IN2(n19212), .IN3(n2149), .IN4(n19197), .Q(
        n8350) );
  OA22X1 U30983 ( .IN1(n2234), .IN2(n19210), .IN3(n2148), .IN4(n19197), .Q(
        n8346) );
  OA22X1 U30984 ( .IN1(n2233), .IN2(n19211), .IN3(n2147), .IN4(n19198), .Q(
        n8342) );
  OA22X1 U30985 ( .IN1(n2232), .IN2(n19215), .IN3(n2146), .IN4(n19198), .Q(
        n8338) );
  OA22X1 U30986 ( .IN1(n2231), .IN2(n19214), .IN3(n2145), .IN4(n19198), .Q(
        n8334) );
  OA22X1 U30987 ( .IN1(n2230), .IN2(n19211), .IN3(n2144), .IN4(n19199), .Q(
        n8330) );
  OA22X1 U30988 ( .IN1(n2229), .IN2(n19211), .IN3(n2143), .IN4(n19199), .Q(
        n8326) );
  OA22X1 U30989 ( .IN1(n2228), .IN2(n19215), .IN3(n2142), .IN4(n19199), .Q(
        n8322) );
  OA22X1 U30990 ( .IN1(n2227), .IN2(n19214), .IN3(n2141), .IN4(n19201), .Q(
        n8314) );
  OA22X1 U30991 ( .IN1(n2226), .IN2(n19214), .IN3(n2140), .IN4(n19191), .Q(
        n8310) );
  OA22X1 U30992 ( .IN1(n2310), .IN2(n19076), .IN3(n2224), .IN4(n19070), .Q(
        n8538) );
  OA22X1 U30993 ( .IN1(n2309), .IN2(n19083), .IN3(n2223), .IN4(n19069), .Q(
        n8574) );
  OA22X1 U30994 ( .IN1(n2308), .IN2(n19083), .IN3(n2222), .IN4(n19069), .Q(
        n8570) );
  OA22X1 U30995 ( .IN1(n2307), .IN2(n19083), .IN3(n2221), .IN4(n19070), .Q(
        n8566) );
  OA22X1 U30996 ( .IN1(n2306), .IN2(n19083), .IN3(n2220), .IN4(n19070), .Q(
        n8562) );
  OA22X1 U30997 ( .IN1(n2305), .IN2(n19076), .IN3(n2219), .IN4(n19053), .Q(
        n8830) );
  OA22X1 U30998 ( .IN1(n2304), .IN2(n19078), .IN3(n2218), .IN4(n19056), .Q(
        n8786) );
  OA22X1 U30999 ( .IN1(n2303), .IN2(n19082), .IN3(n2217), .IN4(n19059), .Q(
        n8742) );
  OA22X1 U31000 ( .IN1(n2302), .IN2(n8539), .IN3(n2216), .IN4(n19059), .Q(
        n8730) );
  OA22X1 U31001 ( .IN1(n2301), .IN2(n19079), .IN3(n2215), .IN4(n19059), .Q(
        n8726) );
  OA22X1 U31002 ( .IN1(n2300), .IN2(n8539), .IN3(n2214), .IN4(n19059), .Q(
        n8722) );
  OA22X1 U31003 ( .IN1(n2299), .IN2(n19080), .IN3(n2213), .IN4(n19059), .Q(
        n8718) );
  OA22X1 U31004 ( .IN1(n2298), .IN2(n19080), .IN3(n2212), .IN4(n19059), .Q(
        n8714) );
  OA22X1 U31005 ( .IN1(n2297), .IN2(n19080), .IN3(n2211), .IN4(n19060), .Q(
        n8710) );
  OA22X1 U31006 ( .IN1(n2296), .IN2(n19080), .IN3(n2210), .IN4(n19060), .Q(
        n8706) );
  OA22X1 U31007 ( .IN1(n2295), .IN2(n19076), .IN3(n2209), .IN4(n19053), .Q(
        n8826) );
  OA22X1 U31008 ( .IN1(n2294), .IN2(n19076), .IN3(n2208), .IN4(n19053), .Q(
        n8822) );
  OA22X1 U31009 ( .IN1(n2293), .IN2(n19076), .IN3(n2207), .IN4(n19054), .Q(
        n8818) );
  OA22X1 U31010 ( .IN1(n2292), .IN2(n19077), .IN3(n2206), .IN4(n19054), .Q(
        n8814) );
  OA22X1 U31011 ( .IN1(n2291), .IN2(n19077), .IN3(n2205), .IN4(n19054), .Q(
        n8810) );
  OA22X1 U31012 ( .IN1(n2290), .IN2(n19077), .IN3(n2204), .IN4(n19055), .Q(
        n8806) );
  OA22X1 U31013 ( .IN1(n2289), .IN2(n19077), .IN3(n2203), .IN4(n19055), .Q(
        n8802) );
  OA22X1 U31014 ( .IN1(n2288), .IN2(n19078), .IN3(n2202), .IN4(n19055), .Q(
        n8798) );
  OA22X1 U31015 ( .IN1(n2287), .IN2(n19078), .IN3(n2201), .IN4(n19056), .Q(
        n8794) );
  OA22X1 U31016 ( .IN1(n2286), .IN2(n19078), .IN3(n2200), .IN4(n19056), .Q(
        n8790) );
  OA22X1 U31017 ( .IN1(n2285), .IN2(n19077), .IN3(n2199), .IN4(n19057), .Q(
        n8782) );
  OA22X1 U31018 ( .IN1(n2284), .IN2(n19077), .IN3(n2198), .IN4(n19057), .Q(
        n8778) );
  OA22X1 U31019 ( .IN1(n2283), .IN2(n19076), .IN3(n2197), .IN4(n19057), .Q(
        n8774) );
  OA22X1 U31020 ( .IN1(n2282), .IN2(n19077), .IN3(n2196), .IN4(n19058), .Q(
        n8770) );
  OA22X1 U31021 ( .IN1(n2281), .IN2(n19079), .IN3(n2195), .IN4(n19058), .Q(
        n8766) );
  OA22X1 U31022 ( .IN1(n2280), .IN2(n19079), .IN3(n2194), .IN4(n19058), .Q(
        n8762) );
  OA22X1 U31023 ( .IN1(n2279), .IN2(n19079), .IN3(n2193), .IN4(n19058), .Q(
        n8758) );
  OA22X1 U31024 ( .IN1(n2278), .IN2(n19079), .IN3(n2192), .IN4(n19058), .Q(
        n8754) );
  OA22X1 U31025 ( .IN1(n2257), .IN2(n19083), .IN3(n2171), .IN4(n19060), .Q(
        n8702) );
  OA22X1 U31026 ( .IN1(n2256), .IN2(n8539), .IN3(n2170), .IN4(n19064), .Q(
        n8658) );
  OA22X1 U31027 ( .IN1(n2255), .IN2(n19082), .IN3(n2169), .IN4(n19068), .Q(
        n8614) );
  OA22X1 U31028 ( .IN1(n2254), .IN2(n8539), .IN3(n2168), .IN4(n19068), .Q(
        n8602) );
  OA22X1 U31029 ( .IN1(n2253), .IN2(n8539), .IN3(n2167), .IN4(n19068), .Q(
        n8598) );
  OA22X1 U31030 ( .IN1(n2252), .IN2(n8539), .IN3(n2166), .IN4(n19068), .Q(
        n8594) );
  OA22X1 U31031 ( .IN1(n2251), .IN2(n19082), .IN3(n2165), .IN4(n19070), .Q(
        n8590) );
  OA22X1 U31032 ( .IN1(n2250), .IN2(n19082), .IN3(n2164), .IN4(n19070), .Q(
        n8586) );
  OA22X1 U31033 ( .IN1(n2249), .IN2(n19082), .IN3(n2163), .IN4(n19070), .Q(
        n8582) );
  OA22X1 U31034 ( .IN1(n2248), .IN2(n19082), .IN3(n2162), .IN4(n19069), .Q(
        n8578) );
  OA22X1 U31035 ( .IN1(n2247), .IN2(n8539), .IN3(n2161), .IN4(n19061), .Q(
        n8698) );
  OA22X1 U31036 ( .IN1(n2246), .IN2(n19080), .IN3(n2160), .IN4(n19061), .Q(
        n8694) );
  OA22X1 U31037 ( .IN1(n2245), .IN2(n19078), .IN3(n2159), .IN4(n19061), .Q(
        n8690) );
  OA22X1 U31038 ( .IN1(n2244), .IN2(n19081), .IN3(n2158), .IN4(n19062), .Q(
        n8686) );
  OA22X1 U31039 ( .IN1(n2243), .IN2(n19081), .IN3(n2157), .IN4(n19062), .Q(
        n8682) );
  OA22X1 U31040 ( .IN1(n2242), .IN2(n19081), .IN3(n2156), .IN4(n19062), .Q(
        n8678) );
  OA22X1 U31041 ( .IN1(n2241), .IN2(n19081), .IN3(n2155), .IN4(n19063), .Q(
        n8674) );
  OA22X1 U31042 ( .IN1(n2240), .IN2(n8539), .IN3(n2154), .IN4(n19063), .Q(
        n8670) );
  OA22X1 U31043 ( .IN1(n2239), .IN2(n8539), .IN3(n2153), .IN4(n19063), .Q(
        n8666) );
  OA22X1 U31044 ( .IN1(n2238), .IN2(n8539), .IN3(n2152), .IN4(n19064), .Q(
        n8662) );
  OA22X1 U31045 ( .IN1(n2237), .IN2(n19081), .IN3(n2151), .IN4(n19064), .Q(
        n8654) );
  OA22X1 U31046 ( .IN1(n2236), .IN2(n19079), .IN3(n2150), .IN4(n19065), .Q(
        n8650) );
  OA22X1 U31047 ( .IN1(n2235), .IN2(n19081), .IN3(n2149), .IN4(n19065), .Q(
        n8646) );
  OA22X1 U31048 ( .IN1(n2234), .IN2(n19076), .IN3(n2148), .IN4(n19065), .Q(
        n8642) );
  OA22X1 U31049 ( .IN1(n2233), .IN2(n19083), .IN3(n2147), .IN4(n19066), .Q(
        n8638) );
  OA22X1 U31050 ( .IN1(n2232), .IN2(n8539), .IN3(n2146), .IN4(n19066), .Q(
        n8634) );
  OA22X1 U31051 ( .IN1(n2231), .IN2(n19080), .IN3(n2145), .IN4(n19066), .Q(
        n8630) );
  OA22X1 U31052 ( .IN1(n2230), .IN2(n19078), .IN3(n2144), .IN4(n19067), .Q(
        n8626) );
  OA22X1 U31053 ( .IN1(n2229), .IN2(n19079), .IN3(n2143), .IN4(n19067), .Q(
        n8622) );
  OA22X1 U31054 ( .IN1(n2228), .IN2(n19083), .IN3(n2142), .IN4(n19067), .Q(
        n8618) );
  OA22X1 U31055 ( .IN1(n2227), .IN2(n19082), .IN3(n2141), .IN4(n19069), .Q(
        n8610) );
  OA22X1 U31056 ( .IN1(n2226), .IN2(n8539), .IN3(n2140), .IN4(n19059), .Q(
        n8606) );
  OA22X1 U31057 ( .IN1(n2310), .IN2(n20790), .IN3(n2224), .IN4(n20784), .Q(
        n4802) );
  OA22X1 U31058 ( .IN1(n2309), .IN2(n20797), .IN3(n2223), .IN4(n20783), .Q(
        n4838) );
  OA22X1 U31059 ( .IN1(n2308), .IN2(n20797), .IN3(n2222), .IN4(n20783), .Q(
        n4834) );
  OA22X1 U31060 ( .IN1(n2307), .IN2(n20797), .IN3(n2221), .IN4(n20784), .Q(
        n4830) );
  OA22X1 U31061 ( .IN1(n2306), .IN2(n20797), .IN3(n2220), .IN4(n20784), .Q(
        n4826) );
  OA22X1 U31062 ( .IN1(n2305), .IN2(n20790), .IN3(n2219), .IN4(n20767), .Q(
        n5094) );
  OA22X1 U31063 ( .IN1(n2304), .IN2(n20792), .IN3(n2218), .IN4(n20770), .Q(
        n5050) );
  OA22X1 U31064 ( .IN1(n2303), .IN2(n20794), .IN3(n2217), .IN4(n20773), .Q(
        n5006) );
  OA22X1 U31065 ( .IN1(n2302), .IN2(n20795), .IN3(n2216), .IN4(n20773), .Q(
        n4994) );
  OA22X1 U31066 ( .IN1(n2301), .IN2(n20793), .IN3(n2215), .IN4(n20773), .Q(
        n4990) );
  OA22X1 U31067 ( .IN1(n2300), .IN2(n20795), .IN3(n2214), .IN4(n20773), .Q(
        n4986) );
  OA22X1 U31068 ( .IN1(n2299), .IN2(n4803), .IN3(n2213), .IN4(n20773), .Q(
        n4982) );
  OA22X1 U31069 ( .IN1(n2298), .IN2(n4803), .IN3(n2212), .IN4(n20773), .Q(
        n4978) );
  OA22X1 U31070 ( .IN1(n2297), .IN2(n4803), .IN3(n2211), .IN4(n20774), .Q(
        n4974) );
  OA22X1 U31071 ( .IN1(n2296), .IN2(n4803), .IN3(n2210), .IN4(n20774), .Q(
        n4970) );
  OA22X1 U31072 ( .IN1(n2295), .IN2(n20790), .IN3(n2209), .IN4(n20767), .Q(
        n5090) );
  OA22X1 U31073 ( .IN1(n2294), .IN2(n20790), .IN3(n2208), .IN4(n20767), .Q(
        n5086) );
  OA22X1 U31074 ( .IN1(n2293), .IN2(n20790), .IN3(n2207), .IN4(n20768), .Q(
        n5082) );
  OA22X1 U31075 ( .IN1(n2292), .IN2(n20791), .IN3(n2206), .IN4(n20768), .Q(
        n5078) );
  OA22X1 U31076 ( .IN1(n2291), .IN2(n20791), .IN3(n2205), .IN4(n20768), .Q(
        n5074) );
  OA22X1 U31077 ( .IN1(n2290), .IN2(n20791), .IN3(n2204), .IN4(n20769), .Q(
        n5070) );
  OA22X1 U31078 ( .IN1(n2289), .IN2(n20791), .IN3(n2203), .IN4(n20769), .Q(
        n5066) );
  OA22X1 U31079 ( .IN1(n2288), .IN2(n20792), .IN3(n2202), .IN4(n20769), .Q(
        n5062) );
  OA22X1 U31080 ( .IN1(n2287), .IN2(n20792), .IN3(n2201), .IN4(n20770), .Q(
        n5058) );
  OA22X1 U31081 ( .IN1(n2286), .IN2(n20792), .IN3(n2200), .IN4(n20770), .Q(
        n5054) );
  OA22X1 U31082 ( .IN1(n2285), .IN2(n20791), .IN3(n2199), .IN4(n20771), .Q(
        n5046) );
  OA22X1 U31083 ( .IN1(n2284), .IN2(n20791), .IN3(n2198), .IN4(n20771), .Q(
        n5042) );
  OA22X1 U31084 ( .IN1(n2283), .IN2(n20790), .IN3(n2197), .IN4(n20771), .Q(
        n5038) );
  OA22X1 U31085 ( .IN1(n2282), .IN2(n20791), .IN3(n2196), .IN4(n20772), .Q(
        n5034) );
  OA22X1 U31086 ( .IN1(n2281), .IN2(n20793), .IN3(n2195), .IN4(n20772), .Q(
        n5030) );
  OA22X1 U31087 ( .IN1(n2280), .IN2(n20793), .IN3(n2194), .IN4(n20772), .Q(
        n5026) );
  OA22X1 U31088 ( .IN1(n2279), .IN2(n20793), .IN3(n2193), .IN4(n20772), .Q(
        n5022) );
  OA22X1 U31089 ( .IN1(n2278), .IN2(n20793), .IN3(n2192), .IN4(n20772), .Q(
        n5018) );
  OA22X1 U31090 ( .IN1(n2257), .IN2(n20794), .IN3(n2171), .IN4(n20774), .Q(
        n4966) );
  OA22X1 U31091 ( .IN1(n2256), .IN2(n20795), .IN3(n2170), .IN4(n20778), .Q(
        n4922) );
  OA22X1 U31092 ( .IN1(n2255), .IN2(n20796), .IN3(n2169), .IN4(n20782), .Q(
        n4878) );
  OA22X1 U31093 ( .IN1(n2254), .IN2(n20793), .IN3(n2168), .IN4(n20782), .Q(
        n4866) );
  OA22X1 U31094 ( .IN1(n2253), .IN2(n20797), .IN3(n2167), .IN4(n20782), .Q(
        n4862) );
  OA22X1 U31095 ( .IN1(n2252), .IN2(n20791), .IN3(n2166), .IN4(n20782), .Q(
        n4858) );
  OA22X1 U31096 ( .IN1(n2251), .IN2(n20796), .IN3(n2165), .IN4(n20784), .Q(
        n4854) );
  OA22X1 U31097 ( .IN1(n2250), .IN2(n20796), .IN3(n2164), .IN4(n20784), .Q(
        n4850) );
  OA22X1 U31098 ( .IN1(n2249), .IN2(n20796), .IN3(n2163), .IN4(n20784), .Q(
        n4846) );
  OA22X1 U31099 ( .IN1(n2248), .IN2(n20796), .IN3(n2162), .IN4(n20783), .Q(
        n4842) );
  OA22X1 U31100 ( .IN1(n2247), .IN2(n20794), .IN3(n2161), .IN4(n20775), .Q(
        n4962) );
  OA22X1 U31101 ( .IN1(n2246), .IN2(n20794), .IN3(n2160), .IN4(n20775), .Q(
        n4958) );
  OA22X1 U31102 ( .IN1(n2245), .IN2(n20794), .IN3(n2159), .IN4(n20775), .Q(
        n4954) );
  OA22X1 U31103 ( .IN1(n2244), .IN2(n20792), .IN3(n2158), .IN4(n20776), .Q(
        n4950) );
  OA22X1 U31104 ( .IN1(n2243), .IN2(n20790), .IN3(n2157), .IN4(n20776), .Q(
        n4946) );
  OA22X1 U31105 ( .IN1(n2242), .IN2(n20795), .IN3(n2156), .IN4(n20776), .Q(
        n4942) );
  OA22X1 U31106 ( .IN1(n2241), .IN2(n20794), .IN3(n2155), .IN4(n20777), .Q(
        n4938) );
  OA22X1 U31107 ( .IN1(n2240), .IN2(n20795), .IN3(n2154), .IN4(n20777), .Q(
        n4934) );
  OA22X1 U31108 ( .IN1(n2239), .IN2(n20795), .IN3(n2153), .IN4(n20777), .Q(
        n4930) );
  OA22X1 U31109 ( .IN1(n2238), .IN2(n20795), .IN3(n2152), .IN4(n20778), .Q(
        n4926) );
  OA22X1 U31110 ( .IN1(n2237), .IN2(n20797), .IN3(n2151), .IN4(n20778), .Q(
        n4918) );
  OA22X1 U31111 ( .IN1(n2236), .IN2(n20790), .IN3(n2150), .IN4(n20779), .Q(
        n4914) );
  OA22X1 U31112 ( .IN1(n2235), .IN2(n20795), .IN3(n2149), .IN4(n20779), .Q(
        n4910) );
  OA22X1 U31113 ( .IN1(n2234), .IN2(n20796), .IN3(n2148), .IN4(n20779), .Q(
        n4906) );
  OA22X1 U31114 ( .IN1(n2233), .IN2(n20796), .IN3(n2147), .IN4(n20780), .Q(
        n4902) );
  OA22X1 U31115 ( .IN1(n2232), .IN2(n20793), .IN3(n2146), .IN4(n20780), .Q(
        n4898) );
  OA22X1 U31116 ( .IN1(n2231), .IN2(n20797), .IN3(n2145), .IN4(n20780), .Q(
        n4894) );
  OA22X1 U31117 ( .IN1(n2230), .IN2(n20794), .IN3(n2144), .IN4(n20781), .Q(
        n4890) );
  OA22X1 U31118 ( .IN1(n2229), .IN2(n20793), .IN3(n2143), .IN4(n20781), .Q(
        n4886) );
  OA22X1 U31119 ( .IN1(n2228), .IN2(n20797), .IN3(n2142), .IN4(n20781), .Q(
        n4882) );
  OA22X1 U31120 ( .IN1(n2227), .IN2(n20794), .IN3(n2141), .IN4(n20783), .Q(
        n4874) );
  OA22X1 U31121 ( .IN1(n2226), .IN2(n4803), .IN3(n2140), .IN4(n20773), .Q(
        n4870) );
  OA22X1 U31122 ( .IN1(n2310), .IN2(n20658), .IN3(n2224), .IN4(n20652), .Q(
        n5098) );
  OA22X1 U31123 ( .IN1(n2309), .IN2(n20665), .IN3(n2223), .IN4(n20651), .Q(
        n5134) );
  OA22X1 U31124 ( .IN1(n2308), .IN2(n20665), .IN3(n2222), .IN4(n20651), .Q(
        n5130) );
  OA22X1 U31125 ( .IN1(n2307), .IN2(n20665), .IN3(n2221), .IN4(n20652), .Q(
        n5126) );
  OA22X1 U31126 ( .IN1(n2306), .IN2(n20665), .IN3(n2220), .IN4(n20652), .Q(
        n5122) );
  OA22X1 U31127 ( .IN1(n2305), .IN2(n20658), .IN3(n2219), .IN4(n20635), .Q(
        n5390) );
  OA22X1 U31128 ( .IN1(n2304), .IN2(n20660), .IN3(n2218), .IN4(n20638), .Q(
        n5346) );
  OA22X1 U31129 ( .IN1(n2303), .IN2(n20663), .IN3(n2217), .IN4(n20642), .Q(
        n5302) );
  OA22X1 U31130 ( .IN1(n2302), .IN2(n20659), .IN3(n2216), .IN4(n20639), .Q(
        n5290) );
  OA22X1 U31131 ( .IN1(n2301), .IN2(n20663), .IN3(n2215), .IN4(n20643), .Q(
        n5286) );
  OA22X1 U31132 ( .IN1(n2300), .IN2(n20664), .IN3(n2214), .IN4(n20644), .Q(
        n5282) );
  OA22X1 U31133 ( .IN1(n2299), .IN2(n20662), .IN3(n2213), .IN4(n20645), .Q(
        n5278) );
  OA22X1 U31134 ( .IN1(n2298), .IN2(n20662), .IN3(n2212), .IN4(n20638), .Q(
        n5274) );
  OA22X1 U31135 ( .IN1(n2297), .IN2(n20662), .IN3(n2211), .IN4(n20643), .Q(
        n5270) );
  OA22X1 U31136 ( .IN1(n2296), .IN2(n20662), .IN3(n2210), .IN4(n20643), .Q(
        n5266) );
  OA22X1 U31137 ( .IN1(n2295), .IN2(n20658), .IN3(n2209), .IN4(n20635), .Q(
        n5386) );
  OA22X1 U31138 ( .IN1(n2294), .IN2(n20658), .IN3(n2208), .IN4(n20635), .Q(
        n5382) );
  OA22X1 U31139 ( .IN1(n2293), .IN2(n20658), .IN3(n2207), .IN4(n20636), .Q(
        n5378) );
  OA22X1 U31140 ( .IN1(n2292), .IN2(n20659), .IN3(n2206), .IN4(n20636), .Q(
        n5374) );
  OA22X1 U31141 ( .IN1(n2291), .IN2(n20659), .IN3(n2205), .IN4(n20636), .Q(
        n5370) );
  OA22X1 U31142 ( .IN1(n2290), .IN2(n20659), .IN3(n2204), .IN4(n20637), .Q(
        n5366) );
  OA22X1 U31143 ( .IN1(n2289), .IN2(n20659), .IN3(n2203), .IN4(n20637), .Q(
        n5362) );
  OA22X1 U31144 ( .IN1(n2288), .IN2(n20660), .IN3(n2202), .IN4(n20637), .Q(
        n5358) );
  OA22X1 U31145 ( .IN1(n2287), .IN2(n20660), .IN3(n2201), .IN4(n20638), .Q(
        n5354) );
  OA22X1 U31146 ( .IN1(n2286), .IN2(n20660), .IN3(n2200), .IN4(n20638), .Q(
        n5350) );
  OA22X1 U31147 ( .IN1(n2285), .IN2(n20659), .IN3(n2199), .IN4(n20639), .Q(
        n5342) );
  OA22X1 U31148 ( .IN1(n2284), .IN2(n20659), .IN3(n2198), .IN4(n20639), .Q(
        n5338) );
  OA22X1 U31149 ( .IN1(n2283), .IN2(n20658), .IN3(n2197), .IN4(n20639), .Q(
        n5334) );
  OA22X1 U31150 ( .IN1(n2282), .IN2(n20659), .IN3(n2196), .IN4(n20640), .Q(
        n5330) );
  OA22X1 U31151 ( .IN1(n2281), .IN2(n20661), .IN3(n2195), .IN4(n20640), .Q(
        n5326) );
  OA22X1 U31152 ( .IN1(n2280), .IN2(n20661), .IN3(n2194), .IN4(n20640), .Q(
        n5322) );
  OA22X1 U31153 ( .IN1(n2279), .IN2(n20661), .IN3(n2193), .IN4(n20641), .Q(
        n5318) );
  OA22X1 U31154 ( .IN1(n2278), .IN2(n20661), .IN3(n2192), .IN4(n20641), .Q(
        n5314) );
  OA22X1 U31155 ( .IN1(n2257), .IN2(n20663), .IN3(n2171), .IN4(n20643), .Q(
        n5262) );
  OA22X1 U31156 ( .IN1(n2256), .IN2(n20661), .IN3(n2170), .IN4(n20645), .Q(
        n5218) );
  OA22X1 U31157 ( .IN1(n2255), .IN2(n20664), .IN3(n2169), .IN4(n20649), .Q(
        n5174) );
  OA22X1 U31158 ( .IN1(n2254), .IN2(n20663), .IN3(n2168), .IN4(n20649), .Q(
        n5162) );
  OA22X1 U31159 ( .IN1(n2253), .IN2(n20665), .IN3(n2167), .IN4(n20649), .Q(
        n5158) );
  OA22X1 U31160 ( .IN1(n2252), .IN2(n20660), .IN3(n2166), .IN4(n20649), .Q(
        n5154) );
  OA22X1 U31161 ( .IN1(n2251), .IN2(n20664), .IN3(n2165), .IN4(n20650), .Q(
        n5150) );
  OA22X1 U31162 ( .IN1(n2250), .IN2(n20664), .IN3(n2164), .IN4(n20650), .Q(
        n5146) );
  OA22X1 U31163 ( .IN1(n2249), .IN2(n20664), .IN3(n2163), .IN4(n20650), .Q(
        n5142) );
  OA22X1 U31164 ( .IN1(n2248), .IN2(n20664), .IN3(n2162), .IN4(n20651), .Q(
        n5138) );
  OA22X1 U31165 ( .IN1(n2247), .IN2(n20663), .IN3(n2161), .IN4(n20644), .Q(
        n5258) );
  OA22X1 U31166 ( .IN1(n2246), .IN2(n20663), .IN3(n2160), .IN4(n20644), .Q(
        n5254) );
  OA22X1 U31167 ( .IN1(n2245), .IN2(n20663), .IN3(n2159), .IN4(n20644), .Q(
        n5250) );
  OA22X1 U31168 ( .IN1(n2244), .IN2(n20660), .IN3(n2158), .IN4(n20645), .Q(
        n5246) );
  OA22X1 U31169 ( .IN1(n2243), .IN2(n20659), .IN3(n2157), .IN4(n20645), .Q(
        n5242) );
  OA22X1 U31170 ( .IN1(n2242), .IN2(n20664), .IN3(n2156), .IN4(n20645), .Q(
        n5238) );
  OA22X1 U31171 ( .IN1(n2241), .IN2(n20661), .IN3(n2155), .IN4(n20640), .Q(
        n5234) );
  OA22X1 U31172 ( .IN1(n2240), .IN2(n20665), .IN3(n2154), .IN4(n20634), .Q(
        n5230) );
  OA22X1 U31173 ( .IN1(n2239), .IN2(n20663), .IN3(n2153), .IN4(n20642), .Q(
        n5226) );
  OA22X1 U31174 ( .IN1(n2238), .IN2(n20658), .IN3(n2152), .IN4(n20641), .Q(
        n5222) );
  OA22X1 U31175 ( .IN1(n2237), .IN2(n20658), .IN3(n2151), .IN4(n20639), .Q(
        n5214) );
  OA22X1 U31176 ( .IN1(n2236), .IN2(n20660), .IN3(n2150), .IN4(n20646), .Q(
        n5210) );
  OA22X1 U31177 ( .IN1(n2235), .IN2(n20662), .IN3(n2149), .IN4(n20646), .Q(
        n5206) );
  OA22X1 U31178 ( .IN1(n2234), .IN2(n20660), .IN3(n2148), .IN4(n20646), .Q(
        n5202) );
  OA22X1 U31179 ( .IN1(n2233), .IN2(n20661), .IN3(n2147), .IN4(n20647), .Q(
        n5198) );
  OA22X1 U31180 ( .IN1(n2232), .IN2(n20665), .IN3(n2146), .IN4(n20647), .Q(
        n5194) );
  OA22X1 U31181 ( .IN1(n2231), .IN2(n20664), .IN3(n2145), .IN4(n20647), .Q(
        n5190) );
  OA22X1 U31182 ( .IN1(n2230), .IN2(n20661), .IN3(n2144), .IN4(n20648), .Q(
        n5186) );
  OA22X1 U31183 ( .IN1(n2229), .IN2(n20661), .IN3(n2143), .IN4(n20648), .Q(
        n5182) );
  OA22X1 U31184 ( .IN1(n2228), .IN2(n20665), .IN3(n2142), .IN4(n20648), .Q(
        n5178) );
  OA22X1 U31185 ( .IN1(n2227), .IN2(n20664), .IN3(n2141), .IN4(n20651), .Q(
        n5170) );
  OA22X1 U31186 ( .IN1(n2226), .IN2(n20662), .IN3(n2140), .IN4(n20649), .Q(
        n5166) );
  OA22X1 U31187 ( .IN1(n2310), .IN2(n20526), .IN3(n2224), .IN4(n20520), .Q(
        n5394) );
  OA22X1 U31188 ( .IN1(n2309), .IN2(n20533), .IN3(n2223), .IN4(n20519), .Q(
        n5430) );
  OA22X1 U31189 ( .IN1(n2308), .IN2(n20533), .IN3(n2222), .IN4(n20519), .Q(
        n5426) );
  OA22X1 U31190 ( .IN1(n2307), .IN2(n20533), .IN3(n2221), .IN4(n20520), .Q(
        n5422) );
  OA22X1 U31191 ( .IN1(n2306), .IN2(n20533), .IN3(n2220), .IN4(n20520), .Q(
        n5418) );
  OA22X1 U31192 ( .IN1(n2305), .IN2(n20526), .IN3(n2219), .IN4(n20503), .Q(
        n5686) );
  OA22X1 U31193 ( .IN1(n2304), .IN2(n20528), .IN3(n2218), .IN4(n20506), .Q(
        n5642) );
  OA22X1 U31194 ( .IN1(n2303), .IN2(n20531), .IN3(n2217), .IN4(n20510), .Q(
        n5598) );
  OA22X1 U31195 ( .IN1(n2302), .IN2(n20527), .IN3(n2216), .IN4(n20507), .Q(
        n5586) );
  OA22X1 U31196 ( .IN1(n2301), .IN2(n20531), .IN3(n2215), .IN4(n20511), .Q(
        n5582) );
  OA22X1 U31197 ( .IN1(n2300), .IN2(n20532), .IN3(n2214), .IN4(n20512), .Q(
        n5578) );
  OA22X1 U31198 ( .IN1(n2299), .IN2(n20530), .IN3(n2213), .IN4(n20513), .Q(
        n5574) );
  OA22X1 U31199 ( .IN1(n2298), .IN2(n20530), .IN3(n2212), .IN4(n20506), .Q(
        n5570) );
  OA22X1 U31200 ( .IN1(n2297), .IN2(n20530), .IN3(n2211), .IN4(n20511), .Q(
        n5566) );
  OA22X1 U31201 ( .IN1(n2296), .IN2(n20530), .IN3(n2210), .IN4(n20511), .Q(
        n5562) );
  OA22X1 U31202 ( .IN1(n2295), .IN2(n20526), .IN3(n2209), .IN4(n20503), .Q(
        n5682) );
  OA22X1 U31203 ( .IN1(n2294), .IN2(n20526), .IN3(n2208), .IN4(n20503), .Q(
        n5678) );
  OA22X1 U31204 ( .IN1(n2293), .IN2(n20526), .IN3(n2207), .IN4(n20504), .Q(
        n5674) );
  OA22X1 U31205 ( .IN1(n2292), .IN2(n20527), .IN3(n2206), .IN4(n20504), .Q(
        n5670) );
  OA22X1 U31206 ( .IN1(n2291), .IN2(n20527), .IN3(n2205), .IN4(n20504), .Q(
        n5666) );
  OA22X1 U31207 ( .IN1(n2290), .IN2(n20527), .IN3(n2204), .IN4(n20505), .Q(
        n5662) );
  OA22X1 U31208 ( .IN1(n2289), .IN2(n20527), .IN3(n2203), .IN4(n20505), .Q(
        n5658) );
  OA22X1 U31209 ( .IN1(n2288), .IN2(n20528), .IN3(n2202), .IN4(n20505), .Q(
        n5654) );
  OA22X1 U31210 ( .IN1(n2287), .IN2(n20528), .IN3(n2201), .IN4(n20506), .Q(
        n5650) );
  OA22X1 U31211 ( .IN1(n2286), .IN2(n20528), .IN3(n2200), .IN4(n20506), .Q(
        n5646) );
  OA22X1 U31212 ( .IN1(n2285), .IN2(n20527), .IN3(n2199), .IN4(n20507), .Q(
        n5638) );
  OA22X1 U31213 ( .IN1(n2284), .IN2(n20527), .IN3(n2198), .IN4(n20507), .Q(
        n5634) );
  OA22X1 U31214 ( .IN1(n2283), .IN2(n20526), .IN3(n2197), .IN4(n20507), .Q(
        n5630) );
  OA22X1 U31215 ( .IN1(n2282), .IN2(n20527), .IN3(n2196), .IN4(n20508), .Q(
        n5626) );
  OA22X1 U31216 ( .IN1(n2281), .IN2(n20529), .IN3(n2195), .IN4(n20508), .Q(
        n5622) );
  OA22X1 U31217 ( .IN1(n2280), .IN2(n20529), .IN3(n2194), .IN4(n20508), .Q(
        n5618) );
  OA22X1 U31218 ( .IN1(n2279), .IN2(n20529), .IN3(n2193), .IN4(n20509), .Q(
        n5614) );
  OA22X1 U31219 ( .IN1(n2278), .IN2(n20529), .IN3(n2192), .IN4(n20509), .Q(
        n5610) );
  OA22X1 U31220 ( .IN1(n2257), .IN2(n20531), .IN3(n2171), .IN4(n20511), .Q(
        n5558) );
  OA22X1 U31221 ( .IN1(n2256), .IN2(n20529), .IN3(n2170), .IN4(n20513), .Q(
        n5514) );
  OA22X1 U31222 ( .IN1(n2255), .IN2(n20532), .IN3(n2169), .IN4(n20517), .Q(
        n5470) );
  OA22X1 U31223 ( .IN1(n2254), .IN2(n20531), .IN3(n2168), .IN4(n20517), .Q(
        n5458) );
  OA22X1 U31224 ( .IN1(n2253), .IN2(n20533), .IN3(n2167), .IN4(n20517), .Q(
        n5454) );
  OA22X1 U31225 ( .IN1(n2252), .IN2(n20528), .IN3(n2166), .IN4(n20517), .Q(
        n5450) );
  OA22X1 U31226 ( .IN1(n2251), .IN2(n20532), .IN3(n2165), .IN4(n20518), .Q(
        n5446) );
  OA22X1 U31227 ( .IN1(n2250), .IN2(n20532), .IN3(n2164), .IN4(n20518), .Q(
        n5442) );
  OA22X1 U31228 ( .IN1(n2249), .IN2(n20532), .IN3(n2163), .IN4(n20518), .Q(
        n5438) );
  OA22X1 U31229 ( .IN1(n2248), .IN2(n20532), .IN3(n2162), .IN4(n20519), .Q(
        n5434) );
  OA22X1 U31230 ( .IN1(n2247), .IN2(n20531), .IN3(n2161), .IN4(n20512), .Q(
        n5554) );
  OA22X1 U31231 ( .IN1(n2246), .IN2(n20531), .IN3(n2160), .IN4(n20512), .Q(
        n5550) );
  OA22X1 U31232 ( .IN1(n2245), .IN2(n20531), .IN3(n2159), .IN4(n20512), .Q(
        n5546) );
  OA22X1 U31233 ( .IN1(n2244), .IN2(n20528), .IN3(n2158), .IN4(n20513), .Q(
        n5542) );
  OA22X1 U31234 ( .IN1(n2243), .IN2(n20527), .IN3(n2157), .IN4(n20513), .Q(
        n5538) );
  OA22X1 U31235 ( .IN1(n2242), .IN2(n20532), .IN3(n2156), .IN4(n20513), .Q(
        n5534) );
  OA22X1 U31236 ( .IN1(n2241), .IN2(n20529), .IN3(n2155), .IN4(n20508), .Q(
        n5530) );
  OA22X1 U31237 ( .IN1(n2240), .IN2(n20533), .IN3(n2154), .IN4(n20502), .Q(
        n5526) );
  OA22X1 U31238 ( .IN1(n2239), .IN2(n20531), .IN3(n2153), .IN4(n20510), .Q(
        n5522) );
  OA22X1 U31239 ( .IN1(n2238), .IN2(n20526), .IN3(n2152), .IN4(n20509), .Q(
        n5518) );
  OA22X1 U31240 ( .IN1(n2237), .IN2(n20526), .IN3(n2151), .IN4(n20507), .Q(
        n5510) );
  OA22X1 U31241 ( .IN1(n2236), .IN2(n20528), .IN3(n2150), .IN4(n20514), .Q(
        n5506) );
  OA22X1 U31242 ( .IN1(n2235), .IN2(n20530), .IN3(n2149), .IN4(n20514), .Q(
        n5502) );
  OA22X1 U31243 ( .IN1(n2234), .IN2(n20528), .IN3(n2148), .IN4(n20514), .Q(
        n5498) );
  OA22X1 U31244 ( .IN1(n2233), .IN2(n20529), .IN3(n2147), .IN4(n20515), .Q(
        n5494) );
  OA22X1 U31245 ( .IN1(n2232), .IN2(n20533), .IN3(n2146), .IN4(n20515), .Q(
        n5490) );
  OA22X1 U31246 ( .IN1(n2231), .IN2(n20532), .IN3(n2145), .IN4(n20515), .Q(
        n5486) );
  OA22X1 U31247 ( .IN1(n2230), .IN2(n20529), .IN3(n2144), .IN4(n20516), .Q(
        n5482) );
  OA22X1 U31248 ( .IN1(n2229), .IN2(n20529), .IN3(n2143), .IN4(n20516), .Q(
        n5478) );
  OA22X1 U31249 ( .IN1(n2228), .IN2(n20533), .IN3(n2142), .IN4(n20516), .Q(
        n5474) );
  OA22X1 U31250 ( .IN1(n2227), .IN2(n20532), .IN3(n2141), .IN4(n20519), .Q(
        n5466) );
  OA22X1 U31251 ( .IN1(n2226), .IN2(n20530), .IN3(n2140), .IN4(n20517), .Q(
        n5462) );
  OA22X1 U31252 ( .IN1(n2310), .IN2(n20394), .IN3(n2224), .IN4(n20388), .Q(
        n5690) );
  OA22X1 U31253 ( .IN1(n2309), .IN2(n20401), .IN3(n2223), .IN4(n20387), .Q(
        n5726) );
  OA22X1 U31254 ( .IN1(n2308), .IN2(n20401), .IN3(n2222), .IN4(n20387), .Q(
        n5722) );
  OA22X1 U31255 ( .IN1(n2307), .IN2(n20401), .IN3(n2221), .IN4(n20388), .Q(
        n5718) );
  OA22X1 U31256 ( .IN1(n2306), .IN2(n20401), .IN3(n2220), .IN4(n20388), .Q(
        n5714) );
  OA22X1 U31257 ( .IN1(n2305), .IN2(n20394), .IN3(n2219), .IN4(n20371), .Q(
        n5982) );
  OA22X1 U31258 ( .IN1(n2304), .IN2(n20396), .IN3(n2218), .IN4(n20374), .Q(
        n5938) );
  OA22X1 U31259 ( .IN1(n2303), .IN2(n20399), .IN3(n2217), .IN4(n20378), .Q(
        n5894) );
  OA22X1 U31260 ( .IN1(n2302), .IN2(n20395), .IN3(n2216), .IN4(n20375), .Q(
        n5882) );
  OA22X1 U31261 ( .IN1(n2301), .IN2(n20399), .IN3(n2215), .IN4(n20379), .Q(
        n5878) );
  OA22X1 U31262 ( .IN1(n2300), .IN2(n20400), .IN3(n2214), .IN4(n20380), .Q(
        n5874) );
  OA22X1 U31263 ( .IN1(n2299), .IN2(n20398), .IN3(n2213), .IN4(n20381), .Q(
        n5870) );
  OA22X1 U31264 ( .IN1(n2298), .IN2(n20398), .IN3(n2212), .IN4(n20374), .Q(
        n5866) );
  OA22X1 U31265 ( .IN1(n2297), .IN2(n20398), .IN3(n2211), .IN4(n20379), .Q(
        n5862) );
  OA22X1 U31266 ( .IN1(n2296), .IN2(n20398), .IN3(n2210), .IN4(n20379), .Q(
        n5858) );
  OA22X1 U31267 ( .IN1(n2295), .IN2(n20394), .IN3(n2209), .IN4(n20371), .Q(
        n5978) );
  OA22X1 U31268 ( .IN1(n2294), .IN2(n20394), .IN3(n2208), .IN4(n20371), .Q(
        n5974) );
  OA22X1 U31269 ( .IN1(n2293), .IN2(n20394), .IN3(n2207), .IN4(n20372), .Q(
        n5970) );
  OA22X1 U31270 ( .IN1(n2292), .IN2(n20395), .IN3(n2206), .IN4(n20372), .Q(
        n5966) );
  OA22X1 U31271 ( .IN1(n2291), .IN2(n20395), .IN3(n2205), .IN4(n20372), .Q(
        n5962) );
  OA22X1 U31272 ( .IN1(n2290), .IN2(n20395), .IN3(n2204), .IN4(n20373), .Q(
        n5958) );
  OA22X1 U31273 ( .IN1(n2289), .IN2(n20395), .IN3(n2203), .IN4(n20373), .Q(
        n5954) );
  OA22X1 U31274 ( .IN1(n2288), .IN2(n20396), .IN3(n2202), .IN4(n20373), .Q(
        n5950) );
  OA22X1 U31275 ( .IN1(n2287), .IN2(n20396), .IN3(n2201), .IN4(n20374), .Q(
        n5946) );
  OA22X1 U31276 ( .IN1(n2286), .IN2(n20396), .IN3(n2200), .IN4(n20374), .Q(
        n5942) );
  OA22X1 U31277 ( .IN1(n2285), .IN2(n20395), .IN3(n2199), .IN4(n20375), .Q(
        n5934) );
  OA22X1 U31278 ( .IN1(n2284), .IN2(n20395), .IN3(n2198), .IN4(n20375), .Q(
        n5930) );
  OA22X1 U31279 ( .IN1(n2283), .IN2(n20394), .IN3(n2197), .IN4(n20375), .Q(
        n5926) );
  OA22X1 U31280 ( .IN1(n2282), .IN2(n20395), .IN3(n2196), .IN4(n20376), .Q(
        n5922) );
  OA22X1 U31281 ( .IN1(n2281), .IN2(n20397), .IN3(n2195), .IN4(n20376), .Q(
        n5918) );
  OA22X1 U31282 ( .IN1(n2280), .IN2(n20397), .IN3(n2194), .IN4(n20376), .Q(
        n5914) );
  OA22X1 U31283 ( .IN1(n2279), .IN2(n20397), .IN3(n2193), .IN4(n20377), .Q(
        n5910) );
  OA22X1 U31284 ( .IN1(n2278), .IN2(n20397), .IN3(n2192), .IN4(n20377), .Q(
        n5906) );
  OA22X1 U31285 ( .IN1(n2257), .IN2(n20399), .IN3(n2171), .IN4(n20379), .Q(
        n5854) );
  OA22X1 U31286 ( .IN1(n2256), .IN2(n20397), .IN3(n2170), .IN4(n20381), .Q(
        n5810) );
  OA22X1 U31287 ( .IN1(n2255), .IN2(n20400), .IN3(n2169), .IN4(n20385), .Q(
        n5766) );
  OA22X1 U31288 ( .IN1(n2254), .IN2(n20399), .IN3(n2168), .IN4(n20385), .Q(
        n5754) );
  OA22X1 U31289 ( .IN1(n2253), .IN2(n20401), .IN3(n2167), .IN4(n20385), .Q(
        n5750) );
  OA22X1 U31290 ( .IN1(n2252), .IN2(n20396), .IN3(n2166), .IN4(n20385), .Q(
        n5746) );
  OA22X1 U31291 ( .IN1(n2251), .IN2(n20400), .IN3(n2165), .IN4(n20386), .Q(
        n5742) );
  OA22X1 U31292 ( .IN1(n2250), .IN2(n20400), .IN3(n2164), .IN4(n20386), .Q(
        n5738) );
  OA22X1 U31293 ( .IN1(n2249), .IN2(n20400), .IN3(n2163), .IN4(n20386), .Q(
        n5734) );
  OA22X1 U31294 ( .IN1(n2248), .IN2(n20400), .IN3(n2162), .IN4(n20387), .Q(
        n5730) );
  OA22X1 U31295 ( .IN1(n2247), .IN2(n20399), .IN3(n2161), .IN4(n20380), .Q(
        n5850) );
  OA22X1 U31296 ( .IN1(n2246), .IN2(n20399), .IN3(n2160), .IN4(n20380), .Q(
        n5846) );
  OA22X1 U31297 ( .IN1(n2245), .IN2(n20399), .IN3(n2159), .IN4(n20380), .Q(
        n5842) );
  OA22X1 U31298 ( .IN1(n2244), .IN2(n20396), .IN3(n2158), .IN4(n20381), .Q(
        n5838) );
  OA22X1 U31299 ( .IN1(n2243), .IN2(n20395), .IN3(n2157), .IN4(n20381), .Q(
        n5834) );
  OA22X1 U31300 ( .IN1(n2242), .IN2(n20400), .IN3(n2156), .IN4(n20381), .Q(
        n5830) );
  OA22X1 U31301 ( .IN1(n2241), .IN2(n20397), .IN3(n2155), .IN4(n20376), .Q(
        n5826) );
  OA22X1 U31302 ( .IN1(n2240), .IN2(n20401), .IN3(n2154), .IN4(n20370), .Q(
        n5822) );
  OA22X1 U31303 ( .IN1(n2239), .IN2(n20399), .IN3(n2153), .IN4(n20378), .Q(
        n5818) );
  OA22X1 U31304 ( .IN1(n2238), .IN2(n20394), .IN3(n2152), .IN4(n20377), .Q(
        n5814) );
  OA22X1 U31305 ( .IN1(n2237), .IN2(n20394), .IN3(n2151), .IN4(n20375), .Q(
        n5806) );
  OA22X1 U31306 ( .IN1(n2236), .IN2(n20396), .IN3(n2150), .IN4(n20382), .Q(
        n5802) );
  OA22X1 U31307 ( .IN1(n2235), .IN2(n20398), .IN3(n2149), .IN4(n20382), .Q(
        n5798) );
  OA22X1 U31308 ( .IN1(n2234), .IN2(n20396), .IN3(n2148), .IN4(n20382), .Q(
        n5794) );
  OA22X1 U31309 ( .IN1(n2233), .IN2(n20397), .IN3(n2147), .IN4(n20383), .Q(
        n5790) );
  OA22X1 U31310 ( .IN1(n2232), .IN2(n20401), .IN3(n2146), .IN4(n20383), .Q(
        n5786) );
  OA22X1 U31311 ( .IN1(n2231), .IN2(n20400), .IN3(n2145), .IN4(n20383), .Q(
        n5782) );
  OA22X1 U31312 ( .IN1(n2230), .IN2(n20397), .IN3(n2144), .IN4(n20384), .Q(
        n5778) );
  OA22X1 U31313 ( .IN1(n2229), .IN2(n20397), .IN3(n2143), .IN4(n20384), .Q(
        n5774) );
  OA22X1 U31314 ( .IN1(n2228), .IN2(n20401), .IN3(n2142), .IN4(n20384), .Q(
        n5770) );
  OA22X1 U31315 ( .IN1(n2227), .IN2(n20400), .IN3(n2141), .IN4(n20387), .Q(
        n5762) );
  OA22X1 U31316 ( .IN1(n2226), .IN2(n20398), .IN3(n2140), .IN4(n20385), .Q(
        n5758) );
  OA22X1 U31317 ( .IN1(n2310), .IN2(n20262), .IN3(n2224), .IN4(n20256), .Q(
        n5986) );
  OA22X1 U31318 ( .IN1(n2309), .IN2(n20269), .IN3(n2223), .IN4(n20255), .Q(
        n6022) );
  OA22X1 U31319 ( .IN1(n2308), .IN2(n20269), .IN3(n2222), .IN4(n20255), .Q(
        n6018) );
  OA22X1 U31320 ( .IN1(n2307), .IN2(n20269), .IN3(n2221), .IN4(n20256), .Q(
        n6014) );
  OA22X1 U31321 ( .IN1(n2306), .IN2(n20269), .IN3(n2220), .IN4(n20256), .Q(
        n6010) );
  OA22X1 U31322 ( .IN1(n2305), .IN2(n20262), .IN3(n2219), .IN4(n20239), .Q(
        n6278) );
  OA22X1 U31323 ( .IN1(n2304), .IN2(n20264), .IN3(n2218), .IN4(n20242), .Q(
        n6234) );
  OA22X1 U31324 ( .IN1(n2303), .IN2(n20267), .IN3(n2217), .IN4(n20246), .Q(
        n6190) );
  OA22X1 U31325 ( .IN1(n2302), .IN2(n20263), .IN3(n2216), .IN4(n20243), .Q(
        n6178) );
  OA22X1 U31326 ( .IN1(n2301), .IN2(n20267), .IN3(n2215), .IN4(n20247), .Q(
        n6174) );
  OA22X1 U31327 ( .IN1(n2300), .IN2(n20268), .IN3(n2214), .IN4(n20248), .Q(
        n6170) );
  OA22X1 U31328 ( .IN1(n2299), .IN2(n20266), .IN3(n2213), .IN4(n20249), .Q(
        n6166) );
  OA22X1 U31329 ( .IN1(n2298), .IN2(n20266), .IN3(n2212), .IN4(n20251), .Q(
        n6162) );
  OA22X1 U31330 ( .IN1(n2297), .IN2(n20266), .IN3(n2211), .IN4(n20247), .Q(
        n6158) );
  OA22X1 U31331 ( .IN1(n2296), .IN2(n20266), .IN3(n2210), .IN4(n20247), .Q(
        n6154) );
  OA22X1 U31332 ( .IN1(n2295), .IN2(n20262), .IN3(n2209), .IN4(n20239), .Q(
        n6274) );
  OA22X1 U31333 ( .IN1(n2294), .IN2(n20262), .IN3(n2208), .IN4(n20239), .Q(
        n6270) );
  OA22X1 U31334 ( .IN1(n2293), .IN2(n20262), .IN3(n2207), .IN4(n20240), .Q(
        n6266) );
  OA22X1 U31335 ( .IN1(n2292), .IN2(n20263), .IN3(n2206), .IN4(n20240), .Q(
        n6262) );
  OA22X1 U31336 ( .IN1(n2291), .IN2(n20263), .IN3(n2205), .IN4(n20240), .Q(
        n6258) );
  OA22X1 U31337 ( .IN1(n2290), .IN2(n20263), .IN3(n2204), .IN4(n20241), .Q(
        n6254) );
  OA22X1 U31338 ( .IN1(n2289), .IN2(n20263), .IN3(n2203), .IN4(n20241), .Q(
        n6250) );
  OA22X1 U31339 ( .IN1(n2288), .IN2(n20264), .IN3(n2202), .IN4(n20241), .Q(
        n6246) );
  OA22X1 U31340 ( .IN1(n2287), .IN2(n20264), .IN3(n2201), .IN4(n20242), .Q(
        n6242) );
  OA22X1 U31341 ( .IN1(n2286), .IN2(n20264), .IN3(n2200), .IN4(n20242), .Q(
        n6238) );
  OA22X1 U31342 ( .IN1(n2285), .IN2(n20263), .IN3(n2199), .IN4(n20243), .Q(
        n6230) );
  OA22X1 U31343 ( .IN1(n2284), .IN2(n20263), .IN3(n2198), .IN4(n20243), .Q(
        n6226) );
  OA22X1 U31344 ( .IN1(n2283), .IN2(n20262), .IN3(n2197), .IN4(n20243), .Q(
        n6222) );
  OA22X1 U31345 ( .IN1(n2282), .IN2(n20263), .IN3(n2196), .IN4(n20244), .Q(
        n6218) );
  OA22X1 U31346 ( .IN1(n2281), .IN2(n20265), .IN3(n2195), .IN4(n20244), .Q(
        n6214) );
  OA22X1 U31347 ( .IN1(n2280), .IN2(n20265), .IN3(n2194), .IN4(n20244), .Q(
        n6210) );
  OA22X1 U31348 ( .IN1(n2279), .IN2(n20265), .IN3(n2193), .IN4(n20245), .Q(
        n6206) );
  OA22X1 U31349 ( .IN1(n2278), .IN2(n20265), .IN3(n2192), .IN4(n20245), .Q(
        n6202) );
  OA22X1 U31350 ( .IN1(n2257), .IN2(n20267), .IN3(n2171), .IN4(n20247), .Q(
        n6150) );
  OA22X1 U31351 ( .IN1(n2256), .IN2(n20265), .IN3(n2170), .IN4(n20249), .Q(
        n6106) );
  OA22X1 U31352 ( .IN1(n2255), .IN2(n20268), .IN3(n2169), .IN4(n20239), .Q(
        n6062) );
  OA22X1 U31353 ( .IN1(n2254), .IN2(n20267), .IN3(n2168), .IN4(n20253), .Q(
        n6050) );
  OA22X1 U31354 ( .IN1(n2253), .IN2(n20269), .IN3(n2167), .IN4(n20253), .Q(
        n6046) );
  OA22X1 U31355 ( .IN1(n2252), .IN2(n20264), .IN3(n2166), .IN4(n20253), .Q(
        n6042) );
  OA22X1 U31356 ( .IN1(n2251), .IN2(n20268), .IN3(n2165), .IN4(n20254), .Q(
        n6038) );
  OA22X1 U31357 ( .IN1(n2250), .IN2(n20268), .IN3(n2164), .IN4(n20254), .Q(
        n6034) );
  OA22X1 U31358 ( .IN1(n2249), .IN2(n20268), .IN3(n2163), .IN4(n20254), .Q(
        n6030) );
  OA22X1 U31359 ( .IN1(n2248), .IN2(n20268), .IN3(n2162), .IN4(n20255), .Q(
        n6026) );
  OA22X1 U31360 ( .IN1(n2247), .IN2(n20267), .IN3(n2161), .IN4(n20248), .Q(
        n6146) );
  OA22X1 U31361 ( .IN1(n2246), .IN2(n20267), .IN3(n2160), .IN4(n20248), .Q(
        n6142) );
  OA22X1 U31362 ( .IN1(n2245), .IN2(n20267), .IN3(n2159), .IN4(n20248), .Q(
        n6138) );
  OA22X1 U31363 ( .IN1(n2244), .IN2(n20264), .IN3(n2158), .IN4(n20249), .Q(
        n6134) );
  OA22X1 U31364 ( .IN1(n2243), .IN2(n20263), .IN3(n2157), .IN4(n20249), .Q(
        n6130) );
  OA22X1 U31365 ( .IN1(n2242), .IN2(n20268), .IN3(n2156), .IN4(n20249), .Q(
        n6126) );
  OA22X1 U31366 ( .IN1(n2241), .IN2(n20265), .IN3(n2155), .IN4(n20252), .Q(
        n6122) );
  OA22X1 U31367 ( .IN1(n2240), .IN2(n20269), .IN3(n2154), .IN4(n20253), .Q(
        n6118) );
  OA22X1 U31368 ( .IN1(n2239), .IN2(n20267), .IN3(n2153), .IN4(n20255), .Q(
        n6114) );
  OA22X1 U31369 ( .IN1(n2238), .IN2(n20262), .IN3(n2152), .IN4(n20250), .Q(
        n6110) );
  OA22X1 U31370 ( .IN1(n2237), .IN2(n20262), .IN3(n2151), .IN4(n20243), .Q(
        n6102) );
  OA22X1 U31371 ( .IN1(n2236), .IN2(n20264), .IN3(n2150), .IN4(n20250), .Q(
        n6098) );
  OA22X1 U31372 ( .IN1(n2235), .IN2(n20266), .IN3(n2149), .IN4(n20250), .Q(
        n6094) );
  OA22X1 U31373 ( .IN1(n2234), .IN2(n20264), .IN3(n2148), .IN4(n20250), .Q(
        n6090) );
  OA22X1 U31374 ( .IN1(n2233), .IN2(n20265), .IN3(n2147), .IN4(n20251), .Q(
        n6086) );
  OA22X1 U31375 ( .IN1(n2232), .IN2(n20269), .IN3(n2146), .IN4(n20251), .Q(
        n6082) );
  OA22X1 U31376 ( .IN1(n2231), .IN2(n20268), .IN3(n2145), .IN4(n20251), .Q(
        n6078) );
  OA22X1 U31377 ( .IN1(n2230), .IN2(n20265), .IN3(n2144), .IN4(n20252), .Q(
        n6074) );
  OA22X1 U31378 ( .IN1(n2229), .IN2(n20265), .IN3(n2143), .IN4(n20252), .Q(
        n6070) );
  OA22X1 U31379 ( .IN1(n2228), .IN2(n20269), .IN3(n2142), .IN4(n20252), .Q(
        n6066) );
  OA22X1 U31380 ( .IN1(n2227), .IN2(n20268), .IN3(n2141), .IN4(n20240), .Q(
        n6058) );
  OA22X1 U31381 ( .IN1(n2226), .IN2(n20266), .IN3(n2140), .IN4(n20241), .Q(
        n6054) );
  OA22X1 U31382 ( .IN1(n2310), .IN2(n20130), .IN3(n2224), .IN4(n20124), .Q(
        n6282) );
  OA22X1 U31383 ( .IN1(n2309), .IN2(n20137), .IN3(n2223), .IN4(n20123), .Q(
        n6318) );
  OA22X1 U31384 ( .IN1(n2308), .IN2(n20137), .IN3(n2222), .IN4(n20123), .Q(
        n6314) );
  OA22X1 U31385 ( .IN1(n2307), .IN2(n20137), .IN3(n2221), .IN4(n20124), .Q(
        n6310) );
  OA22X1 U31386 ( .IN1(n2306), .IN2(n20137), .IN3(n2220), .IN4(n20124), .Q(
        n6306) );
  OA22X1 U31387 ( .IN1(n2305), .IN2(n20130), .IN3(n2219), .IN4(n20107), .Q(
        n6574) );
  OA22X1 U31388 ( .IN1(n2304), .IN2(n20132), .IN3(n2218), .IN4(n20110), .Q(
        n6530) );
  OA22X1 U31389 ( .IN1(n2303), .IN2(n20136), .IN3(n2217), .IN4(n20113), .Q(
        n6486) );
  OA22X1 U31390 ( .IN1(n2302), .IN2(n6283), .IN3(n2216), .IN4(n20113), .Q(
        n6474) );
  OA22X1 U31391 ( .IN1(n2301), .IN2(n20133), .IN3(n2215), .IN4(n20113), .Q(
        n6470) );
  OA22X1 U31392 ( .IN1(n2300), .IN2(n6283), .IN3(n2214), .IN4(n20113), .Q(
        n6466) );
  OA22X1 U31393 ( .IN1(n2299), .IN2(n20134), .IN3(n2213), .IN4(n20113), .Q(
        n6462) );
  OA22X1 U31394 ( .IN1(n2298), .IN2(n20134), .IN3(n2212), .IN4(n20113), .Q(
        n6458) );
  OA22X1 U31395 ( .IN1(n2297), .IN2(n20134), .IN3(n2211), .IN4(n20114), .Q(
        n6454) );
  OA22X1 U31396 ( .IN1(n2296), .IN2(n20134), .IN3(n2210), .IN4(n20114), .Q(
        n6450) );
  OA22X1 U31397 ( .IN1(n2295), .IN2(n20130), .IN3(n2209), .IN4(n20107), .Q(
        n6570) );
  OA22X1 U31398 ( .IN1(n2294), .IN2(n20130), .IN3(n2208), .IN4(n20107), .Q(
        n6566) );
  OA22X1 U31399 ( .IN1(n2293), .IN2(n20130), .IN3(n2207), .IN4(n20108), .Q(
        n6562) );
  OA22X1 U31400 ( .IN1(n2292), .IN2(n20131), .IN3(n2206), .IN4(n20108), .Q(
        n6558) );
  OA22X1 U31401 ( .IN1(n2291), .IN2(n20131), .IN3(n2205), .IN4(n20108), .Q(
        n6554) );
  OA22X1 U31402 ( .IN1(n2290), .IN2(n20131), .IN3(n2204), .IN4(n20109), .Q(
        n6550) );
  OA22X1 U31403 ( .IN1(n2289), .IN2(n20131), .IN3(n2203), .IN4(n20109), .Q(
        n6546) );
  OA22X1 U31404 ( .IN1(n2288), .IN2(n20132), .IN3(n2202), .IN4(n20109), .Q(
        n6542) );
  OA22X1 U31405 ( .IN1(n2287), .IN2(n20132), .IN3(n2201), .IN4(n20110), .Q(
        n6538) );
  OA22X1 U31406 ( .IN1(n2286), .IN2(n20132), .IN3(n2200), .IN4(n20110), .Q(
        n6534) );
  OA22X1 U31407 ( .IN1(n2285), .IN2(n20131), .IN3(n2199), .IN4(n20111), .Q(
        n6526) );
  OA22X1 U31408 ( .IN1(n2284), .IN2(n20131), .IN3(n2198), .IN4(n20111), .Q(
        n6522) );
  OA22X1 U31409 ( .IN1(n2283), .IN2(n20130), .IN3(n2197), .IN4(n20111), .Q(
        n6518) );
  OA22X1 U31410 ( .IN1(n2282), .IN2(n20131), .IN3(n2196), .IN4(n20112), .Q(
        n6514) );
  OA22X1 U31411 ( .IN1(n2281), .IN2(n20133), .IN3(n2195), .IN4(n20112), .Q(
        n6510) );
  OA22X1 U31412 ( .IN1(n2280), .IN2(n20133), .IN3(n2194), .IN4(n20112), .Q(
        n6506) );
  OA22X1 U31413 ( .IN1(n2279), .IN2(n20133), .IN3(n2193), .IN4(n20112), .Q(
        n6502) );
  OA22X1 U31414 ( .IN1(n2278), .IN2(n20133), .IN3(n2192), .IN4(n20112), .Q(
        n6498) );
  OA22X1 U31415 ( .IN1(n2257), .IN2(n20137), .IN3(n2171), .IN4(n20114), .Q(
        n6446) );
  OA22X1 U31416 ( .IN1(n2256), .IN2(n6283), .IN3(n2170), .IN4(n20118), .Q(
        n6402) );
  OA22X1 U31417 ( .IN1(n2255), .IN2(n20136), .IN3(n2169), .IN4(n20122), .Q(
        n6358) );
  OA22X1 U31418 ( .IN1(n2254), .IN2(n20136), .IN3(n2168), .IN4(n20122), .Q(
        n6346) );
  OA22X1 U31419 ( .IN1(n2253), .IN2(n20137), .IN3(n2167), .IN4(n20122), .Q(
        n6342) );
  OA22X1 U31420 ( .IN1(n2252), .IN2(n20131), .IN3(n2166), .IN4(n20122), .Q(
        n6338) );
  OA22X1 U31421 ( .IN1(n2251), .IN2(n20136), .IN3(n2165), .IN4(n20124), .Q(
        n6334) );
  OA22X1 U31422 ( .IN1(n2250), .IN2(n20136), .IN3(n2164), .IN4(n20124), .Q(
        n6330) );
  OA22X1 U31423 ( .IN1(n2249), .IN2(n20136), .IN3(n2163), .IN4(n20124), .Q(
        n6326) );
  OA22X1 U31424 ( .IN1(n2248), .IN2(n20136), .IN3(n2162), .IN4(n20123), .Q(
        n6322) );
  OA22X1 U31425 ( .IN1(n2247), .IN2(n20130), .IN3(n2161), .IN4(n20115), .Q(
        n6442) );
  OA22X1 U31426 ( .IN1(n2246), .IN2(n20134), .IN3(n2160), .IN4(n20115), .Q(
        n6438) );
  OA22X1 U31427 ( .IN1(n2245), .IN2(n20132), .IN3(n2159), .IN4(n20115), .Q(
        n6434) );
  OA22X1 U31428 ( .IN1(n2244), .IN2(n20135), .IN3(n2158), .IN4(n20116), .Q(
        n6430) );
  OA22X1 U31429 ( .IN1(n2243), .IN2(n20135), .IN3(n2157), .IN4(n20116), .Q(
        n6426) );
  OA22X1 U31430 ( .IN1(n2242), .IN2(n20135), .IN3(n2156), .IN4(n20116), .Q(
        n6422) );
  OA22X1 U31431 ( .IN1(n2241), .IN2(n20135), .IN3(n2155), .IN4(n20117), .Q(
        n6418) );
  OA22X1 U31432 ( .IN1(n2240), .IN2(n6283), .IN3(n2154), .IN4(n20117), .Q(
        n6414) );
  OA22X1 U31433 ( .IN1(n2239), .IN2(n6283), .IN3(n2153), .IN4(n20117), .Q(
        n6410) );
  OA22X1 U31434 ( .IN1(n2238), .IN2(n6283), .IN3(n2152), .IN4(n20118), .Q(
        n6406) );
  OA22X1 U31435 ( .IN1(n2237), .IN2(n20135), .IN3(n2151), .IN4(n20118), .Q(
        n6398) );
  OA22X1 U31436 ( .IN1(n2236), .IN2(n20133), .IN3(n2150), .IN4(n20119), .Q(
        n6394) );
  OA22X1 U31437 ( .IN1(n2235), .IN2(n20135), .IN3(n2149), .IN4(n20119), .Q(
        n6390) );
  OA22X1 U31438 ( .IN1(n2234), .IN2(n20130), .IN3(n2148), .IN4(n20119), .Q(
        n6386) );
  OA22X1 U31439 ( .IN1(n2233), .IN2(n20137), .IN3(n2147), .IN4(n20120), .Q(
        n6382) );
  OA22X1 U31440 ( .IN1(n2232), .IN2(n20133), .IN3(n2146), .IN4(n20120), .Q(
        n6378) );
  OA22X1 U31441 ( .IN1(n2231), .IN2(n20134), .IN3(n2145), .IN4(n20120), .Q(
        n6374) );
  OA22X1 U31442 ( .IN1(n2230), .IN2(n20132), .IN3(n2144), .IN4(n20121), .Q(
        n6370) );
  OA22X1 U31443 ( .IN1(n2229), .IN2(n20133), .IN3(n2143), .IN4(n20121), .Q(
        n6366) );
  OA22X1 U31444 ( .IN1(n2228), .IN2(n20137), .IN3(n2142), .IN4(n20121), .Q(
        n6362) );
  OA22X1 U31445 ( .IN1(n2227), .IN2(n20136), .IN3(n2141), .IN4(n20123), .Q(
        n6354) );
  OA22X1 U31446 ( .IN1(n2226), .IN2(n20135), .IN3(n2140), .IN4(n20113), .Q(
        n6350) );
  OA22X1 U31447 ( .IN1(n2310), .IN2(n19999), .IN3(n2224), .IN4(n19993), .Q(
        n6578) );
  OA22X1 U31448 ( .IN1(n2309), .IN2(n20006), .IN3(n2223), .IN4(n19992), .Q(
        n6614) );
  OA22X1 U31449 ( .IN1(n2308), .IN2(n20006), .IN3(n2222), .IN4(n19992), .Q(
        n6610) );
  OA22X1 U31450 ( .IN1(n2307), .IN2(n20006), .IN3(n2221), .IN4(n19993), .Q(
        n6606) );
  OA22X1 U31451 ( .IN1(n2306), .IN2(n20006), .IN3(n2220), .IN4(n19993), .Q(
        n6602) );
  OA22X1 U31452 ( .IN1(n2305), .IN2(n19999), .IN3(n2219), .IN4(n19976), .Q(
        n6870) );
  OA22X1 U31453 ( .IN1(n2304), .IN2(n20001), .IN3(n2218), .IN4(n19979), .Q(
        n6826) );
  OA22X1 U31454 ( .IN1(n2303), .IN2(n20003), .IN3(n2217), .IN4(n19982), .Q(
        n6782) );
  OA22X1 U31455 ( .IN1(n2302), .IN2(n20004), .IN3(n2216), .IN4(n19982), .Q(
        n6770) );
  OA22X1 U31456 ( .IN1(n2301), .IN2(n20002), .IN3(n2215), .IN4(n19982), .Q(
        n6766) );
  OA22X1 U31457 ( .IN1(n2300), .IN2(n20004), .IN3(n2214), .IN4(n19982), .Q(
        n6762) );
  OA22X1 U31458 ( .IN1(n2299), .IN2(n6579), .IN3(n2213), .IN4(n19982), .Q(
        n6758) );
  OA22X1 U31459 ( .IN1(n2298), .IN2(n6579), .IN3(n2212), .IN4(n19982), .Q(
        n6754) );
  OA22X1 U31460 ( .IN1(n2297), .IN2(n6579), .IN3(n2211), .IN4(n19983), .Q(
        n6750) );
  OA22X1 U31461 ( .IN1(n2296), .IN2(n6579), .IN3(n2210), .IN4(n19983), .Q(
        n6746) );
  OA22X1 U31462 ( .IN1(n2295), .IN2(n19999), .IN3(n2209), .IN4(n19976), .Q(
        n6866) );
  OA22X1 U31463 ( .IN1(n2294), .IN2(n19999), .IN3(n2208), .IN4(n19976), .Q(
        n6862) );
  OA22X1 U31464 ( .IN1(n2293), .IN2(n19999), .IN3(n2207), .IN4(n19977), .Q(
        n6858) );
  OA22X1 U31465 ( .IN1(n2292), .IN2(n20000), .IN3(n2206), .IN4(n19977), .Q(
        n6854) );
  OA22X1 U31466 ( .IN1(n2291), .IN2(n20000), .IN3(n2205), .IN4(n19977), .Q(
        n6850) );
  OA22X1 U31467 ( .IN1(n2290), .IN2(n20000), .IN3(n2204), .IN4(n19978), .Q(
        n6846) );
  OA22X1 U31468 ( .IN1(n2289), .IN2(n20000), .IN3(n2203), .IN4(n19978), .Q(
        n6842) );
  OA22X1 U31469 ( .IN1(n2288), .IN2(n20001), .IN3(n2202), .IN4(n19978), .Q(
        n6838) );
  OA22X1 U31470 ( .IN1(n2287), .IN2(n20001), .IN3(n2201), .IN4(n19979), .Q(
        n6834) );
  OA22X1 U31471 ( .IN1(n2286), .IN2(n20001), .IN3(n2200), .IN4(n19979), .Q(
        n6830) );
  OA22X1 U31472 ( .IN1(n2285), .IN2(n20000), .IN3(n2199), .IN4(n19980), .Q(
        n6822) );
  OA22X1 U31473 ( .IN1(n2284), .IN2(n20000), .IN3(n2198), .IN4(n19980), .Q(
        n6818) );
  OA22X1 U31474 ( .IN1(n2283), .IN2(n19999), .IN3(n2197), .IN4(n19980), .Q(
        n6814) );
  OA22X1 U31475 ( .IN1(n2282), .IN2(n20000), .IN3(n2196), .IN4(n19981), .Q(
        n6810) );
  OA22X1 U31476 ( .IN1(n2281), .IN2(n20002), .IN3(n2195), .IN4(n19981), .Q(
        n6806) );
  OA22X1 U31477 ( .IN1(n2280), .IN2(n20002), .IN3(n2194), .IN4(n19981), .Q(
        n6802) );
  OA22X1 U31478 ( .IN1(n2279), .IN2(n20002), .IN3(n2193), .IN4(n19981), .Q(
        n6798) );
  OA22X1 U31479 ( .IN1(n2278), .IN2(n20002), .IN3(n2192), .IN4(n19981), .Q(
        n6794) );
  OA22X1 U31480 ( .IN1(n2257), .IN2(n20003), .IN3(n2171), .IN4(n19983), .Q(
        n6742) );
  OA22X1 U31481 ( .IN1(n2256), .IN2(n20004), .IN3(n2170), .IN4(n19987), .Q(
        n6698) );
  OA22X1 U31482 ( .IN1(n2255), .IN2(n20005), .IN3(n2169), .IN4(n19991), .Q(
        n6654) );
  OA22X1 U31483 ( .IN1(n2254), .IN2(n20002), .IN3(n2168), .IN4(n19991), .Q(
        n6642) );
  OA22X1 U31484 ( .IN1(n2253), .IN2(n20006), .IN3(n2167), .IN4(n19991), .Q(
        n6638) );
  OA22X1 U31485 ( .IN1(n2252), .IN2(n20000), .IN3(n2166), .IN4(n19991), .Q(
        n6634) );
  OA22X1 U31486 ( .IN1(n2251), .IN2(n20005), .IN3(n2165), .IN4(n19993), .Q(
        n6630) );
  OA22X1 U31487 ( .IN1(n2250), .IN2(n20005), .IN3(n2164), .IN4(n19993), .Q(
        n6626) );
  OA22X1 U31488 ( .IN1(n2249), .IN2(n20005), .IN3(n2163), .IN4(n19993), .Q(
        n6622) );
  OA22X1 U31489 ( .IN1(n2248), .IN2(n20005), .IN3(n2162), .IN4(n19992), .Q(
        n6618) );
  OA22X1 U31490 ( .IN1(n2247), .IN2(n20003), .IN3(n2161), .IN4(n19984), .Q(
        n6738) );
  OA22X1 U31491 ( .IN1(n2246), .IN2(n20003), .IN3(n2160), .IN4(n19984), .Q(
        n6734) );
  OA22X1 U31492 ( .IN1(n2245), .IN2(n20003), .IN3(n2159), .IN4(n19984), .Q(
        n6730) );
  OA22X1 U31493 ( .IN1(n2244), .IN2(n20001), .IN3(n2158), .IN4(n19985), .Q(
        n6726) );
  OA22X1 U31494 ( .IN1(n2243), .IN2(n19999), .IN3(n2157), .IN4(n19985), .Q(
        n6722) );
  OA22X1 U31495 ( .IN1(n2242), .IN2(n20004), .IN3(n2156), .IN4(n19985), .Q(
        n6718) );
  OA22X1 U31496 ( .IN1(n2241), .IN2(n20003), .IN3(n2155), .IN4(n19986), .Q(
        n6714) );
  OA22X1 U31497 ( .IN1(n2240), .IN2(n20004), .IN3(n2154), .IN4(n19986), .Q(
        n6710) );
  OA22X1 U31498 ( .IN1(n2239), .IN2(n20004), .IN3(n2153), .IN4(n19986), .Q(
        n6706) );
  OA22X1 U31499 ( .IN1(n2238), .IN2(n20004), .IN3(n2152), .IN4(n19987), .Q(
        n6702) );
  OA22X1 U31500 ( .IN1(n2237), .IN2(n20006), .IN3(n2151), .IN4(n19987), .Q(
        n6694) );
  OA22X1 U31501 ( .IN1(n2236), .IN2(n19999), .IN3(n2150), .IN4(n19988), .Q(
        n6690) );
  OA22X1 U31502 ( .IN1(n2235), .IN2(n20004), .IN3(n2149), .IN4(n19988), .Q(
        n6686) );
  OA22X1 U31503 ( .IN1(n2234), .IN2(n20005), .IN3(n2148), .IN4(n19988), .Q(
        n6682) );
  OA22X1 U31504 ( .IN1(n2233), .IN2(n20005), .IN3(n2147), .IN4(n19989), .Q(
        n6678) );
  OA22X1 U31505 ( .IN1(n2232), .IN2(n20002), .IN3(n2146), .IN4(n19989), .Q(
        n6674) );
  OA22X1 U31506 ( .IN1(n2231), .IN2(n20006), .IN3(n2145), .IN4(n19989), .Q(
        n6670) );
  OA22X1 U31507 ( .IN1(n2230), .IN2(n20003), .IN3(n2144), .IN4(n19990), .Q(
        n6666) );
  OA22X1 U31508 ( .IN1(n2229), .IN2(n20002), .IN3(n2143), .IN4(n19990), .Q(
        n6662) );
  OA22X1 U31509 ( .IN1(n2228), .IN2(n20006), .IN3(n2142), .IN4(n19990), .Q(
        n6658) );
  OA22X1 U31510 ( .IN1(n2227), .IN2(n20003), .IN3(n2141), .IN4(n19992), .Q(
        n6650) );
  OA22X1 U31511 ( .IN1(n2226), .IN2(n6579), .IN3(n2140), .IN4(n19982), .Q(
        n6646) );
  OA22X1 U31512 ( .IN1(n2310), .IN2(n19868), .IN3(n2224), .IN4(n19862), .Q(
        n6874) );
  OA22X1 U31513 ( .IN1(n2309), .IN2(n19875), .IN3(n2223), .IN4(n19861), .Q(
        n6910) );
  OA22X1 U31514 ( .IN1(n2308), .IN2(n19875), .IN3(n2222), .IN4(n19861), .Q(
        n6906) );
  OA22X1 U31515 ( .IN1(n2307), .IN2(n19875), .IN3(n2221), .IN4(n19862), .Q(
        n6902) );
  OA22X1 U31516 ( .IN1(n2306), .IN2(n19875), .IN3(n2220), .IN4(n19862), .Q(
        n6898) );
  OA22X1 U31517 ( .IN1(n2305), .IN2(n19868), .IN3(n2219), .IN4(n19845), .Q(
        n7166) );
  OA22X1 U31518 ( .IN1(n2304), .IN2(n19870), .IN3(n2218), .IN4(n19848), .Q(
        n7122) );
  OA22X1 U31519 ( .IN1(n2303), .IN2(n19874), .IN3(n2217), .IN4(n19851), .Q(
        n7078) );
  OA22X1 U31520 ( .IN1(n2302), .IN2(n6875), .IN3(n2216), .IN4(n19851), .Q(
        n7066) );
  OA22X1 U31521 ( .IN1(n2301), .IN2(n19871), .IN3(n2215), .IN4(n19851), .Q(
        n7062) );
  OA22X1 U31522 ( .IN1(n2300), .IN2(n6875), .IN3(n2214), .IN4(n19851), .Q(
        n7058) );
  OA22X1 U31523 ( .IN1(n2299), .IN2(n19872), .IN3(n2213), .IN4(n19851), .Q(
        n7054) );
  OA22X1 U31524 ( .IN1(n2298), .IN2(n19872), .IN3(n2212), .IN4(n19851), .Q(
        n7050) );
  OA22X1 U31525 ( .IN1(n2297), .IN2(n19872), .IN3(n2211), .IN4(n19852), .Q(
        n7046) );
  OA22X1 U31526 ( .IN1(n2296), .IN2(n19872), .IN3(n2210), .IN4(n19852), .Q(
        n7042) );
  OA22X1 U31527 ( .IN1(n2295), .IN2(n19868), .IN3(n2209), .IN4(n19845), .Q(
        n7162) );
  OA22X1 U31528 ( .IN1(n2294), .IN2(n19868), .IN3(n2208), .IN4(n19845), .Q(
        n7158) );
  OA22X1 U31529 ( .IN1(n2293), .IN2(n19868), .IN3(n2207), .IN4(n19846), .Q(
        n7154) );
  OA22X1 U31530 ( .IN1(n2292), .IN2(n19869), .IN3(n2206), .IN4(n19846), .Q(
        n7150) );
  OA22X1 U31531 ( .IN1(n2291), .IN2(n19869), .IN3(n2205), .IN4(n19846), .Q(
        n7146) );
  OA22X1 U31532 ( .IN1(n2290), .IN2(n19869), .IN3(n2204), .IN4(n19847), .Q(
        n7142) );
  OA22X1 U31533 ( .IN1(n2289), .IN2(n19869), .IN3(n2203), .IN4(n19847), .Q(
        n7138) );
  OA22X1 U31534 ( .IN1(n2288), .IN2(n19870), .IN3(n2202), .IN4(n19847), .Q(
        n7134) );
  OA22X1 U31535 ( .IN1(n2287), .IN2(n19870), .IN3(n2201), .IN4(n19848), .Q(
        n7130) );
  OA22X1 U31536 ( .IN1(n2286), .IN2(n19870), .IN3(n2200), .IN4(n19848), .Q(
        n7126) );
  OA22X1 U31537 ( .IN1(n2285), .IN2(n19869), .IN3(n2199), .IN4(n19849), .Q(
        n7118) );
  OA22X1 U31538 ( .IN1(n2284), .IN2(n19869), .IN3(n2198), .IN4(n19849), .Q(
        n7114) );
  OA22X1 U31539 ( .IN1(n2283), .IN2(n19868), .IN3(n2197), .IN4(n19849), .Q(
        n7110) );
  OA22X1 U31540 ( .IN1(n2282), .IN2(n19869), .IN3(n2196), .IN4(n19850), .Q(
        n7106) );
  OA22X1 U31541 ( .IN1(n2281), .IN2(n19871), .IN3(n2195), .IN4(n19850), .Q(
        n7102) );
  OA22X1 U31542 ( .IN1(n2280), .IN2(n19871), .IN3(n2194), .IN4(n19850), .Q(
        n7098) );
  OA22X1 U31543 ( .IN1(n2279), .IN2(n19871), .IN3(n2193), .IN4(n19850), .Q(
        n7094) );
  OA22X1 U31544 ( .IN1(n2278), .IN2(n19871), .IN3(n2192), .IN4(n19850), .Q(
        n7090) );
  OA22X1 U31545 ( .IN1(n2257), .IN2(n19875), .IN3(n2171), .IN4(n19852), .Q(
        n7038) );
  OA22X1 U31546 ( .IN1(n2256), .IN2(n6875), .IN3(n2170), .IN4(n19856), .Q(
        n6994) );
  OA22X1 U31547 ( .IN1(n2255), .IN2(n19874), .IN3(n2169), .IN4(n19860), .Q(
        n6950) );
  OA22X1 U31548 ( .IN1(n2254), .IN2(n6875), .IN3(n2168), .IN4(n19860), .Q(
        n6938) );
  OA22X1 U31549 ( .IN1(n2253), .IN2(n6875), .IN3(n2167), .IN4(n19860), .Q(
        n6934) );
  OA22X1 U31550 ( .IN1(n2252), .IN2(n6875), .IN3(n2166), .IN4(n19860), .Q(
        n6930) );
  OA22X1 U31551 ( .IN1(n2251), .IN2(n19874), .IN3(n2165), .IN4(n19862), .Q(
        n6926) );
  OA22X1 U31552 ( .IN1(n2250), .IN2(n19874), .IN3(n2164), .IN4(n19862), .Q(
        n6922) );
  OA22X1 U31553 ( .IN1(n2249), .IN2(n19874), .IN3(n2163), .IN4(n19862), .Q(
        n6918) );
  OA22X1 U31554 ( .IN1(n2248), .IN2(n19874), .IN3(n2162), .IN4(n19861), .Q(
        n6914) );
  OA22X1 U31555 ( .IN1(n2247), .IN2(n6875), .IN3(n2161), .IN4(n19853), .Q(
        n7034) );
  OA22X1 U31556 ( .IN1(n2246), .IN2(n19872), .IN3(n2160), .IN4(n19853), .Q(
        n7030) );
  OA22X1 U31557 ( .IN1(n2245), .IN2(n19870), .IN3(n2159), .IN4(n19853), .Q(
        n7026) );
  OA22X1 U31558 ( .IN1(n2244), .IN2(n19873), .IN3(n2158), .IN4(n19854), .Q(
        n7022) );
  OA22X1 U31559 ( .IN1(n2243), .IN2(n19873), .IN3(n2157), .IN4(n19854), .Q(
        n7018) );
  OA22X1 U31560 ( .IN1(n2242), .IN2(n19873), .IN3(n2156), .IN4(n19854), .Q(
        n7014) );
  OA22X1 U31561 ( .IN1(n2241), .IN2(n19873), .IN3(n2155), .IN4(n19855), .Q(
        n7010) );
  OA22X1 U31562 ( .IN1(n2240), .IN2(n6875), .IN3(n2154), .IN4(n19855), .Q(
        n7006) );
  OA22X1 U31563 ( .IN1(n2239), .IN2(n6875), .IN3(n2153), .IN4(n19855), .Q(
        n7002) );
  OA22X1 U31564 ( .IN1(n2238), .IN2(n6875), .IN3(n2152), .IN4(n19856), .Q(
        n6998) );
  OA22X1 U31565 ( .IN1(n2237), .IN2(n19873), .IN3(n2151), .IN4(n19856), .Q(
        n6990) );
  OA22X1 U31566 ( .IN1(n2236), .IN2(n19871), .IN3(n2150), .IN4(n19857), .Q(
        n6986) );
  OA22X1 U31567 ( .IN1(n2235), .IN2(n19873), .IN3(n2149), .IN4(n19857), .Q(
        n6982) );
  OA22X1 U31568 ( .IN1(n2234), .IN2(n19868), .IN3(n2148), .IN4(n19857), .Q(
        n6978) );
  OA22X1 U31569 ( .IN1(n2233), .IN2(n19875), .IN3(n2147), .IN4(n19858), .Q(
        n6974) );
  OA22X1 U31570 ( .IN1(n2232), .IN2(n6875), .IN3(n2146), .IN4(n19858), .Q(
        n6970) );
  OA22X1 U31571 ( .IN1(n2231), .IN2(n19872), .IN3(n2145), .IN4(n19858), .Q(
        n6966) );
  OA22X1 U31572 ( .IN1(n2230), .IN2(n19870), .IN3(n2144), .IN4(n19859), .Q(
        n6962) );
  OA22X1 U31573 ( .IN1(n2229), .IN2(n19871), .IN3(n2143), .IN4(n19859), .Q(
        n6958) );
  OA22X1 U31574 ( .IN1(n2228), .IN2(n19875), .IN3(n2142), .IN4(n19859), .Q(
        n6954) );
  OA22X1 U31575 ( .IN1(n2227), .IN2(n19874), .IN3(n2141), .IN4(n19861), .Q(
        n6946) );
  OA22X1 U31576 ( .IN1(n2226), .IN2(n6875), .IN3(n2140), .IN4(n19851), .Q(
        n6942) );
  OA22X1 U31577 ( .IN1(n2310), .IN2(n18944), .IN3(n2224), .IN4(n18938), .Q(
        n8834) );
  OA22X1 U31578 ( .IN1(n2309), .IN2(n18951), .IN3(n2223), .IN4(n18937), .Q(
        n8870) );
  OA22X1 U31579 ( .IN1(n2308), .IN2(n18951), .IN3(n2222), .IN4(n18937), .Q(
        n8866) );
  OA22X1 U31580 ( .IN1(n2307), .IN2(n18951), .IN3(n2221), .IN4(n18938), .Q(
        n8862) );
  OA22X1 U31581 ( .IN1(n2306), .IN2(n18951), .IN3(n2220), .IN4(n18938), .Q(
        n8858) );
  OA22X1 U31582 ( .IN1(n2305), .IN2(n18944), .IN3(n2219), .IN4(n18921), .Q(
        n9126) );
  OA22X1 U31583 ( .IN1(n2304), .IN2(n18946), .IN3(n2218), .IN4(n18924), .Q(
        n9082) );
  OA22X1 U31584 ( .IN1(n2303), .IN2(n18950), .IN3(n2217), .IN4(n18927), .Q(
        n9038) );
  OA22X1 U31585 ( .IN1(n2302), .IN2(n8835), .IN3(n2216), .IN4(n18927), .Q(
        n9026) );
  OA22X1 U31586 ( .IN1(n2301), .IN2(n18947), .IN3(n2215), .IN4(n18927), .Q(
        n9022) );
  OA22X1 U31587 ( .IN1(n2300), .IN2(n8835), .IN3(n2214), .IN4(n18927), .Q(
        n9018) );
  OA22X1 U31588 ( .IN1(n2299), .IN2(n18948), .IN3(n2213), .IN4(n18927), .Q(
        n9014) );
  OA22X1 U31589 ( .IN1(n2298), .IN2(n18948), .IN3(n2212), .IN4(n18927), .Q(
        n9010) );
  OA22X1 U31590 ( .IN1(n2297), .IN2(n18948), .IN3(n2211), .IN4(n18928), .Q(
        n9006) );
  OA22X1 U31591 ( .IN1(n2296), .IN2(n18948), .IN3(n2210), .IN4(n18928), .Q(
        n9002) );
  OA22X1 U31592 ( .IN1(n2295), .IN2(n18944), .IN3(n2209), .IN4(n18921), .Q(
        n9122) );
  OA22X1 U31593 ( .IN1(n2294), .IN2(n18944), .IN3(n2208), .IN4(n18921), .Q(
        n9118) );
  OA22X1 U31594 ( .IN1(n2293), .IN2(n18944), .IN3(n2207), .IN4(n18922), .Q(
        n9114) );
  OA22X1 U31595 ( .IN1(n2292), .IN2(n18945), .IN3(n2206), .IN4(n18922), .Q(
        n9110) );
  OA22X1 U31596 ( .IN1(n2291), .IN2(n18945), .IN3(n2205), .IN4(n18922), .Q(
        n9106) );
  OA22X1 U31597 ( .IN1(n2290), .IN2(n18945), .IN3(n2204), .IN4(n18923), .Q(
        n9102) );
  OA22X1 U31598 ( .IN1(n2289), .IN2(n18945), .IN3(n2203), .IN4(n18923), .Q(
        n9098) );
  OA22X1 U31599 ( .IN1(n2288), .IN2(n18946), .IN3(n2202), .IN4(n18923), .Q(
        n9094) );
  OA22X1 U31600 ( .IN1(n2287), .IN2(n18946), .IN3(n2201), .IN4(n18924), .Q(
        n9090) );
  OA22X1 U31601 ( .IN1(n2286), .IN2(n18946), .IN3(n2200), .IN4(n18924), .Q(
        n9086) );
  OA22X1 U31602 ( .IN1(n2285), .IN2(n18945), .IN3(n2199), .IN4(n18925), .Q(
        n9078) );
  OA22X1 U31603 ( .IN1(n2284), .IN2(n18945), .IN3(n2198), .IN4(n18925), .Q(
        n9074) );
  OA22X1 U31604 ( .IN1(n2283), .IN2(n18944), .IN3(n2197), .IN4(n18925), .Q(
        n9070) );
  OA22X1 U31605 ( .IN1(n2282), .IN2(n18945), .IN3(n2196), .IN4(n18926), .Q(
        n9066) );
  OA22X1 U31606 ( .IN1(n2281), .IN2(n18947), .IN3(n2195), .IN4(n18926), .Q(
        n9062) );
  OA22X1 U31607 ( .IN1(n2280), .IN2(n18947), .IN3(n2194), .IN4(n18926), .Q(
        n9058) );
  OA22X1 U31608 ( .IN1(n2279), .IN2(n18947), .IN3(n2193), .IN4(n18926), .Q(
        n9054) );
  OA22X1 U31609 ( .IN1(n2278), .IN2(n18947), .IN3(n2192), .IN4(n18926), .Q(
        n9050) );
  OA22X1 U31610 ( .IN1(n2257), .IN2(n18951), .IN3(n2171), .IN4(n18928), .Q(
        n8998) );
  OA22X1 U31611 ( .IN1(n2256), .IN2(n8835), .IN3(n2170), .IN4(n18932), .Q(
        n8954) );
  OA22X1 U31612 ( .IN1(n2255), .IN2(n18950), .IN3(n2169), .IN4(n18936), .Q(
        n8910) );
  OA22X1 U31613 ( .IN1(n2254), .IN2(n8835), .IN3(n2168), .IN4(n18936), .Q(
        n8898) );
  OA22X1 U31614 ( .IN1(n2253), .IN2(n8835), .IN3(n2167), .IN4(n18936), .Q(
        n8894) );
  OA22X1 U31615 ( .IN1(n2252), .IN2(n8835), .IN3(n2166), .IN4(n18936), .Q(
        n8890) );
  OA22X1 U31616 ( .IN1(n2251), .IN2(n18950), .IN3(n2165), .IN4(n18938), .Q(
        n8886) );
  OA22X1 U31617 ( .IN1(n2250), .IN2(n18950), .IN3(n2164), .IN4(n18938), .Q(
        n8882) );
  OA22X1 U31618 ( .IN1(n2249), .IN2(n18950), .IN3(n2163), .IN4(n18938), .Q(
        n8878) );
  OA22X1 U31619 ( .IN1(n2248), .IN2(n18950), .IN3(n2162), .IN4(n18937), .Q(
        n8874) );
  OA22X1 U31620 ( .IN1(n2247), .IN2(n8835), .IN3(n2161), .IN4(n18929), .Q(
        n8994) );
  OA22X1 U31621 ( .IN1(n2246), .IN2(n18948), .IN3(n2160), .IN4(n18929), .Q(
        n8990) );
  OA22X1 U31622 ( .IN1(n2245), .IN2(n18946), .IN3(n2159), .IN4(n18929), .Q(
        n8986) );
  OA22X1 U31623 ( .IN1(n2244), .IN2(n18949), .IN3(n2158), .IN4(n18930), .Q(
        n8982) );
  OA22X1 U31624 ( .IN1(n2243), .IN2(n18949), .IN3(n2157), .IN4(n18930), .Q(
        n8978) );
  OA22X1 U31625 ( .IN1(n2242), .IN2(n18949), .IN3(n2156), .IN4(n18930), .Q(
        n8974) );
  OA22X1 U31626 ( .IN1(n2241), .IN2(n18949), .IN3(n2155), .IN4(n18931), .Q(
        n8970) );
  OA22X1 U31627 ( .IN1(n2240), .IN2(n8835), .IN3(n2154), .IN4(n18931), .Q(
        n8966) );
  OA22X1 U31628 ( .IN1(n2239), .IN2(n8835), .IN3(n2153), .IN4(n18931), .Q(
        n8962) );
  OA22X1 U31629 ( .IN1(n2238), .IN2(n8835), .IN3(n2152), .IN4(n18932), .Q(
        n8958) );
  OA22X1 U31630 ( .IN1(n2237), .IN2(n18949), .IN3(n2151), .IN4(n18932), .Q(
        n8950) );
  OA22X1 U31631 ( .IN1(n2236), .IN2(n18947), .IN3(n2150), .IN4(n18933), .Q(
        n8946) );
  OA22X1 U31632 ( .IN1(n2235), .IN2(n18949), .IN3(n2149), .IN4(n18933), .Q(
        n8942) );
  OA22X1 U31633 ( .IN1(n2234), .IN2(n18944), .IN3(n2148), .IN4(n18933), .Q(
        n8938) );
  OA22X1 U31634 ( .IN1(n2233), .IN2(n18951), .IN3(n2147), .IN4(n18934), .Q(
        n8934) );
  OA22X1 U31635 ( .IN1(n2232), .IN2(n8835), .IN3(n2146), .IN4(n18934), .Q(
        n8930) );
  OA22X1 U31636 ( .IN1(n2231), .IN2(n18948), .IN3(n2145), .IN4(n18934), .Q(
        n8926) );
  OA22X1 U31637 ( .IN1(n2230), .IN2(n18946), .IN3(n2144), .IN4(n18935), .Q(
        n8922) );
  OA22X1 U31638 ( .IN1(n2229), .IN2(n18947), .IN3(n2143), .IN4(n18935), .Q(
        n8918) );
  OA22X1 U31639 ( .IN1(n2228), .IN2(n18951), .IN3(n2142), .IN4(n18935), .Q(
        n8914) );
  OA22X1 U31640 ( .IN1(n2227), .IN2(n18950), .IN3(n2141), .IN4(n18937), .Q(
        n8906) );
  OA22X1 U31641 ( .IN1(n2226), .IN2(n8835), .IN3(n2140), .IN4(n18927), .Q(
        n8902) );
  OA22X1 U31642 ( .IN1(n2311), .IN2(n7367), .IN3(n2225), .IN4(n7368), .Q(n7366) );
  OA22X1 U31643 ( .IN1(n2311), .IN2(n7663), .IN3(n2225), .IN4(n7664), .Q(n7662) );
  OA22X1 U31644 ( .IN1(n2311), .IN2(n7959), .IN3(n2225), .IN4(n7960), .Q(n7958) );
  OA22X1 U31645 ( .IN1(n2311), .IN2(n8255), .IN3(n2225), .IN4(n8256), .Q(n8254) );
  OA22X1 U31646 ( .IN1(n2311), .IN2(n8551), .IN3(n2225), .IN4(n8552), .Q(n8550) );
  OA22X1 U31647 ( .IN1(n20862), .IN2(n2310), .IN3(n20858), .IN4(n2224), .Q(
        n4506) );
  OA22X1 U31648 ( .IN1(n2311), .IN2(n4815), .IN3(n2225), .IN4(n4816), .Q(n4814) );
  OA22X1 U31649 ( .IN1(n2311), .IN2(n5111), .IN3(n2225), .IN4(n5112), .Q(n5110) );
  OA22X1 U31650 ( .IN1(n2311), .IN2(n5407), .IN3(n2225), .IN4(n5408), .Q(n5406) );
  OA22X1 U31651 ( .IN1(n2311), .IN2(n5703), .IN3(n2225), .IN4(n5704), .Q(n5702) );
  OA22X1 U31652 ( .IN1(n2311), .IN2(n5999), .IN3(n2225), .IN4(n6000), .Q(n5998) );
  OA22X1 U31653 ( .IN1(n2311), .IN2(n6295), .IN3(n2225), .IN4(n6296), .Q(n6294) );
  OA22X1 U31654 ( .IN1(n2311), .IN2(n6591), .IN3(n2225), .IN4(n6592), .Q(n6590) );
  OA22X1 U31655 ( .IN1(n2311), .IN2(n6887), .IN3(n2225), .IN4(n6888), .Q(n6886) );
  OA22X1 U31656 ( .IN1(n2311), .IN2(n8847), .IN3(n2225), .IN4(n8848), .Q(n8846) );
  OA22X1 U31657 ( .IN1(n20869), .IN2(n2309), .IN3(n20860), .IN4(n2223), .Q(
        n4542) );
  OA22X1 U31658 ( .IN1(n20869), .IN2(n2308), .IN3(n20860), .IN4(n2222), .Q(
        n4538) );
  OA22X1 U31659 ( .IN1(n20869), .IN2(n2307), .IN3(n20860), .IN4(n2221), .Q(
        n4534) );
  OA22X1 U31660 ( .IN1(n20869), .IN2(n2306), .IN3(n20860), .IN4(n2220), .Q(
        n4530) );
  OA22X1 U31661 ( .IN1(n20862), .IN2(n2305), .IN3(n20853), .IN4(n2219), .Q(
        n4798) );
  OA22X1 U31662 ( .IN1(n20864), .IN2(n2304), .IN3(n20855), .IN4(n2218), .Q(
        n4754) );
  OA22X1 U31663 ( .IN1(n20864), .IN2(n2303), .IN3(n20857), .IN4(n2217), .Q(
        n4710) );
  OA22X1 U31664 ( .IN1(n20865), .IN2(n2302), .IN3(n20856), .IN4(n2216), .Q(
        n4698) );
  OA22X1 U31665 ( .IN1(n20864), .IN2(n2301), .IN3(n20856), .IN4(n2215), .Q(
        n4694) );
  OA22X1 U31666 ( .IN1(n20866), .IN2(n2300), .IN3(n20857), .IN4(n2214), .Q(
        n4690) );
  OA22X1 U31667 ( .IN1(n20865), .IN2(n2299), .IN3(n20858), .IN4(n2213), .Q(
        n4686) );
  OA22X1 U31668 ( .IN1(n20865), .IN2(n2298), .IN3(n20858), .IN4(n2212), .Q(
        n4682) );
  OA22X1 U31669 ( .IN1(n20865), .IN2(n2297), .IN3(n20858), .IN4(n2211), .Q(
        n4678) );
  OA22X1 U31670 ( .IN1(n20865), .IN2(n2296), .IN3(n20858), .IN4(n2210), .Q(
        n4674) );
  OA22X1 U31671 ( .IN1(n20862), .IN2(n2295), .IN3(n20853), .IN4(n2209), .Q(
        n4794) );
  OA22X1 U31672 ( .IN1(n20862), .IN2(n2294), .IN3(n20853), .IN4(n2208), .Q(
        n4790) );
  OA22X1 U31673 ( .IN1(n20862), .IN2(n2293), .IN3(n20853), .IN4(n2207), .Q(
        n4786) );
  OA22X1 U31674 ( .IN1(n20863), .IN2(n2292), .IN3(n20854), .IN4(n2206), .Q(
        n4782) );
  OA22X1 U31675 ( .IN1(n20863), .IN2(n2291), .IN3(n20854), .IN4(n2205), .Q(
        n4778) );
  OA22X1 U31676 ( .IN1(n20863), .IN2(n2290), .IN3(n20854), .IN4(n2204), .Q(
        n4774) );
  OA22X1 U31677 ( .IN1(n20863), .IN2(n2289), .IN3(n20854), .IN4(n2203), .Q(
        n4770) );
  OA22X1 U31678 ( .IN1(n20864), .IN2(n2288), .IN3(n20855), .IN4(n2202), .Q(
        n4766) );
  OA22X1 U31679 ( .IN1(n20864), .IN2(n2287), .IN3(n20855), .IN4(n2201), .Q(
        n4762) );
  OA22X1 U31680 ( .IN1(n20864), .IN2(n2286), .IN3(n20855), .IN4(n2200), .Q(
        n4758) );
  OA22X1 U31681 ( .IN1(n20869), .IN2(n2285), .IN3(n20860), .IN4(n2199), .Q(
        n4750) );
  OA22X1 U31682 ( .IN1(n20865), .IN2(n2284), .IN3(n20853), .IN4(n2198), .Q(
        n4746) );
  OA22X1 U31683 ( .IN1(n20866), .IN2(n2283), .IN3(n20854), .IN4(n2197), .Q(
        n4742) );
  OA22X1 U31684 ( .IN1(n20863), .IN2(n2282), .IN3(n20860), .IN4(n2196), .Q(
        n4738) );
  OA22X1 U31685 ( .IN1(n4507), .IN2(n2281), .IN3(n20856), .IN4(n2195), .Q(
        n4734) );
  OA22X1 U31686 ( .IN1(n20867), .IN2(n2280), .IN3(n20856), .IN4(n2194), .Q(
        n4730) );
  OA22X1 U31687 ( .IN1(n20868), .IN2(n2279), .IN3(n20856), .IN4(n2193), .Q(
        n4726) );
  OA22X1 U31688 ( .IN1(n20863), .IN2(n2278), .IN3(n20856), .IN4(n2192), .Q(
        n4722) );
  OA22X1 U31689 ( .IN1(n20863), .IN2(n2277), .IN3(n20857), .IN4(n2191), .Q(
        n4718) );
  OA22X1 U31690 ( .IN1(n20869), .IN2(n2276), .IN3(n20857), .IN4(n2190), .Q(
        n4714) );
  OA22X1 U31691 ( .IN1(n20869), .IN2(n2275), .IN3(n20857), .IN4(n2189), .Q(
        n4706) );
  OA22X1 U31692 ( .IN1(n4507), .IN2(n2274), .IN3(n20857), .IN4(n2188), .Q(
        n4702) );
  OA22X1 U31693 ( .IN1(n20866), .IN2(n2257), .IN3(n4508), .IN4(n2171), .Q(
        n4670) );
  OA22X1 U31694 ( .IN1(n20867), .IN2(n2256), .IN3(n4508), .IN4(n2170), .Q(
        n4626) );
  OA22X1 U31695 ( .IN1(n4507), .IN2(n2255), .IN3(n20859), .IN4(n2169), .Q(
        n4582) );
  OA22X1 U31696 ( .IN1(n20862), .IN2(n2254), .IN3(n4508), .IN4(n2168), .Q(
        n4570) );
  OA22X1 U31697 ( .IN1(n4507), .IN2(n2253), .IN3(n20855), .IN4(n2167), .Q(
        n4566) );
  OA22X1 U31698 ( .IN1(n20867), .IN2(n2252), .IN3(n20854), .IN4(n2166), .Q(
        n4562) );
  OA22X1 U31699 ( .IN1(n4507), .IN2(n2251), .IN3(n20854), .IN4(n2165), .Q(
        n4558) );
  OA22X1 U31700 ( .IN1(n4507), .IN2(n2250), .IN3(n20858), .IN4(n2164), .Q(
        n4554) );
  OA22X1 U31701 ( .IN1(n4507), .IN2(n2249), .IN3(n20860), .IN4(n2163), .Q(
        n4550) );
  OA22X1 U31702 ( .IN1(n4507), .IN2(n2248), .IN3(n20856), .IN4(n2162), .Q(
        n4546) );
  OA22X1 U31703 ( .IN1(n20866), .IN2(n2247), .IN3(n4508), .IN4(n2161), .Q(
        n4666) );
  OA22X1 U31704 ( .IN1(n20866), .IN2(n2246), .IN3(n4508), .IN4(n2160), .Q(
        n4662) );
  OA22X1 U31705 ( .IN1(n20866), .IN2(n2245), .IN3(n4508), .IN4(n2159), .Q(
        n4658) );
  OA22X1 U31706 ( .IN1(n4507), .IN2(n2244), .IN3(n20859), .IN4(n2158), .Q(
        n4654) );
  OA22X1 U31707 ( .IN1(n4507), .IN2(n2243), .IN3(n20859), .IN4(n2157), .Q(
        n4650) );
  OA22X1 U31708 ( .IN1(n4507), .IN2(n2242), .IN3(n20859), .IN4(n2156), .Q(
        n4646) );
  OA22X1 U31709 ( .IN1(n4507), .IN2(n2241), .IN3(n20859), .IN4(n2155), .Q(
        n4642) );
  OA22X1 U31710 ( .IN1(n20867), .IN2(n2240), .IN3(n4508), .IN4(n2154), .Q(
        n4638) );
  OA22X1 U31711 ( .IN1(n20867), .IN2(n2239), .IN3(n4508), .IN4(n2153), .Q(
        n4634) );
  OA22X1 U31712 ( .IN1(n20867), .IN2(n2238), .IN3(n4508), .IN4(n2152), .Q(
        n4630) );
  OA22X1 U31713 ( .IN1(n20868), .IN2(n2237), .IN3(n20855), .IN4(n2151), .Q(
        n4622) );
  OA22X1 U31714 ( .IN1(n20868), .IN2(n2236), .IN3(n20859), .IN4(n2150), .Q(
        n4618) );
  OA22X1 U31715 ( .IN1(n20868), .IN2(n2235), .IN3(n4508), .IN4(n2149), .Q(
        n4614) );
  OA22X1 U31716 ( .IN1(n20868), .IN2(n2234), .IN3(n20853), .IN4(n2148), .Q(
        n4610) );
  OA22X1 U31717 ( .IN1(n4507), .IN2(n2233), .IN3(n20855), .IN4(n2147), .Q(
        n4606) );
  OA22X1 U31718 ( .IN1(n20865), .IN2(n2232), .IN3(n20859), .IN4(n2146), .Q(
        n4602) );
  OA22X1 U31719 ( .IN1(n20864), .IN2(n2231), .IN3(n4508), .IN4(n2145), .Q(
        n4598) );
  OA22X1 U31720 ( .IN1(n20866), .IN2(n2230), .IN3(n20853), .IN4(n2144), .Q(
        n4594) );
  OA22X1 U31721 ( .IN1(n20867), .IN2(n2229), .IN3(n4508), .IN4(n2143), .Q(
        n4590) );
  OA22X1 U31722 ( .IN1(n20868), .IN2(n2228), .IN3(n20857), .IN4(n2142), .Q(
        n4586) );
  OA22X1 U31723 ( .IN1(n20862), .IN2(n2227), .IN3(n20858), .IN4(n2141), .Q(
        n4578) );
  OA22X1 U31724 ( .IN1(n20868), .IN2(n2226), .IN3(n4508), .IN4(n2140), .Q(
        n4574) );
  OA22X1 U31725 ( .IN1(n4519), .IN2(n2311), .IN3(n4520), .IN4(n2225), .Q(n4518) );
  OA22X1 U31726 ( .IN1(n2277), .IN2(n19742), .IN3(n2191), .IN4(n19721), .Q(
        n7286) );
  OA22X1 U31727 ( .IN1(n2276), .IN2(n19742), .IN3(n2190), .IN4(n19722), .Q(
        n7282) );
  OA22X1 U31728 ( .IN1(n2275), .IN2(n19738), .IN3(n2189), .IN4(n19721), .Q(
        n7278) );
  OA22X1 U31729 ( .IN1(n2274), .IN2(n19742), .IN3(n2188), .IN4(n19724), .Q(
        n7274) );
  OA22X1 U31730 ( .IN1(n2277), .IN2(n19608), .IN3(n2191), .IN4(n19587), .Q(
        n7566) );
  OA22X1 U31731 ( .IN1(n2276), .IN2(n19606), .IN3(n2190), .IN4(n19588), .Q(
        n7562) );
  OA22X1 U31732 ( .IN1(n2275), .IN2(n19608), .IN3(n2189), .IN4(n19588), .Q(
        n7554) );
  OA22X1 U31733 ( .IN1(n2274), .IN2(n19608), .IN3(n2188), .IN4(n19588), .Q(
        n7550) );
  OA22X1 U31734 ( .IN1(n2277), .IN2(n19476), .IN3(n2191), .IN4(n19452), .Q(
        n7862) );
  OA22X1 U31735 ( .IN1(n2276), .IN2(n19474), .IN3(n2190), .IN4(n19455), .Q(
        n7858) );
  OA22X1 U31736 ( .IN1(n2275), .IN2(n19476), .IN3(n2189), .IN4(n19455), .Q(
        n7850) );
  OA22X1 U31737 ( .IN1(n2274), .IN2(n19473), .IN3(n2188), .IN4(n19455), .Q(
        n7846) );
  OA22X1 U31738 ( .IN1(n2277), .IN2(n19344), .IN3(n2191), .IN4(n19320), .Q(
        n8158) );
  OA22X1 U31739 ( .IN1(n2276), .IN2(n19342), .IN3(n2190), .IN4(n19323), .Q(
        n8154) );
  OA22X1 U31740 ( .IN1(n2275), .IN2(n19344), .IN3(n2189), .IN4(n19323), .Q(
        n8146) );
  OA22X1 U31741 ( .IN1(n2274), .IN2(n19341), .IN3(n2188), .IN4(n19323), .Q(
        n8142) );
  OA22X1 U31742 ( .IN1(n2277), .IN2(n19212), .IN3(n2191), .IN4(n19188), .Q(
        n8454) );
  OA22X1 U31743 ( .IN1(n2276), .IN2(n19210), .IN3(n2190), .IN4(n19191), .Q(
        n8450) );
  OA22X1 U31744 ( .IN1(n2275), .IN2(n19212), .IN3(n2189), .IN4(n19191), .Q(
        n8442) );
  OA22X1 U31745 ( .IN1(n2274), .IN2(n19209), .IN3(n2188), .IN4(n19191), .Q(
        n8438) );
  OA22X1 U31746 ( .IN1(n2277), .IN2(n8539), .IN3(n2191), .IN4(n19056), .Q(
        n8750) );
  OA22X1 U31747 ( .IN1(n2276), .IN2(n19078), .IN3(n2190), .IN4(n19059), .Q(
        n8746) );
  OA22X1 U31748 ( .IN1(n2275), .IN2(n19080), .IN3(n2189), .IN4(n19059), .Q(
        n8738) );
  OA22X1 U31749 ( .IN1(n2274), .IN2(n19081), .IN3(n2188), .IN4(n19059), .Q(
        n8734) );
  OA22X1 U31750 ( .IN1(n2277), .IN2(n20796), .IN3(n2191), .IN4(n20770), .Q(
        n5014) );
  OA22X1 U31751 ( .IN1(n2276), .IN2(n20792), .IN3(n2190), .IN4(n20773), .Q(
        n5010) );
  OA22X1 U31752 ( .IN1(n2275), .IN2(n4803), .IN3(n2189), .IN4(n20773), .Q(
        n5002) );
  OA22X1 U31753 ( .IN1(n2274), .IN2(n20792), .IN3(n2188), .IN4(n20773), .Q(
        n4998) );
  OA22X1 U31754 ( .IN1(n2277), .IN2(n20662), .IN3(n2191), .IN4(n20641), .Q(
        n5310) );
  OA22X1 U31755 ( .IN1(n2276), .IN2(n20660), .IN3(n2190), .IN4(n20642), .Q(
        n5306) );
  OA22X1 U31756 ( .IN1(n2275), .IN2(n20662), .IN3(n2189), .IN4(n20642), .Q(
        n5298) );
  OA22X1 U31757 ( .IN1(n2274), .IN2(n20662), .IN3(n2188), .IN4(n20642), .Q(
        n5294) );
  OA22X1 U31758 ( .IN1(n2277), .IN2(n20530), .IN3(n2191), .IN4(n20509), .Q(
        n5606) );
  OA22X1 U31759 ( .IN1(n2276), .IN2(n20528), .IN3(n2190), .IN4(n20510), .Q(
        n5602) );
  OA22X1 U31760 ( .IN1(n2275), .IN2(n20530), .IN3(n2189), .IN4(n20510), .Q(
        n5594) );
  OA22X1 U31761 ( .IN1(n2274), .IN2(n20530), .IN3(n2188), .IN4(n20510), .Q(
        n5590) );
  OA22X1 U31762 ( .IN1(n2277), .IN2(n20398), .IN3(n2191), .IN4(n20377), .Q(
        n5902) );
  OA22X1 U31763 ( .IN1(n2276), .IN2(n20396), .IN3(n2190), .IN4(n20378), .Q(
        n5898) );
  OA22X1 U31764 ( .IN1(n2275), .IN2(n20398), .IN3(n2189), .IN4(n20378), .Q(
        n5890) );
  OA22X1 U31765 ( .IN1(n2274), .IN2(n20398), .IN3(n2188), .IN4(n20378), .Q(
        n5886) );
  OA22X1 U31766 ( .IN1(n2277), .IN2(n20266), .IN3(n2191), .IN4(n20245), .Q(
        n6198) );
  OA22X1 U31767 ( .IN1(n2276), .IN2(n20264), .IN3(n2190), .IN4(n20246), .Q(
        n6194) );
  OA22X1 U31768 ( .IN1(n2275), .IN2(n20266), .IN3(n2189), .IN4(n20246), .Q(
        n6186) );
  OA22X1 U31769 ( .IN1(n2274), .IN2(n20266), .IN3(n2188), .IN4(n20246), .Q(
        n6182) );
  OA22X1 U31770 ( .IN1(n2277), .IN2(n20134), .IN3(n2191), .IN4(n20110), .Q(
        n6494) );
  OA22X1 U31771 ( .IN1(n2276), .IN2(n20132), .IN3(n2190), .IN4(n20113), .Q(
        n6490) );
  OA22X1 U31772 ( .IN1(n2275), .IN2(n20134), .IN3(n2189), .IN4(n20113), .Q(
        n6482) );
  OA22X1 U31773 ( .IN1(n2274), .IN2(n20135), .IN3(n2188), .IN4(n20113), .Q(
        n6478) );
  OA22X1 U31774 ( .IN1(n2277), .IN2(n20005), .IN3(n2191), .IN4(n19979), .Q(
        n6790) );
  OA22X1 U31775 ( .IN1(n2276), .IN2(n20001), .IN3(n2190), .IN4(n19982), .Q(
        n6786) );
  OA22X1 U31776 ( .IN1(n2275), .IN2(n6579), .IN3(n2189), .IN4(n19982), .Q(
        n6778) );
  OA22X1 U31777 ( .IN1(n2274), .IN2(n20001), .IN3(n2188), .IN4(n19982), .Q(
        n6774) );
  OA22X1 U31778 ( .IN1(n2277), .IN2(n6875), .IN3(n2191), .IN4(n19848), .Q(
        n7086) );
  OA22X1 U31779 ( .IN1(n2276), .IN2(n19870), .IN3(n2190), .IN4(n19851), .Q(
        n7082) );
  OA22X1 U31780 ( .IN1(n2275), .IN2(n19872), .IN3(n2189), .IN4(n19851), .Q(
        n7074) );
  OA22X1 U31781 ( .IN1(n2274), .IN2(n19873), .IN3(n2188), .IN4(n19851), .Q(
        n7070) );
  OA22X1 U31782 ( .IN1(n2277), .IN2(n8835), .IN3(n2191), .IN4(n18924), .Q(
        n9046) );
  OA22X1 U31783 ( .IN1(n2276), .IN2(n18946), .IN3(n2190), .IN4(n18927), .Q(
        n9042) );
  OA22X1 U31784 ( .IN1(n2275), .IN2(n18948), .IN3(n2189), .IN4(n18927), .Q(
        n9034) );
  OA22X1 U31785 ( .IN1(n2274), .IN2(n18949), .IN3(n2188), .IN4(n18927), .Q(
        n9030) );
  OA22X1 U31786 ( .IN1(n18794), .IN2(n2728), .IN3(n18791), .IN4(n2693), .Q(
        n14810) );
  OA22X1 U31787 ( .IN1(n18782), .IN2(n2588), .IN3(n18779), .IN4(n2553), .Q(
        n14811) );
  OA22X1 U31788 ( .IN1(n18770), .IN2(n2378), .IN3(n18767), .IN4(n2343), .Q(
        n14812) );
  OA22X1 U31789 ( .IN1(n18795), .IN2(n2727), .IN3(n14523), .IN4(n2692), .Q(
        n14711) );
  OA22X1 U31790 ( .IN1(n18783), .IN2(n2587), .IN3(n18780), .IN4(n2552), .Q(
        n14712) );
  OA22X1 U31791 ( .IN1(n18771), .IN2(n2377), .IN3(n18768), .IN4(n2342), .Q(
        n14713) );
  OA22X1 U31792 ( .IN1(n18794), .IN2(n2726), .IN3(n18792), .IN4(n2691), .Q(
        n14612) );
  OA22X1 U31793 ( .IN1(n18783), .IN2(n2586), .IN3(n18781), .IN4(n2551), .Q(
        n14613) );
  OA22X1 U31794 ( .IN1(n18772), .IN2(n2376), .IN3(n14533), .IN4(n2341), .Q(
        n14614) );
  OA22X1 U31795 ( .IN1(n18796), .IN2(n2725), .IN3(n18792), .IN4(n2690), .Q(
        n14585) );
  OA22X1 U31796 ( .IN1(n18784), .IN2(n2585), .IN3(n18781), .IN4(n2550), .Q(
        n14586) );
  OA22X1 U31797 ( .IN1(n18770), .IN2(n2375), .IN3(n18768), .IN4(n2340), .Q(
        n14587) );
  OA22X1 U31798 ( .IN1(n18794), .IN2(n2724), .IN3(n18792), .IN4(n2689), .Q(
        n14576) );
  OA22X1 U31799 ( .IN1(n18782), .IN2(n2584), .IN3(n18781), .IN4(n2549), .Q(
        n14577) );
  OA22X1 U31800 ( .IN1(n18771), .IN2(n2374), .IN3(n18768), .IN4(n2339), .Q(
        n14578) );
  OA22X1 U31801 ( .IN1(n18795), .IN2(n2723), .IN3(n18792), .IN4(n2688), .Q(
        n14567) );
  OA22X1 U31802 ( .IN1(n18782), .IN2(n2583), .IN3(n18779), .IN4(n2548), .Q(
        n14568) );
  OA22X1 U31803 ( .IN1(n18772), .IN2(n2373), .IN3(n18768), .IN4(n2338), .Q(
        n14569) );
  OA22X1 U31804 ( .IN1(n18796), .IN2(n2722), .IN3(n18792), .IN4(n2687), .Q(
        n14558) );
  OA22X1 U31805 ( .IN1(n18784), .IN2(n2582), .IN3(n18781), .IN4(n2547), .Q(
        n14559) );
  OA22X1 U31806 ( .IN1(n18772), .IN2(n2372), .IN3(n18768), .IN4(n2337), .Q(
        n14560) );
  OA22X1 U31807 ( .IN1(n18796), .IN2(n2721), .IN3(n18792), .IN4(n2686), .Q(
        n14549) );
  OA22X1 U31808 ( .IN1(n18784), .IN2(n2581), .IN3(n18781), .IN4(n2546), .Q(
        n14550) );
  OA22X1 U31809 ( .IN1(n18772), .IN2(n2371), .IN3(n18768), .IN4(n2336), .Q(
        n14551) );
  OA22X1 U31810 ( .IN1(n18796), .IN2(n2720), .IN3(n18792), .IN4(n2685), .Q(
        n14540) );
  OA22X1 U31811 ( .IN1(n18784), .IN2(n2580), .IN3(n18781), .IN4(n2545), .Q(
        n14541) );
  OA22X1 U31812 ( .IN1(n18772), .IN2(n2370), .IN3(n18768), .IN4(n2335), .Q(
        n14542) );
  OA22X1 U31813 ( .IN1(n18796), .IN2(n2719), .IN3(n18792), .IN4(n2684), .Q(
        n14521) );
  OA22X1 U31814 ( .IN1(n18784), .IN2(n2579), .IN3(n18781), .IN4(n2544), .Q(
        n14526) );
  OA22X1 U31815 ( .IN1(n18772), .IN2(n2369), .IN3(n18768), .IN4(n2334), .Q(
        n14531) );
  OA22X1 U31816 ( .IN1(n18794), .IN2(n2718), .IN3(n18791), .IN4(n2683), .Q(
        n14801) );
  OA22X1 U31817 ( .IN1(n18782), .IN2(n2578), .IN3(n18779), .IN4(n2543), .Q(
        n14802) );
  OA22X1 U31818 ( .IN1(n18770), .IN2(n2368), .IN3(n18767), .IN4(n2333), .Q(
        n14803) );
  OA22X1 U31819 ( .IN1(n18794), .IN2(n2717), .IN3(n18791), .IN4(n2682), .Q(
        n14792) );
  OA22X1 U31820 ( .IN1(n18782), .IN2(n2577), .IN3(n18779), .IN4(n2542), .Q(
        n14793) );
  OA22X1 U31821 ( .IN1(n18770), .IN2(n2367), .IN3(n18767), .IN4(n2332), .Q(
        n14794) );
  OA22X1 U31822 ( .IN1(n18796), .IN2(n2716), .IN3(n18791), .IN4(n2681), .Q(
        n14783) );
  OA22X1 U31823 ( .IN1(n18782), .IN2(n2576), .IN3(n18779), .IN4(n2541), .Q(
        n14784) );
  OA22X1 U31824 ( .IN1(n18770), .IN2(n2366), .IN3(n18767), .IN4(n2331), .Q(
        n14785) );
  OA22X1 U31825 ( .IN1(n18796), .IN2(n2715), .IN3(n18791), .IN4(n2680), .Q(
        n14774) );
  OA22X1 U31826 ( .IN1(n18784), .IN2(n2575), .IN3(n18780), .IN4(n2540), .Q(
        n14775) );
  OA22X1 U31827 ( .IN1(n18770), .IN2(n2365), .IN3(n14533), .IN4(n2330), .Q(
        n14776) );
  OA22X1 U31828 ( .IN1(n18796), .IN2(n2714), .IN3(n18791), .IN4(n2679), .Q(
        n14765) );
  OA22X1 U31829 ( .IN1(n18782), .IN2(n2574), .IN3(n18780), .IN4(n2539), .Q(
        n14766) );
  OA22X1 U31830 ( .IN1(n18771), .IN2(n2364), .IN3(n14533), .IN4(n2329), .Q(
        n14767) );
  OA22X1 U31831 ( .IN1(n18795), .IN2(n2713), .IN3(n14523), .IN4(n2678), .Q(
        n14756) );
  OA22X1 U31832 ( .IN1(n18783), .IN2(n2573), .IN3(n18780), .IN4(n2538), .Q(
        n14757) );
  OA22X1 U31833 ( .IN1(n18772), .IN2(n2363), .IN3(n14533), .IN4(n2328), .Q(
        n14758) );
  OA22X1 U31834 ( .IN1(n18796), .IN2(n2712), .IN3(n14523), .IN4(n2677), .Q(
        n14747) );
  OA22X1 U31835 ( .IN1(n18784), .IN2(n2572), .IN3(n18780), .IN4(n2537), .Q(
        n14748) );
  OA22X1 U31836 ( .IN1(n18772), .IN2(n2362), .IN3(n14533), .IN4(n2327), .Q(
        n14749) );
  OA22X1 U31837 ( .IN1(n18796), .IN2(n2711), .IN3(n14523), .IN4(n2676), .Q(
        n14738) );
  OA22X1 U31838 ( .IN1(n18784), .IN2(n2571), .IN3(n18781), .IN4(n2536), .Q(
        n14739) );
  OA22X1 U31839 ( .IN1(n18771), .IN2(n2361), .IN3(n14533), .IN4(n2326), .Q(
        n14740) );
  OA22X1 U31840 ( .IN1(n18795), .IN2(n2710), .IN3(n14523), .IN4(n2675), .Q(
        n14729) );
  OA22X1 U31841 ( .IN1(n18782), .IN2(n2570), .IN3(n18779), .IN4(n2535), .Q(
        n14730) );
  OA22X1 U31842 ( .IN1(n18771), .IN2(n2360), .IN3(n14533), .IN4(n2325), .Q(
        n14731) );
  OA22X1 U31843 ( .IN1(n18795), .IN2(n2709), .IN3(n14523), .IN4(n2674), .Q(
        n14720) );
  OA22X1 U31844 ( .IN1(n18784), .IN2(n2569), .IN3(n18780), .IN4(n2534), .Q(
        n14721) );
  OA22X1 U31845 ( .IN1(n18771), .IN2(n2359), .IN3(n14533), .IN4(n2324), .Q(
        n14722) );
  OA22X1 U31846 ( .IN1(n18794), .IN2(n2708), .IN3(n14523), .IN4(n2673), .Q(
        n14702) );
  OA22X1 U31847 ( .IN1(n18784), .IN2(n2568), .IN3(n18779), .IN4(n2533), .Q(
        n14703) );
  OA22X1 U31848 ( .IN1(n18770), .IN2(n2358), .IN3(n18767), .IN4(n2323), .Q(
        n14704) );
  OA22X1 U31849 ( .IN1(n18794), .IN2(n2707), .IN3(n18791), .IN4(n2672), .Q(
        n14693) );
  OA22X1 U31850 ( .IN1(n18784), .IN2(n2567), .IN3(n18780), .IN4(n2532), .Q(
        n14694) );
  OA22X1 U31851 ( .IN1(n18770), .IN2(n2357), .IN3(n18768), .IN4(n2322), .Q(
        n14695) );
  OA22X1 U31852 ( .IN1(n18794), .IN2(n2706), .IN3(n18791), .IN4(n2671), .Q(
        n14684) );
  OA22X1 U31853 ( .IN1(n18782), .IN2(n2566), .IN3(n18781), .IN4(n2531), .Q(
        n14685) );
  OA22X1 U31854 ( .IN1(n18771), .IN2(n2356), .IN3(n18767), .IN4(n2321), .Q(
        n14686) );
  OA22X1 U31855 ( .IN1(n18794), .IN2(n2705), .IN3(n14523), .IN4(n2670), .Q(
        n14675) );
  OA22X1 U31856 ( .IN1(n18783), .IN2(n2565), .IN3(n18779), .IN4(n2530), .Q(
        n14676) );
  OA22X1 U31857 ( .IN1(n18771), .IN2(n2355), .IN3(n14533), .IN4(n2320), .Q(
        n14677) );
  OA22X1 U31858 ( .IN1(n18795), .IN2(n2704), .IN3(n18791), .IN4(n2669), .Q(
        n14666) );
  OA22X1 U31859 ( .IN1(n18783), .IN2(n2564), .IN3(n18779), .IN4(n2529), .Q(
        n14667) );
  OA22X1 U31860 ( .IN1(n18771), .IN2(n2354), .IN3(n18767), .IN4(n2319), .Q(
        n14668) );
  OA22X1 U31861 ( .IN1(n18795), .IN2(n2703), .IN3(n18791), .IN4(n2668), .Q(
        n14657) );
  OA22X1 U31862 ( .IN1(n18783), .IN2(n2563), .IN3(n18780), .IN4(n2528), .Q(
        n14658) );
  OA22X1 U31863 ( .IN1(n18772), .IN2(n2353), .IN3(n18767), .IN4(n2318), .Q(
        n14659) );
  OA22X1 U31864 ( .IN1(n18795), .IN2(n2702), .IN3(n14523), .IN4(n2667), .Q(
        n14648) );
  OA22X1 U31865 ( .IN1(n18783), .IN2(n2562), .IN3(n18781), .IN4(n2527), .Q(
        n14649) );
  OA22X1 U31866 ( .IN1(n18771), .IN2(n2352), .IN3(n14533), .IN4(n2317), .Q(
        n14650) );
  OA22X1 U31867 ( .IN1(n18795), .IN2(n2701), .IN3(n14523), .IN4(n2666), .Q(
        n14639) );
  OA22X1 U31868 ( .IN1(n18783), .IN2(n2561), .IN3(n18779), .IN4(n2526), .Q(
        n14640) );
  OA22X1 U31869 ( .IN1(n18770), .IN2(n2351), .IN3(n18767), .IN4(n2316), .Q(
        n14641) );
  OA22X1 U31870 ( .IN1(n18794), .IN2(n2700), .IN3(n14523), .IN4(n2665), .Q(
        n14630) );
  OA22X1 U31871 ( .IN1(n18783), .IN2(n2560), .IN3(n18779), .IN4(n2525), .Q(
        n14631) );
  OA22X1 U31872 ( .IN1(n18772), .IN2(n2350), .IN3(n14533), .IN4(n2315), .Q(
        n14632) );
  OA22X1 U31873 ( .IN1(n18794), .IN2(n2699), .IN3(n18792), .IN4(n2664), .Q(
        n14621) );
  OA22X1 U31874 ( .IN1(n18783), .IN2(n2559), .IN3(n18780), .IN4(n2524), .Q(
        n14622) );
  OA22X1 U31875 ( .IN1(n18770), .IN2(n2349), .IN3(n14533), .IN4(n2314), .Q(
        n14623) );
  OA22X1 U31876 ( .IN1(n18795), .IN2(n2698), .IN3(n18792), .IN4(n2663), .Q(
        n14603) );
  OA22X1 U31877 ( .IN1(n18783), .IN2(n2558), .IN3(n18781), .IN4(n2523), .Q(
        n14604) );
  OA22X1 U31878 ( .IN1(n18772), .IN2(n2348), .IN3(n14533), .IN4(n2313), .Q(
        n14605) );
  OA22X1 U31879 ( .IN1(n18795), .IN2(n2697), .IN3(n14523), .IN4(n2662), .Q(
        n14594) );
  OA22X1 U31880 ( .IN1(n18782), .IN2(n2557), .IN3(n18780), .IN4(n2522), .Q(
        n14595) );
  OA22X1 U31881 ( .IN1(n18770), .IN2(n2347), .IN3(n14533), .IN4(n2312), .Q(
        n14596) );
  OA22X1 U31882 ( .IN1(n18746), .IN2(n2728), .IN3(n18743), .IN4(n2693), .Q(
        n15161) );
  OA22X1 U31883 ( .IN1(n18734), .IN2(n2588), .IN3(n14910), .IN4(n2553), .Q(
        n15162) );
  OA22X1 U31884 ( .IN1(n18724), .IN2(n2378), .IN3(n18719), .IN4(n2343), .Q(
        n15163) );
  OA22X1 U31885 ( .IN1(n18748), .IN2(n2727), .IN3(n14905), .IN4(n2692), .Q(
        n15073) );
  OA22X1 U31886 ( .IN1(n18736), .IN2(n2587), .IN3(n18732), .IN4(n2552), .Q(
        n15074) );
  OA22X1 U31887 ( .IN1(n18722), .IN2(n2377), .IN3(n14915), .IN4(n2342), .Q(
        n15075) );
  OA22X1 U31888 ( .IN1(n18746), .IN2(n2726), .IN3(n18744), .IN4(n2691), .Q(
        n14985) );
  OA22X1 U31889 ( .IN1(n18734), .IN2(n2586), .IN3(n18732), .IN4(n2551), .Q(
        n14986) );
  OA22X1 U31890 ( .IN1(n18724), .IN2(n2376), .IN3(n18720), .IN4(n2341), .Q(
        n14987) );
  OA22X1 U31891 ( .IN1(n18747), .IN2(n2725), .IN3(n18743), .IN4(n2690), .Q(
        n14961) );
  OA22X1 U31892 ( .IN1(n18736), .IN2(n2585), .IN3(n18732), .IN4(n2550), .Q(
        n14962) );
  OA22X1 U31893 ( .IN1(n18723), .IN2(n2375), .IN3(n14915), .IN4(n2340), .Q(
        n14963) );
  OA22X1 U31894 ( .IN1(n18748), .IN2(n2724), .IN3(n18744), .IN4(n2689), .Q(
        n14953) );
  OA22X1 U31895 ( .IN1(n18734), .IN2(n2584), .IN3(n18731), .IN4(n2549), .Q(
        n14954) );
  OA22X1 U31896 ( .IN1(n18722), .IN2(n2374), .IN3(n18720), .IN4(n2339), .Q(
        n14955) );
  OA22X1 U31897 ( .IN1(n18748), .IN2(n2723), .IN3(n14905), .IN4(n2688), .Q(
        n14945) );
  OA22X1 U31898 ( .IN1(n18735), .IN2(n2583), .IN3(n14910), .IN4(n2548), .Q(
        n14946) );
  OA22X1 U31899 ( .IN1(n18722), .IN2(n2373), .IN3(n14915), .IN4(n2338), .Q(
        n14947) );
  OA22X1 U31900 ( .IN1(n18746), .IN2(n2722), .IN3(n18744), .IN4(n2687), .Q(
        n14937) );
  OA22X1 U31901 ( .IN1(n18736), .IN2(n2582), .IN3(n18732), .IN4(n2547), .Q(
        n14938) );
  OA22X1 U31902 ( .IN1(n18724), .IN2(n2372), .IN3(n18720), .IN4(n2337), .Q(
        n14939) );
  OA22X1 U31903 ( .IN1(n18748), .IN2(n2721), .IN3(n18744), .IN4(n2686), .Q(
        n14929) );
  OA22X1 U31904 ( .IN1(n18736), .IN2(n2581), .IN3(n18732), .IN4(n2546), .Q(
        n14930) );
  OA22X1 U31905 ( .IN1(n18724), .IN2(n2371), .IN3(n18720), .IN4(n2336), .Q(
        n14931) );
  OA22X1 U31906 ( .IN1(n18746), .IN2(n2720), .IN3(n18744), .IN4(n2685), .Q(
        n14921) );
  OA22X1 U31907 ( .IN1(n18736), .IN2(n2580), .IN3(n18732), .IN4(n2545), .Q(
        n14922) );
  OA22X1 U31908 ( .IN1(n18724), .IN2(n2370), .IN3(n18720), .IN4(n2335), .Q(
        n14923) );
  OA22X1 U31909 ( .IN1(n18746), .IN2(n2719), .IN3(n18744), .IN4(n2684), .Q(
        n14903) );
  OA22X1 U31910 ( .IN1(n18736), .IN2(n2579), .IN3(n18732), .IN4(n2544), .Q(
        n14908) );
  OA22X1 U31911 ( .IN1(n18724), .IN2(n2369), .IN3(n18720), .IN4(n2334), .Q(
        n14913) );
  OA22X1 U31912 ( .IN1(n18746), .IN2(n2718), .IN3(n18743), .IN4(n2683), .Q(
        n15153) );
  OA22X1 U31913 ( .IN1(n18735), .IN2(n2578), .IN3(n14910), .IN4(n2543), .Q(
        n15154) );
  OA22X1 U31914 ( .IN1(n18722), .IN2(n2368), .IN3(n18719), .IN4(n2333), .Q(
        n15155) );
  OA22X1 U31915 ( .IN1(n18746), .IN2(n2717), .IN3(n18743), .IN4(n2682), .Q(
        n15145) );
  OA22X1 U31916 ( .IN1(n18734), .IN2(n2577), .IN3(n14910), .IN4(n2542), .Q(
        n15146) );
  OA22X1 U31917 ( .IN1(n18723), .IN2(n2367), .IN3(n18719), .IN4(n2332), .Q(
        n15147) );
  OA22X1 U31918 ( .IN1(n18746), .IN2(n2716), .IN3(n18743), .IN4(n2681), .Q(
        n15137) );
  OA22X1 U31919 ( .IN1(n18735), .IN2(n2576), .IN3(n14910), .IN4(n2541), .Q(
        n15138) );
  OA22X1 U31920 ( .IN1(n18724), .IN2(n2366), .IN3(n18719), .IN4(n2331), .Q(
        n15139) );
  OA22X1 U31921 ( .IN1(n18747), .IN2(n2715), .IN3(n14905), .IN4(n2680), .Q(
        n15129) );
  OA22X1 U31922 ( .IN1(n18734), .IN2(n2575), .IN3(n18731), .IN4(n2540), .Q(
        n15130) );
  OA22X1 U31923 ( .IN1(n18722), .IN2(n2365), .IN3(n14915), .IN4(n2330), .Q(
        n15131) );
  OA22X1 U31924 ( .IN1(n18747), .IN2(n2714), .IN3(n14905), .IN4(n2679), .Q(
        n15121) );
  OA22X1 U31925 ( .IN1(n18734), .IN2(n2574), .IN3(n18731), .IN4(n2539), .Q(
        n15122) );
  OA22X1 U31926 ( .IN1(n18722), .IN2(n2364), .IN3(n14915), .IN4(n2329), .Q(
        n15123) );
  OA22X1 U31927 ( .IN1(n18747), .IN2(n2713), .IN3(n14905), .IN4(n2678), .Q(
        n15113) );
  OA22X1 U31928 ( .IN1(n18734), .IN2(n2573), .IN3(n18731), .IN4(n2538), .Q(
        n15114) );
  OA22X1 U31929 ( .IN1(n18722), .IN2(n2363), .IN3(n14915), .IN4(n2328), .Q(
        n15115) );
  OA22X1 U31930 ( .IN1(n18747), .IN2(n2712), .IN3(n14905), .IN4(n2677), .Q(
        n15105) );
  OA22X1 U31931 ( .IN1(n18734), .IN2(n2572), .IN3(n18731), .IN4(n2537), .Q(
        n15106) );
  OA22X1 U31932 ( .IN1(n18722), .IN2(n2362), .IN3(n14915), .IN4(n2327), .Q(
        n15107) );
  OA22X1 U31933 ( .IN1(n18748), .IN2(n2711), .IN3(n14905), .IN4(n2676), .Q(
        n15097) );
  OA22X1 U31934 ( .IN1(n18735), .IN2(n2571), .IN3(n18731), .IN4(n2536), .Q(
        n15098) );
  OA22X1 U31935 ( .IN1(n18723), .IN2(n2361), .IN3(n18719), .IN4(n2326), .Q(
        n15099) );
  OA22X1 U31936 ( .IN1(n18748), .IN2(n2710), .IN3(n14905), .IN4(n2675), .Q(
        n15089) );
  OA22X1 U31937 ( .IN1(n18735), .IN2(n2570), .IN3(n18732), .IN4(n2535), .Q(
        n15090) );
  OA22X1 U31938 ( .IN1(n18722), .IN2(n2360), .IN3(n14915), .IN4(n2325), .Q(
        n15091) );
  OA22X1 U31939 ( .IN1(n18748), .IN2(n2709), .IN3(n14905), .IN4(n2674), .Q(
        n15081) );
  OA22X1 U31940 ( .IN1(n18734), .IN2(n2569), .IN3(n18732), .IN4(n2534), .Q(
        n15082) );
  OA22X1 U31941 ( .IN1(n18723), .IN2(n2359), .IN3(n14915), .IN4(n2324), .Q(
        n15083) );
  OA22X1 U31942 ( .IN1(n18746), .IN2(n2708), .IN3(n18743), .IN4(n2673), .Q(
        n15065) );
  OA22X1 U31943 ( .IN1(n18735), .IN2(n2568), .IN3(n14910), .IN4(n2533), .Q(
        n15066) );
  OA22X1 U31944 ( .IN1(n18723), .IN2(n2358), .IN3(n14915), .IN4(n2323), .Q(
        n15067) );
  OA22X1 U31945 ( .IN1(n18747), .IN2(n2707), .IN3(n14905), .IN4(n2672), .Q(
        n15057) );
  OA22X1 U31946 ( .IN1(n18735), .IN2(n2567), .IN3(n14910), .IN4(n2532), .Q(
        n15058) );
  OA22X1 U31947 ( .IN1(n18723), .IN2(n2357), .IN3(n18720), .IN4(n2322), .Q(
        n15059) );
  OA22X1 U31948 ( .IN1(n18747), .IN2(n2706), .IN3(n18743), .IN4(n2671), .Q(
        n15049) );
  OA22X1 U31949 ( .IN1(n18735), .IN2(n2566), .IN3(n14910), .IN4(n2531), .Q(
        n15050) );
  OA22X1 U31950 ( .IN1(n18722), .IN2(n2356), .IN3(n18719), .IN4(n2321), .Q(
        n15051) );
  OA22X1 U31951 ( .IN1(n18748), .IN2(n2705), .IN3(n18743), .IN4(n2670), .Q(
        n15041) );
  OA22X1 U31952 ( .IN1(n18735), .IN2(n2565), .IN3(n14910), .IN4(n2530), .Q(
        n15042) );
  OA22X1 U31953 ( .IN1(n18722), .IN2(n2355), .IN3(n14915), .IN4(n2320), .Q(
        n15043) );
  OA22X1 U31954 ( .IN1(n18748), .IN2(n2704), .IN3(n18743), .IN4(n2669), .Q(
        n15033) );
  OA22X1 U31955 ( .IN1(n18735), .IN2(n2564), .IN3(n18731), .IN4(n2529), .Q(
        n15034) );
  OA22X1 U31956 ( .IN1(n18723), .IN2(n2354), .IN3(n18719), .IN4(n2319), .Q(
        n15035) );
  OA22X1 U31957 ( .IN1(n18746), .IN2(n2703), .IN3(n18743), .IN4(n2668), .Q(
        n15025) );
  OA22X1 U31958 ( .IN1(n18736), .IN2(n2563), .IN3(n18731), .IN4(n2528), .Q(
        n15026) );
  OA22X1 U31959 ( .IN1(n18723), .IN2(n2353), .IN3(n18719), .IN4(n2318), .Q(
        n15027) );
  OA22X1 U31960 ( .IN1(n18747), .IN2(n2702), .IN3(n14905), .IN4(n2667), .Q(
        n15017) );
  OA22X1 U31961 ( .IN1(n18735), .IN2(n2562), .IN3(n14910), .IN4(n2527), .Q(
        n15018) );
  OA22X1 U31962 ( .IN1(n18723), .IN2(n2352), .IN3(n18720), .IN4(n2317), .Q(
        n15019) );
  OA22X1 U31963 ( .IN1(n18747), .IN2(n2701), .IN3(n18744), .IN4(n2666), .Q(
        n15009) );
  OA22X1 U31964 ( .IN1(n18734), .IN2(n2561), .IN3(n14910), .IN4(n2526), .Q(
        n15010) );
  OA22X1 U31965 ( .IN1(n18723), .IN2(n2351), .IN3(n18719), .IN4(n2316), .Q(
        n15011) );
  OA22X1 U31966 ( .IN1(n18747), .IN2(n2700), .IN3(n18744), .IN4(n2665), .Q(
        n15001) );
  OA22X1 U31967 ( .IN1(n18736), .IN2(n2560), .IN3(n14910), .IN4(n2525), .Q(
        n15002) );
  OA22X1 U31968 ( .IN1(n18724), .IN2(n2350), .IN3(n14915), .IN4(n2315), .Q(
        n15003) );
  OA22X1 U31969 ( .IN1(n18748), .IN2(n2699), .IN3(n14905), .IN4(n2664), .Q(
        n14993) );
  OA22X1 U31970 ( .IN1(n18734), .IN2(n2559), .IN3(n18731), .IN4(n2524), .Q(
        n14994) );
  OA22X1 U31971 ( .IN1(n18723), .IN2(n2349), .IN3(n14915), .IN4(n2314), .Q(
        n14995) );
  OA22X1 U31972 ( .IN1(n18746), .IN2(n2698), .IN3(n18744), .IN4(n2663), .Q(
        n14977) );
  OA22X1 U31973 ( .IN1(n18736), .IN2(n2558), .IN3(n18732), .IN4(n2523), .Q(
        n14978) );
  OA22X1 U31974 ( .IN1(n18724), .IN2(n2348), .IN3(n14915), .IN4(n2313), .Q(
        n14979) );
  OA22X1 U31975 ( .IN1(n18747), .IN2(n2697), .IN3(n18744), .IN4(n2662), .Q(
        n14969) );
  OA22X1 U31976 ( .IN1(n18736), .IN2(n2557), .IN3(n18731), .IN4(n2522), .Q(
        n14970) );
  OA22X1 U31977 ( .IN1(n18724), .IN2(n2347), .IN3(n18720), .IN4(n2312), .Q(
        n14971) );
  OA22X1 U31978 ( .IN1(n18698), .IN2(n2728), .IN3(n18695), .IN4(n2693), .Q(
        n15466) );
  OA22X1 U31979 ( .IN1(n18687), .IN2(n2588), .IN3(n18683), .IN4(n2553), .Q(
        n15467) );
  OA22X1 U31980 ( .IN1(n18674), .IN2(n2378), .IN3(n18671), .IN4(n2343), .Q(
        n15468) );
  OA22X1 U31981 ( .IN1(n18700), .IN2(n2727), .IN3(n15210), .IN4(n2692), .Q(
        n15378) );
  OA22X1 U31982 ( .IN1(n18686), .IN2(n2587), .IN3(n18684), .IN4(n2552), .Q(
        n15379) );
  OA22X1 U31983 ( .IN1(n18675), .IN2(n2377), .IN3(n18672), .IN4(n2342), .Q(
        n15380) );
  OA22X1 U31984 ( .IN1(n18699), .IN2(n2726), .IN3(n18696), .IN4(n2691), .Q(
        n15290) );
  OA22X1 U31985 ( .IN1(n18687), .IN2(n2586), .IN3(n18685), .IN4(n2551), .Q(
        n15291) );
  OA22X1 U31986 ( .IN1(n18676), .IN2(n2376), .IN3(n15220), .IN4(n2341), .Q(
        n15292) );
  OA22X1 U31987 ( .IN1(n18698), .IN2(n2725), .IN3(n18696), .IN4(n2690), .Q(
        n15266) );
  OA22X1 U31988 ( .IN1(n18686), .IN2(n2585), .IN3(n18685), .IN4(n2550), .Q(
        n15267) );
  OA22X1 U31989 ( .IN1(n18674), .IN2(n2375), .IN3(n18672), .IN4(n2340), .Q(
        n15268) );
  OA22X1 U31990 ( .IN1(n18699), .IN2(n2724), .IN3(n18696), .IN4(n2689), .Q(
        n15258) );
  OA22X1 U31991 ( .IN1(n18688), .IN2(n2584), .IN3(n18685), .IN4(n2549), .Q(
        n15259) );
  OA22X1 U31992 ( .IN1(n18675), .IN2(n2374), .IN3(n18672), .IN4(n2339), .Q(
        n15260) );
  OA22X1 U31993 ( .IN1(n18700), .IN2(n2723), .IN3(n18696), .IN4(n2688), .Q(
        n15250) );
  OA22X1 U31994 ( .IN1(n18687), .IN2(n2583), .IN3(n18683), .IN4(n2548), .Q(
        n15251) );
  OA22X1 U31995 ( .IN1(n18676), .IN2(n2373), .IN3(n18672), .IN4(n2338), .Q(
        n15252) );
  OA22X1 U31996 ( .IN1(n18700), .IN2(n2722), .IN3(n18696), .IN4(n2687), .Q(
        n15242) );
  OA22X1 U31997 ( .IN1(n18688), .IN2(n2582), .IN3(n18685), .IN4(n2547), .Q(
        n15243) );
  OA22X1 U31998 ( .IN1(n18676), .IN2(n2372), .IN3(n18672), .IN4(n2337), .Q(
        n15244) );
  OA22X1 U31999 ( .IN1(n18700), .IN2(n2721), .IN3(n18696), .IN4(n2686), .Q(
        n15234) );
  OA22X1 U32000 ( .IN1(n18688), .IN2(n2581), .IN3(n18685), .IN4(n2546), .Q(
        n15235) );
  OA22X1 U32001 ( .IN1(n18676), .IN2(n2371), .IN3(n18672), .IN4(n2336), .Q(
        n15236) );
  OA22X1 U32002 ( .IN1(n18700), .IN2(n2720), .IN3(n18696), .IN4(n2685), .Q(
        n15226) );
  OA22X1 U32003 ( .IN1(n18688), .IN2(n2580), .IN3(n18685), .IN4(n2545), .Q(
        n15227) );
  OA22X1 U32004 ( .IN1(n18676), .IN2(n2370), .IN3(n18672), .IN4(n2335), .Q(
        n15228) );
  OA22X1 U32005 ( .IN1(n18700), .IN2(n2719), .IN3(n18696), .IN4(n2684), .Q(
        n15208) );
  OA22X1 U32006 ( .IN1(n18688), .IN2(n2579), .IN3(n18685), .IN4(n2544), .Q(
        n15213) );
  OA22X1 U32007 ( .IN1(n18676), .IN2(n2369), .IN3(n18672), .IN4(n2334), .Q(
        n15218) );
  OA22X1 U32008 ( .IN1(n18698), .IN2(n2718), .IN3(n18695), .IN4(n2683), .Q(
        n15458) );
  OA22X1 U32009 ( .IN1(n18688), .IN2(n2578), .IN3(n18683), .IN4(n2543), .Q(
        n15459) );
  OA22X1 U32010 ( .IN1(n18674), .IN2(n2368), .IN3(n18671), .IN4(n2333), .Q(
        n15460) );
  OA22X1 U32011 ( .IN1(n18698), .IN2(n2717), .IN3(n18695), .IN4(n2682), .Q(
        n15450) );
  OA22X1 U32012 ( .IN1(n18686), .IN2(n2577), .IN3(n18683), .IN4(n2542), .Q(
        n15451) );
  OA22X1 U32013 ( .IN1(n18674), .IN2(n2367), .IN3(n18671), .IN4(n2332), .Q(
        n15452) );
  OA22X1 U32014 ( .IN1(n18698), .IN2(n2716), .IN3(n18695), .IN4(n2681), .Q(
        n15442) );
  OA22X1 U32015 ( .IN1(n18686), .IN2(n2576), .IN3(n18683), .IN4(n2541), .Q(
        n15443) );
  OA22X1 U32016 ( .IN1(n18674), .IN2(n2366), .IN3(n18671), .IN4(n2331), .Q(
        n15444) );
  OA22X1 U32017 ( .IN1(n18698), .IN2(n2715), .IN3(n15210), .IN4(n2680), .Q(
        n15434) );
  OA22X1 U32018 ( .IN1(n18686), .IN2(n2575), .IN3(n18684), .IN4(n2540), .Q(
        n15435) );
  OA22X1 U32019 ( .IN1(n18674), .IN2(n2365), .IN3(n15220), .IN4(n2330), .Q(
        n15436) );
  OA22X1 U32020 ( .IN1(n18698), .IN2(n2714), .IN3(n15210), .IN4(n2679), .Q(
        n15426) );
  OA22X1 U32021 ( .IN1(n18688), .IN2(n2574), .IN3(n18684), .IN4(n2539), .Q(
        n15427) );
  OA22X1 U32022 ( .IN1(n18675), .IN2(n2364), .IN3(n15220), .IN4(n2329), .Q(
        n15428) );
  OA22X1 U32023 ( .IN1(n18700), .IN2(n2713), .IN3(n15210), .IN4(n2678), .Q(
        n15418) );
  OA22X1 U32024 ( .IN1(n18688), .IN2(n2573), .IN3(n18684), .IN4(n2538), .Q(
        n15419) );
  OA22X1 U32025 ( .IN1(n18676), .IN2(n2363), .IN3(n15220), .IN4(n2328), .Q(
        n15420) );
  OA22X1 U32026 ( .IN1(n18698), .IN2(n2712), .IN3(n15210), .IN4(n2677), .Q(
        n15410) );
  OA22X1 U32027 ( .IN1(n18688), .IN2(n2572), .IN3(n18684), .IN4(n2537), .Q(
        n15411) );
  OA22X1 U32028 ( .IN1(n18676), .IN2(n2362), .IN3(n15220), .IN4(n2327), .Q(
        n15412) );
  OA22X1 U32029 ( .IN1(n18698), .IN2(n2711), .IN3(n15210), .IN4(n2676), .Q(
        n15402) );
  OA22X1 U32030 ( .IN1(n18687), .IN2(n2571), .IN3(n18685), .IN4(n2536), .Q(
        n15403) );
  OA22X1 U32031 ( .IN1(n18675), .IN2(n2361), .IN3(n15220), .IN4(n2326), .Q(
        n15404) );
  OA22X1 U32032 ( .IN1(n18700), .IN2(n2710), .IN3(n15210), .IN4(n2675), .Q(
        n15394) );
  OA22X1 U32033 ( .IN1(n18688), .IN2(n2570), .IN3(n18683), .IN4(n2535), .Q(
        n15395) );
  OA22X1 U32034 ( .IN1(n18675), .IN2(n2360), .IN3(n15220), .IN4(n2325), .Q(
        n15396) );
  OA22X1 U32035 ( .IN1(n18698), .IN2(n2709), .IN3(n15210), .IN4(n2674), .Q(
        n15386) );
  OA22X1 U32036 ( .IN1(n18686), .IN2(n2569), .IN3(n18684), .IN4(n2534), .Q(
        n15387) );
  OA22X1 U32037 ( .IN1(n18675), .IN2(n2359), .IN3(n15220), .IN4(n2324), .Q(
        n15388) );
  OA22X1 U32038 ( .IN1(n18699), .IN2(n2708), .IN3(n18695), .IN4(n2673), .Q(
        n15370) );
  OA22X1 U32039 ( .IN1(n18686), .IN2(n2568), .IN3(n18683), .IN4(n2533), .Q(
        n15371) );
  OA22X1 U32040 ( .IN1(n18674), .IN2(n2358), .IN3(n18671), .IN4(n2323), .Q(
        n15372) );
  OA22X1 U32041 ( .IN1(n18699), .IN2(n2707), .IN3(n15210), .IN4(n2672), .Q(
        n15362) );
  OA22X1 U32042 ( .IN1(n18686), .IN2(n2567), .IN3(n18684), .IN4(n2532), .Q(
        n15363) );
  OA22X1 U32043 ( .IN1(n18674), .IN2(n2357), .IN3(n18672), .IN4(n2322), .Q(
        n15364) );
  OA22X1 U32044 ( .IN1(n18699), .IN2(n2706), .IN3(n18695), .IN4(n2671), .Q(
        n15354) );
  OA22X1 U32045 ( .IN1(n18686), .IN2(n2566), .IN3(n18685), .IN4(n2531), .Q(
        n15355) );
  OA22X1 U32046 ( .IN1(n18675), .IN2(n2356), .IN3(n18671), .IN4(n2321), .Q(
        n15356) );
  OA22X1 U32047 ( .IN1(n18699), .IN2(n2705), .IN3(n18695), .IN4(n2670), .Q(
        n15346) );
  OA22X1 U32048 ( .IN1(n18686), .IN2(n2565), .IN3(n18683), .IN4(n2530), .Q(
        n15347) );
  OA22X1 U32049 ( .IN1(n18675), .IN2(n2355), .IN3(n15220), .IN4(n2320), .Q(
        n15348) );
  OA22X1 U32050 ( .IN1(n18699), .IN2(n2704), .IN3(n18695), .IN4(n2669), .Q(
        n15338) );
  OA22X1 U32051 ( .IN1(n18687), .IN2(n2564), .IN3(n18683), .IN4(n2529), .Q(
        n15339) );
  OA22X1 U32052 ( .IN1(n18675), .IN2(n2354), .IN3(n18671), .IN4(n2319), .Q(
        n15340) );
  OA22X1 U32053 ( .IN1(n18700), .IN2(n2703), .IN3(n18695), .IN4(n2668), .Q(
        n15330) );
  OA22X1 U32054 ( .IN1(n18687), .IN2(n2563), .IN3(n18684), .IN4(n2528), .Q(
        n15331) );
  OA22X1 U32055 ( .IN1(n18676), .IN2(n2353), .IN3(n18671), .IN4(n2318), .Q(
        n15332) );
  OA22X1 U32056 ( .IN1(n18699), .IN2(n2702), .IN3(n15210), .IN4(n2667), .Q(
        n15322) );
  OA22X1 U32057 ( .IN1(n18687), .IN2(n2562), .IN3(n18685), .IN4(n2527), .Q(
        n15323) );
  OA22X1 U32058 ( .IN1(n18675), .IN2(n2352), .IN3(n15220), .IN4(n2317), .Q(
        n15324) );
  OA22X1 U32059 ( .IN1(n18700), .IN2(n2701), .IN3(n18695), .IN4(n2666), .Q(
        n15314) );
  OA22X1 U32060 ( .IN1(n18687), .IN2(n2561), .IN3(n18683), .IN4(n2526), .Q(
        n15315) );
  OA22X1 U32061 ( .IN1(n18674), .IN2(n2351), .IN3(n18671), .IN4(n2316), .Q(
        n15316) );
  OA22X1 U32062 ( .IN1(n18699), .IN2(n2700), .IN3(n18696), .IN4(n2665), .Q(
        n15306) );
  OA22X1 U32063 ( .IN1(n18687), .IN2(n2560), .IN3(n18683), .IN4(n2525), .Q(
        n15307) );
  OA22X1 U32064 ( .IN1(n18676), .IN2(n2350), .IN3(n15220), .IN4(n2315), .Q(
        n15308) );
  OA22X1 U32065 ( .IN1(n18699), .IN2(n2699), .IN3(n15210), .IN4(n2664), .Q(
        n15298) );
  OA22X1 U32066 ( .IN1(n18687), .IN2(n2559), .IN3(n18684), .IN4(n2524), .Q(
        n15299) );
  OA22X1 U32067 ( .IN1(n18674), .IN2(n2349), .IN3(n15220), .IN4(n2314), .Q(
        n15300) );
  OA22X1 U32068 ( .IN1(n18700), .IN2(n2698), .IN3(n18696), .IN4(n2663), .Q(
        n15282) );
  OA22X1 U32069 ( .IN1(n18687), .IN2(n2558), .IN3(n18685), .IN4(n2523), .Q(
        n15283) );
  OA22X1 U32070 ( .IN1(n18676), .IN2(n2348), .IN3(n15220), .IN4(n2313), .Q(
        n15284) );
  OA22X1 U32071 ( .IN1(n18699), .IN2(n2697), .IN3(n15210), .IN4(n2662), .Q(
        n15274) );
  OA22X1 U32072 ( .IN1(n18686), .IN2(n2557), .IN3(n18684), .IN4(n2522), .Q(
        n15275) );
  OA22X1 U32073 ( .IN1(n18674), .IN2(n2347), .IN3(n15220), .IN4(n2312), .Q(
        n15276) );
  OA22X1 U32074 ( .IN1(n18650), .IN2(n2728), .IN3(n18647), .IN4(n2693), .Q(
        n15771) );
  OA22X1 U32075 ( .IN1(n18638), .IN2(n2588), .IN3(n15520), .IN4(n2553), .Q(
        n15772) );
  OA22X1 U32076 ( .IN1(n18628), .IN2(n2378), .IN3(n18623), .IN4(n2343), .Q(
        n15773) );
  OA22X1 U32077 ( .IN1(n18652), .IN2(n2727), .IN3(n15515), .IN4(n2692), .Q(
        n15683) );
  OA22X1 U32078 ( .IN1(n18640), .IN2(n2587), .IN3(n18636), .IN4(n2552), .Q(
        n15684) );
  OA22X1 U32079 ( .IN1(n18626), .IN2(n2377), .IN3(n15525), .IN4(n2342), .Q(
        n15685) );
  OA22X1 U32080 ( .IN1(n18650), .IN2(n2726), .IN3(n18648), .IN4(n2691), .Q(
        n15595) );
  OA22X1 U32081 ( .IN1(n18638), .IN2(n2586), .IN3(n18636), .IN4(n2551), .Q(
        n15596) );
  OA22X1 U32082 ( .IN1(n18628), .IN2(n2376), .IN3(n18624), .IN4(n2341), .Q(
        n15597) );
  OA22X1 U32083 ( .IN1(n18651), .IN2(n2725), .IN3(n18648), .IN4(n2690), .Q(
        n15571) );
  OA22X1 U32084 ( .IN1(n18640), .IN2(n2585), .IN3(n18636), .IN4(n2550), .Q(
        n15572) );
  OA22X1 U32085 ( .IN1(n18627), .IN2(n2375), .IN3(n15525), .IN4(n2340), .Q(
        n15573) );
  OA22X1 U32086 ( .IN1(n18652), .IN2(n2724), .IN3(n18648), .IN4(n2689), .Q(
        n15563) );
  OA22X1 U32087 ( .IN1(n18638), .IN2(n2584), .IN3(n18635), .IN4(n2549), .Q(
        n15564) );
  OA22X1 U32088 ( .IN1(n18626), .IN2(n2374), .IN3(n18624), .IN4(n2339), .Q(
        n15565) );
  OA22X1 U32089 ( .IN1(n18650), .IN2(n2723), .IN3(n18648), .IN4(n2688), .Q(
        n15555) );
  OA22X1 U32090 ( .IN1(n18639), .IN2(n2583), .IN3(n15520), .IN4(n2548), .Q(
        n15556) );
  OA22X1 U32091 ( .IN1(n18626), .IN2(n2373), .IN3(n15525), .IN4(n2338), .Q(
        n15557) );
  OA22X1 U32092 ( .IN1(n18652), .IN2(n2722), .IN3(n18648), .IN4(n2687), .Q(
        n15547) );
  OA22X1 U32093 ( .IN1(n18640), .IN2(n2582), .IN3(n18636), .IN4(n2547), .Q(
        n15548) );
  OA22X1 U32094 ( .IN1(n18628), .IN2(n2372), .IN3(n18624), .IN4(n2337), .Q(
        n15549) );
  OA22X1 U32095 ( .IN1(n18650), .IN2(n2721), .IN3(n18648), .IN4(n2686), .Q(
        n15539) );
  OA22X1 U32096 ( .IN1(n18640), .IN2(n2581), .IN3(n18636), .IN4(n2546), .Q(
        n15540) );
  OA22X1 U32097 ( .IN1(n18628), .IN2(n2371), .IN3(n18624), .IN4(n2336), .Q(
        n15541) );
  OA22X1 U32098 ( .IN1(n18651), .IN2(n2720), .IN3(n18648), .IN4(n2685), .Q(
        n15531) );
  OA22X1 U32099 ( .IN1(n18640), .IN2(n2580), .IN3(n18636), .IN4(n2545), .Q(
        n15532) );
  OA22X1 U32100 ( .IN1(n18628), .IN2(n2370), .IN3(n18624), .IN4(n2335), .Q(
        n15533) );
  OA22X1 U32101 ( .IN1(n18652), .IN2(n2719), .IN3(n18648), .IN4(n2684), .Q(
        n15513) );
  OA22X1 U32102 ( .IN1(n18640), .IN2(n2579), .IN3(n18636), .IN4(n2544), .Q(
        n15518) );
  OA22X1 U32103 ( .IN1(n18628), .IN2(n2369), .IN3(n18624), .IN4(n2334), .Q(
        n15523) );
  OA22X1 U32104 ( .IN1(n18650), .IN2(n2718), .IN3(n18647), .IN4(n2683), .Q(
        n15763) );
  OA22X1 U32105 ( .IN1(n18639), .IN2(n2578), .IN3(n15520), .IN4(n2543), .Q(
        n15764) );
  OA22X1 U32106 ( .IN1(n18626), .IN2(n2368), .IN3(n18623), .IN4(n2333), .Q(
        n15765) );
  OA22X1 U32107 ( .IN1(n18650), .IN2(n2717), .IN3(n18647), .IN4(n2682), .Q(
        n15755) );
  OA22X1 U32108 ( .IN1(n18638), .IN2(n2577), .IN3(n15520), .IN4(n2542), .Q(
        n15756) );
  OA22X1 U32109 ( .IN1(n18627), .IN2(n2367), .IN3(n18623), .IN4(n2332), .Q(
        n15757) );
  OA22X1 U32110 ( .IN1(n18650), .IN2(n2716), .IN3(n18647), .IN4(n2681), .Q(
        n15747) );
  OA22X1 U32111 ( .IN1(n18639), .IN2(n2576), .IN3(n15520), .IN4(n2541), .Q(
        n15748) );
  OA22X1 U32112 ( .IN1(n18628), .IN2(n2366), .IN3(n18623), .IN4(n2331), .Q(
        n15749) );
  OA22X1 U32113 ( .IN1(n18651), .IN2(n2715), .IN3(n18647), .IN4(n2680), .Q(
        n15739) );
  OA22X1 U32114 ( .IN1(n18638), .IN2(n2575), .IN3(n18635), .IN4(n2540), .Q(
        n15740) );
  OA22X1 U32115 ( .IN1(n18626), .IN2(n2365), .IN3(n15525), .IN4(n2330), .Q(
        n15741) );
  OA22X1 U32116 ( .IN1(n18651), .IN2(n2714), .IN3(n18647), .IN4(n2679), .Q(
        n15731) );
  OA22X1 U32117 ( .IN1(n18638), .IN2(n2574), .IN3(n18635), .IN4(n2539), .Q(
        n15732) );
  OA22X1 U32118 ( .IN1(n18626), .IN2(n2364), .IN3(n15525), .IN4(n2329), .Q(
        n15733) );
  OA22X1 U32119 ( .IN1(n18651), .IN2(n2713), .IN3(n15515), .IN4(n2678), .Q(
        n15723) );
  OA22X1 U32120 ( .IN1(n18638), .IN2(n2573), .IN3(n18635), .IN4(n2538), .Q(
        n15724) );
  OA22X1 U32121 ( .IN1(n18626), .IN2(n2363), .IN3(n15525), .IN4(n2328), .Q(
        n15725) );
  OA22X1 U32122 ( .IN1(n18651), .IN2(n2712), .IN3(n15515), .IN4(n2677), .Q(
        n15715) );
  OA22X1 U32123 ( .IN1(n18638), .IN2(n2572), .IN3(n18635), .IN4(n2537), .Q(
        n15716) );
  OA22X1 U32124 ( .IN1(n18626), .IN2(n2362), .IN3(n15525), .IN4(n2327), .Q(
        n15717) );
  OA22X1 U32125 ( .IN1(n18652), .IN2(n2711), .IN3(n15515), .IN4(n2676), .Q(
        n15707) );
  OA22X1 U32126 ( .IN1(n18639), .IN2(n2571), .IN3(n18635), .IN4(n2536), .Q(
        n15708) );
  OA22X1 U32127 ( .IN1(n18627), .IN2(n2361), .IN3(n18623), .IN4(n2326), .Q(
        n15709) );
  OA22X1 U32128 ( .IN1(n18652), .IN2(n2710), .IN3(n15515), .IN4(n2675), .Q(
        n15699) );
  OA22X1 U32129 ( .IN1(n18639), .IN2(n2570), .IN3(n18636), .IN4(n2535), .Q(
        n15700) );
  OA22X1 U32130 ( .IN1(n18626), .IN2(n2360), .IN3(n15525), .IN4(n2325), .Q(
        n15701) );
  OA22X1 U32131 ( .IN1(n18652), .IN2(n2709), .IN3(n15515), .IN4(n2674), .Q(
        n15691) );
  OA22X1 U32132 ( .IN1(n18638), .IN2(n2569), .IN3(n18636), .IN4(n2534), .Q(
        n15692) );
  OA22X1 U32133 ( .IN1(n18627), .IN2(n2359), .IN3(n15525), .IN4(n2324), .Q(
        n15693) );
  OA22X1 U32134 ( .IN1(n18651), .IN2(n2708), .IN3(n15515), .IN4(n2673), .Q(
        n15675) );
  OA22X1 U32135 ( .IN1(n18639), .IN2(n2568), .IN3(n15520), .IN4(n2533), .Q(
        n15676) );
  OA22X1 U32136 ( .IN1(n18627), .IN2(n2358), .IN3(n15525), .IN4(n2323), .Q(
        n15677) );
  OA22X1 U32137 ( .IN1(n18651), .IN2(n2707), .IN3(n18648), .IN4(n2672), .Q(
        n15667) );
  OA22X1 U32138 ( .IN1(n18639), .IN2(n2567), .IN3(n15520), .IN4(n2532), .Q(
        n15668) );
  OA22X1 U32139 ( .IN1(n18627), .IN2(n2357), .IN3(n18624), .IN4(n2322), .Q(
        n15669) );
  OA22X1 U32140 ( .IN1(n18651), .IN2(n2706), .IN3(n18647), .IN4(n2671), .Q(
        n15659) );
  OA22X1 U32141 ( .IN1(n18639), .IN2(n2566), .IN3(n15520), .IN4(n2531), .Q(
        n15660) );
  OA22X1 U32142 ( .IN1(n18626), .IN2(n2356), .IN3(n18623), .IN4(n2321), .Q(
        n15661) );
  OA22X1 U32143 ( .IN1(n18652), .IN2(n2705), .IN3(n15515), .IN4(n2670), .Q(
        n15651) );
  OA22X1 U32144 ( .IN1(n18639), .IN2(n2565), .IN3(n15520), .IN4(n2530), .Q(
        n15652) );
  OA22X1 U32145 ( .IN1(n18626), .IN2(n2355), .IN3(n15525), .IN4(n2320), .Q(
        n15653) );
  OA22X1 U32146 ( .IN1(n18650), .IN2(n2704), .IN3(n18647), .IN4(n2669), .Q(
        n15643) );
  OA22X1 U32147 ( .IN1(n18639), .IN2(n2564), .IN3(n18635), .IN4(n2529), .Q(
        n15644) );
  OA22X1 U32148 ( .IN1(n18627), .IN2(n2354), .IN3(n18623), .IN4(n2319), .Q(
        n15645) );
  OA22X1 U32149 ( .IN1(n18650), .IN2(n2703), .IN3(n18647), .IN4(n2668), .Q(
        n15635) );
  OA22X1 U32150 ( .IN1(n18640), .IN2(n2563), .IN3(n18635), .IN4(n2528), .Q(
        n15636) );
  OA22X1 U32151 ( .IN1(n18627), .IN2(n2353), .IN3(n18623), .IN4(n2318), .Q(
        n15637) );
  OA22X1 U32152 ( .IN1(n18650), .IN2(n2702), .IN3(n15515), .IN4(n2667), .Q(
        n15627) );
  OA22X1 U32153 ( .IN1(n18639), .IN2(n2562), .IN3(n15520), .IN4(n2527), .Q(
        n15628) );
  OA22X1 U32154 ( .IN1(n18627), .IN2(n2352), .IN3(n18624), .IN4(n2317), .Q(
        n15629) );
  OA22X1 U32155 ( .IN1(n18652), .IN2(n2701), .IN3(n18647), .IN4(n2666), .Q(
        n15619) );
  OA22X1 U32156 ( .IN1(n18638), .IN2(n2561), .IN3(n15520), .IN4(n2526), .Q(
        n15620) );
  OA22X1 U32157 ( .IN1(n18627), .IN2(n2351), .IN3(n18623), .IN4(n2316), .Q(
        n15621) );
  OA22X1 U32158 ( .IN1(n18651), .IN2(n2700), .IN3(n15515), .IN4(n2665), .Q(
        n15611) );
  OA22X1 U32159 ( .IN1(n18640), .IN2(n2560), .IN3(n15520), .IN4(n2525), .Q(
        n15612) );
  OA22X1 U32160 ( .IN1(n18628), .IN2(n2350), .IN3(n15525), .IN4(n2315), .Q(
        n15613) );
  OA22X1 U32161 ( .IN1(n18652), .IN2(n2699), .IN3(n15515), .IN4(n2664), .Q(
        n15603) );
  OA22X1 U32162 ( .IN1(n18638), .IN2(n2559), .IN3(n18635), .IN4(n2524), .Q(
        n15604) );
  OA22X1 U32163 ( .IN1(n18627), .IN2(n2349), .IN3(n15525), .IN4(n2314), .Q(
        n15605) );
  OA22X1 U32164 ( .IN1(n18650), .IN2(n2698), .IN3(n15515), .IN4(n2663), .Q(
        n15587) );
  OA22X1 U32165 ( .IN1(n18640), .IN2(n2558), .IN3(n18636), .IN4(n2523), .Q(
        n15588) );
  OA22X1 U32166 ( .IN1(n18628), .IN2(n2348), .IN3(n15525), .IN4(n2313), .Q(
        n15589) );
  OA22X1 U32167 ( .IN1(n18651), .IN2(n2697), .IN3(n18648), .IN4(n2662), .Q(
        n15579) );
  OA22X1 U32168 ( .IN1(n18640), .IN2(n2557), .IN3(n18635), .IN4(n2522), .Q(
        n15580) );
  OA22X1 U32169 ( .IN1(n18628), .IN2(n2347), .IN3(n18624), .IN4(n2312), .Q(
        n15581) );
  OA22X1 U32170 ( .IN1(n18602), .IN2(n2728), .IN3(n18599), .IN4(n2693), .Q(
        n16076) );
  OA22X1 U32171 ( .IN1(n18590), .IN2(n2588), .IN3(n18587), .IN4(n2553), .Q(
        n16077) );
  OA22X1 U32172 ( .IN1(n18578), .IN2(n2378), .IN3(n18575), .IN4(n2343), .Q(
        n16078) );
  OA22X1 U32173 ( .IN1(n18604), .IN2(n2727), .IN3(n15820), .IN4(n2692), .Q(
        n15988) );
  OA22X1 U32174 ( .IN1(n18591), .IN2(n2587), .IN3(n18588), .IN4(n2552), .Q(
        n15989) );
  OA22X1 U32175 ( .IN1(n18579), .IN2(n2377), .IN3(n18576), .IN4(n2342), .Q(
        n15990) );
  OA22X1 U32176 ( .IN1(n18603), .IN2(n2726), .IN3(n18600), .IN4(n2691), .Q(
        n15900) );
  OA22X1 U32177 ( .IN1(n18591), .IN2(n2586), .IN3(n18589), .IN4(n2551), .Q(
        n15901) );
  OA22X1 U32178 ( .IN1(n18580), .IN2(n2376), .IN3(n15830), .IN4(n2341), .Q(
        n15902) );
  OA22X1 U32179 ( .IN1(n18602), .IN2(n2725), .IN3(n18600), .IN4(n2690), .Q(
        n15876) );
  OA22X1 U32180 ( .IN1(n18592), .IN2(n2585), .IN3(n18589), .IN4(n2550), .Q(
        n15877) );
  OA22X1 U32181 ( .IN1(n18578), .IN2(n2375), .IN3(n18576), .IN4(n2340), .Q(
        n15878) );
  OA22X1 U32182 ( .IN1(n18603), .IN2(n2724), .IN3(n18600), .IN4(n2689), .Q(
        n15868) );
  OA22X1 U32183 ( .IN1(n18590), .IN2(n2584), .IN3(n18589), .IN4(n2549), .Q(
        n15869) );
  OA22X1 U32184 ( .IN1(n18579), .IN2(n2374), .IN3(n18576), .IN4(n2339), .Q(
        n15870) );
  OA22X1 U32185 ( .IN1(n18604), .IN2(n2723), .IN3(n18600), .IN4(n2688), .Q(
        n15860) );
  OA22X1 U32186 ( .IN1(n18590), .IN2(n2583), .IN3(n18587), .IN4(n2548), .Q(
        n15861) );
  OA22X1 U32187 ( .IN1(n18580), .IN2(n2373), .IN3(n18576), .IN4(n2338), .Q(
        n15862) );
  OA22X1 U32188 ( .IN1(n18604), .IN2(n2722), .IN3(n18600), .IN4(n2687), .Q(
        n15852) );
  OA22X1 U32189 ( .IN1(n18592), .IN2(n2582), .IN3(n18589), .IN4(n2547), .Q(
        n15853) );
  OA22X1 U32190 ( .IN1(n18580), .IN2(n2372), .IN3(n18576), .IN4(n2337), .Q(
        n15854) );
  OA22X1 U32191 ( .IN1(n18604), .IN2(n2721), .IN3(n18600), .IN4(n2686), .Q(
        n15844) );
  OA22X1 U32192 ( .IN1(n18592), .IN2(n2581), .IN3(n18589), .IN4(n2546), .Q(
        n15845) );
  OA22X1 U32193 ( .IN1(n18580), .IN2(n2371), .IN3(n18576), .IN4(n2336), .Q(
        n15846) );
  OA22X1 U32194 ( .IN1(n18604), .IN2(n2720), .IN3(n18600), .IN4(n2685), .Q(
        n15836) );
  OA22X1 U32195 ( .IN1(n18592), .IN2(n2580), .IN3(n18589), .IN4(n2545), .Q(
        n15837) );
  OA22X1 U32196 ( .IN1(n18580), .IN2(n2370), .IN3(n18576), .IN4(n2335), .Q(
        n15838) );
  OA22X1 U32197 ( .IN1(n18604), .IN2(n2719), .IN3(n18600), .IN4(n2684), .Q(
        n15818) );
  OA22X1 U32198 ( .IN1(n18592), .IN2(n2579), .IN3(n18589), .IN4(n2544), .Q(
        n15823) );
  OA22X1 U32199 ( .IN1(n18580), .IN2(n2369), .IN3(n18576), .IN4(n2334), .Q(
        n15828) );
  OA22X1 U32200 ( .IN1(n18602), .IN2(n2718), .IN3(n18599), .IN4(n2683), .Q(
        n16068) );
  OA22X1 U32201 ( .IN1(n18590), .IN2(n2578), .IN3(n18587), .IN4(n2543), .Q(
        n16069) );
  OA22X1 U32202 ( .IN1(n18578), .IN2(n2368), .IN3(n18575), .IN4(n2333), .Q(
        n16070) );
  OA22X1 U32203 ( .IN1(n18602), .IN2(n2717), .IN3(n18599), .IN4(n2682), .Q(
        n16060) );
  OA22X1 U32204 ( .IN1(n18590), .IN2(n2577), .IN3(n18587), .IN4(n2542), .Q(
        n16061) );
  OA22X1 U32205 ( .IN1(n18578), .IN2(n2367), .IN3(n18575), .IN4(n2332), .Q(
        n16062) );
  OA22X1 U32206 ( .IN1(n18602), .IN2(n2716), .IN3(n18599), .IN4(n2681), .Q(
        n16052) );
  OA22X1 U32207 ( .IN1(n18590), .IN2(n2576), .IN3(n18587), .IN4(n2541), .Q(
        n16053) );
  OA22X1 U32208 ( .IN1(n18578), .IN2(n2366), .IN3(n18575), .IN4(n2331), .Q(
        n16054) );
  OA22X1 U32209 ( .IN1(n18602), .IN2(n2715), .IN3(n15820), .IN4(n2680), .Q(
        n16044) );
  OA22X1 U32210 ( .IN1(n18592), .IN2(n2575), .IN3(n18588), .IN4(n2540), .Q(
        n16045) );
  OA22X1 U32211 ( .IN1(n18578), .IN2(n2365), .IN3(n15830), .IN4(n2330), .Q(
        n16046) );
  OA22X1 U32212 ( .IN1(n18602), .IN2(n2714), .IN3(n15820), .IN4(n2679), .Q(
        n16036) );
  OA22X1 U32213 ( .IN1(n18590), .IN2(n2574), .IN3(n18588), .IN4(n2539), .Q(
        n16037) );
  OA22X1 U32214 ( .IN1(n18579), .IN2(n2364), .IN3(n15830), .IN4(n2329), .Q(
        n16038) );
  OA22X1 U32215 ( .IN1(n18604), .IN2(n2713), .IN3(n15820), .IN4(n2678), .Q(
        n16028) );
  OA22X1 U32216 ( .IN1(n18591), .IN2(n2573), .IN3(n18588), .IN4(n2538), .Q(
        n16029) );
  OA22X1 U32217 ( .IN1(n18580), .IN2(n2363), .IN3(n15830), .IN4(n2328), .Q(
        n16030) );
  OA22X1 U32218 ( .IN1(n18602), .IN2(n2712), .IN3(n15820), .IN4(n2677), .Q(
        n16020) );
  OA22X1 U32219 ( .IN1(n18592), .IN2(n2572), .IN3(n18588), .IN4(n2537), .Q(
        n16021) );
  OA22X1 U32220 ( .IN1(n18580), .IN2(n2362), .IN3(n15830), .IN4(n2327), .Q(
        n16022) );
  OA22X1 U32221 ( .IN1(n18602), .IN2(n2711), .IN3(n15820), .IN4(n2676), .Q(
        n16012) );
  OA22X1 U32222 ( .IN1(n18592), .IN2(n2571), .IN3(n18589), .IN4(n2536), .Q(
        n16013) );
  OA22X1 U32223 ( .IN1(n18579), .IN2(n2361), .IN3(n15830), .IN4(n2326), .Q(
        n16014) );
  OA22X1 U32224 ( .IN1(n18604), .IN2(n2710), .IN3(n15820), .IN4(n2675), .Q(
        n16004) );
  OA22X1 U32225 ( .IN1(n18590), .IN2(n2570), .IN3(n18587), .IN4(n2535), .Q(
        n16005) );
  OA22X1 U32226 ( .IN1(n18579), .IN2(n2360), .IN3(n15830), .IN4(n2325), .Q(
        n16006) );
  OA22X1 U32227 ( .IN1(n18602), .IN2(n2709), .IN3(n15820), .IN4(n2674), .Q(
        n15996) );
  OA22X1 U32228 ( .IN1(n18592), .IN2(n2569), .IN3(n18588), .IN4(n2534), .Q(
        n15997) );
  OA22X1 U32229 ( .IN1(n18579), .IN2(n2359), .IN3(n15830), .IN4(n2324), .Q(
        n15998) );
  OA22X1 U32230 ( .IN1(n18603), .IN2(n2708), .IN3(n18599), .IN4(n2673), .Q(
        n15980) );
  OA22X1 U32231 ( .IN1(n18592), .IN2(n2568), .IN3(n18587), .IN4(n2533), .Q(
        n15981) );
  OA22X1 U32232 ( .IN1(n18578), .IN2(n2358), .IN3(n18575), .IN4(n2323), .Q(
        n15982) );
  OA22X1 U32233 ( .IN1(n18603), .IN2(n2707), .IN3(n15820), .IN4(n2672), .Q(
        n15972) );
  OA22X1 U32234 ( .IN1(n18592), .IN2(n2567), .IN3(n18588), .IN4(n2532), .Q(
        n15973) );
  OA22X1 U32235 ( .IN1(n18578), .IN2(n2357), .IN3(n18576), .IN4(n2322), .Q(
        n15974) );
  OA22X1 U32236 ( .IN1(n18603), .IN2(n2706), .IN3(n18599), .IN4(n2671), .Q(
        n15964) );
  OA22X1 U32237 ( .IN1(n18590), .IN2(n2566), .IN3(n18589), .IN4(n2531), .Q(
        n15965) );
  OA22X1 U32238 ( .IN1(n18579), .IN2(n2356), .IN3(n18575), .IN4(n2321), .Q(
        n15966) );
  OA22X1 U32239 ( .IN1(n18603), .IN2(n2705), .IN3(n18599), .IN4(n2670), .Q(
        n15956) );
  OA22X1 U32240 ( .IN1(n18591), .IN2(n2565), .IN3(n18587), .IN4(n2530), .Q(
        n15957) );
  OA22X1 U32241 ( .IN1(n18579), .IN2(n2355), .IN3(n15830), .IN4(n2320), .Q(
        n15958) );
  OA22X1 U32242 ( .IN1(n18603), .IN2(n2704), .IN3(n18599), .IN4(n2669), .Q(
        n15948) );
  OA22X1 U32243 ( .IN1(n18591), .IN2(n2564), .IN3(n18587), .IN4(n2529), .Q(
        n15949) );
  OA22X1 U32244 ( .IN1(n18579), .IN2(n2354), .IN3(n18575), .IN4(n2319), .Q(
        n15950) );
  OA22X1 U32245 ( .IN1(n18604), .IN2(n2703), .IN3(n18599), .IN4(n2668), .Q(
        n15940) );
  OA22X1 U32246 ( .IN1(n18591), .IN2(n2563), .IN3(n18588), .IN4(n2528), .Q(
        n15941) );
  OA22X1 U32247 ( .IN1(n18580), .IN2(n2353), .IN3(n18575), .IN4(n2318), .Q(
        n15942) );
  OA22X1 U32248 ( .IN1(n18603), .IN2(n2702), .IN3(n15820), .IN4(n2667), .Q(
        n15932) );
  OA22X1 U32249 ( .IN1(n18591), .IN2(n2562), .IN3(n18589), .IN4(n2527), .Q(
        n15933) );
  OA22X1 U32250 ( .IN1(n18579), .IN2(n2352), .IN3(n15830), .IN4(n2317), .Q(
        n15934) );
  OA22X1 U32251 ( .IN1(n18604), .IN2(n2701), .IN3(n18599), .IN4(n2666), .Q(
        n15924) );
  OA22X1 U32252 ( .IN1(n18591), .IN2(n2561), .IN3(n18587), .IN4(n2526), .Q(
        n15925) );
  OA22X1 U32253 ( .IN1(n18578), .IN2(n2351), .IN3(n18575), .IN4(n2316), .Q(
        n15926) );
  OA22X1 U32254 ( .IN1(n18603), .IN2(n2700), .IN3(n18600), .IN4(n2665), .Q(
        n15916) );
  OA22X1 U32255 ( .IN1(n18591), .IN2(n2560), .IN3(n18587), .IN4(n2525), .Q(
        n15917) );
  OA22X1 U32256 ( .IN1(n18580), .IN2(n2350), .IN3(n15830), .IN4(n2315), .Q(
        n15918) );
  OA22X1 U32257 ( .IN1(n18603), .IN2(n2699), .IN3(n15820), .IN4(n2664), .Q(
        n15908) );
  OA22X1 U32258 ( .IN1(n18591), .IN2(n2559), .IN3(n18588), .IN4(n2524), .Q(
        n15909) );
  OA22X1 U32259 ( .IN1(n18578), .IN2(n2349), .IN3(n15830), .IN4(n2314), .Q(
        n15910) );
  OA22X1 U32260 ( .IN1(n18604), .IN2(n2698), .IN3(n18600), .IN4(n2663), .Q(
        n15892) );
  OA22X1 U32261 ( .IN1(n18591), .IN2(n2558), .IN3(n18589), .IN4(n2523), .Q(
        n15893) );
  OA22X1 U32262 ( .IN1(n18580), .IN2(n2348), .IN3(n15830), .IN4(n2313), .Q(
        n15894) );
  OA22X1 U32263 ( .IN1(n18603), .IN2(n2697), .IN3(n15820), .IN4(n2662), .Q(
        n15884) );
  OA22X1 U32264 ( .IN1(n18590), .IN2(n2557), .IN3(n18588), .IN4(n2522), .Q(
        n15885) );
  OA22X1 U32265 ( .IN1(n18578), .IN2(n2347), .IN3(n15830), .IN4(n2312), .Q(
        n15886) );
  OA22X1 U32266 ( .IN1(n18554), .IN2(n2728), .IN3(n18551), .IN4(n2693), .Q(
        n16381) );
  OA22X1 U32267 ( .IN1(n18542), .IN2(n2588), .IN3(n16130), .IN4(n2553), .Q(
        n16382) );
  OA22X1 U32268 ( .IN1(n18532), .IN2(n2378), .IN3(n18527), .IN4(n2343), .Q(
        n16383) );
  OA22X1 U32269 ( .IN1(n18556), .IN2(n2727), .IN3(n16125), .IN4(n2692), .Q(
        n16293) );
  OA22X1 U32270 ( .IN1(n18544), .IN2(n2587), .IN3(n18540), .IN4(n2552), .Q(
        n16294) );
  OA22X1 U32271 ( .IN1(n18530), .IN2(n2377), .IN3(n16135), .IN4(n2342), .Q(
        n16295) );
  OA22X1 U32272 ( .IN1(n18554), .IN2(n2726), .IN3(n18552), .IN4(n2691), .Q(
        n16205) );
  OA22X1 U32273 ( .IN1(n18542), .IN2(n2586), .IN3(n18540), .IN4(n2551), .Q(
        n16206) );
  OA22X1 U32274 ( .IN1(n18532), .IN2(n2376), .IN3(n18528), .IN4(n2341), .Q(
        n16207) );
  OA22X1 U32275 ( .IN1(n18555), .IN2(n2725), .IN3(n18552), .IN4(n2690), .Q(
        n16181) );
  OA22X1 U32276 ( .IN1(n18544), .IN2(n2585), .IN3(n18540), .IN4(n2550), .Q(
        n16182) );
  OA22X1 U32277 ( .IN1(n18531), .IN2(n2375), .IN3(n16135), .IN4(n2340), .Q(
        n16183) );
  OA22X1 U32278 ( .IN1(n18556), .IN2(n2724), .IN3(n18552), .IN4(n2689), .Q(
        n16173) );
  OA22X1 U32279 ( .IN1(n18542), .IN2(n2584), .IN3(n18539), .IN4(n2549), .Q(
        n16174) );
  OA22X1 U32280 ( .IN1(n18530), .IN2(n2374), .IN3(n18528), .IN4(n2339), .Q(
        n16175) );
  OA22X1 U32281 ( .IN1(n18554), .IN2(n2723), .IN3(n18552), .IN4(n2688), .Q(
        n16165) );
  OA22X1 U32282 ( .IN1(n18543), .IN2(n2583), .IN3(n16130), .IN4(n2548), .Q(
        n16166) );
  OA22X1 U32283 ( .IN1(n18530), .IN2(n2373), .IN3(n16135), .IN4(n2338), .Q(
        n16167) );
  OA22X1 U32284 ( .IN1(n18556), .IN2(n2722), .IN3(n18552), .IN4(n2687), .Q(
        n16157) );
  OA22X1 U32285 ( .IN1(n18544), .IN2(n2582), .IN3(n18540), .IN4(n2547), .Q(
        n16158) );
  OA22X1 U32286 ( .IN1(n18532), .IN2(n2372), .IN3(n18528), .IN4(n2337), .Q(
        n16159) );
  OA22X1 U32287 ( .IN1(n18554), .IN2(n2721), .IN3(n18552), .IN4(n2686), .Q(
        n16149) );
  OA22X1 U32288 ( .IN1(n18544), .IN2(n2581), .IN3(n18540), .IN4(n2546), .Q(
        n16150) );
  OA22X1 U32289 ( .IN1(n18532), .IN2(n2371), .IN3(n18528), .IN4(n2336), .Q(
        n16151) );
  OA22X1 U32290 ( .IN1(n18555), .IN2(n2720), .IN3(n18552), .IN4(n2685), .Q(
        n16141) );
  OA22X1 U32291 ( .IN1(n18544), .IN2(n2580), .IN3(n18540), .IN4(n2545), .Q(
        n16142) );
  OA22X1 U32292 ( .IN1(n18532), .IN2(n2370), .IN3(n18528), .IN4(n2335), .Q(
        n16143) );
  OA22X1 U32293 ( .IN1(n18556), .IN2(n2719), .IN3(n18552), .IN4(n2684), .Q(
        n16123) );
  OA22X1 U32294 ( .IN1(n18544), .IN2(n2579), .IN3(n18540), .IN4(n2544), .Q(
        n16128) );
  OA22X1 U32295 ( .IN1(n18532), .IN2(n2369), .IN3(n18528), .IN4(n2334), .Q(
        n16133) );
  OA22X1 U32296 ( .IN1(n18554), .IN2(n2718), .IN3(n18551), .IN4(n2683), .Q(
        n16373) );
  OA22X1 U32297 ( .IN1(n18543), .IN2(n2578), .IN3(n16130), .IN4(n2543), .Q(
        n16374) );
  OA22X1 U32298 ( .IN1(n18530), .IN2(n2368), .IN3(n18527), .IN4(n2333), .Q(
        n16375) );
  OA22X1 U32299 ( .IN1(n18554), .IN2(n2717), .IN3(n18551), .IN4(n2682), .Q(
        n16365) );
  OA22X1 U32300 ( .IN1(n18542), .IN2(n2577), .IN3(n16130), .IN4(n2542), .Q(
        n16366) );
  OA22X1 U32301 ( .IN1(n18531), .IN2(n2367), .IN3(n18527), .IN4(n2332), .Q(
        n16367) );
  OA22X1 U32302 ( .IN1(n18554), .IN2(n2716), .IN3(n18551), .IN4(n2681), .Q(
        n16357) );
  OA22X1 U32303 ( .IN1(n18543), .IN2(n2576), .IN3(n16130), .IN4(n2541), .Q(
        n16358) );
  OA22X1 U32304 ( .IN1(n18532), .IN2(n2366), .IN3(n18527), .IN4(n2331), .Q(
        n16359) );
  OA22X1 U32305 ( .IN1(n18555), .IN2(n2715), .IN3(n18551), .IN4(n2680), .Q(
        n16349) );
  OA22X1 U32306 ( .IN1(n18542), .IN2(n2575), .IN3(n18539), .IN4(n2540), .Q(
        n16350) );
  OA22X1 U32307 ( .IN1(n18530), .IN2(n2365), .IN3(n16135), .IN4(n2330), .Q(
        n16351) );
  OA22X1 U32308 ( .IN1(n18555), .IN2(n2714), .IN3(n18551), .IN4(n2679), .Q(
        n16341) );
  OA22X1 U32309 ( .IN1(n18542), .IN2(n2574), .IN3(n18539), .IN4(n2539), .Q(
        n16342) );
  OA22X1 U32310 ( .IN1(n18530), .IN2(n2364), .IN3(n16135), .IN4(n2329), .Q(
        n16343) );
  OA22X1 U32311 ( .IN1(n18555), .IN2(n2713), .IN3(n16125), .IN4(n2678), .Q(
        n16333) );
  OA22X1 U32312 ( .IN1(n18542), .IN2(n2573), .IN3(n18539), .IN4(n2538), .Q(
        n16334) );
  OA22X1 U32313 ( .IN1(n18530), .IN2(n2363), .IN3(n16135), .IN4(n2328), .Q(
        n16335) );
  OA22X1 U32314 ( .IN1(n18555), .IN2(n2712), .IN3(n16125), .IN4(n2677), .Q(
        n16325) );
  OA22X1 U32315 ( .IN1(n18542), .IN2(n2572), .IN3(n18539), .IN4(n2537), .Q(
        n16326) );
  OA22X1 U32316 ( .IN1(n18530), .IN2(n2362), .IN3(n16135), .IN4(n2327), .Q(
        n16327) );
  OA22X1 U32317 ( .IN1(n18556), .IN2(n2711), .IN3(n16125), .IN4(n2676), .Q(
        n16317) );
  OA22X1 U32318 ( .IN1(n18543), .IN2(n2571), .IN3(n18539), .IN4(n2536), .Q(
        n16318) );
  OA22X1 U32319 ( .IN1(n18531), .IN2(n2361), .IN3(n18527), .IN4(n2326), .Q(
        n16319) );
  OA22X1 U32320 ( .IN1(n18556), .IN2(n2710), .IN3(n16125), .IN4(n2675), .Q(
        n16309) );
  OA22X1 U32321 ( .IN1(n18543), .IN2(n2570), .IN3(n18540), .IN4(n2535), .Q(
        n16310) );
  OA22X1 U32322 ( .IN1(n18530), .IN2(n2360), .IN3(n16135), .IN4(n2325), .Q(
        n16311) );
  OA22X1 U32323 ( .IN1(n18556), .IN2(n2709), .IN3(n16125), .IN4(n2674), .Q(
        n16301) );
  OA22X1 U32324 ( .IN1(n18542), .IN2(n2569), .IN3(n18540), .IN4(n2534), .Q(
        n16302) );
  OA22X1 U32325 ( .IN1(n18531), .IN2(n2359), .IN3(n16135), .IN4(n2324), .Q(
        n16303) );
  OA22X1 U32326 ( .IN1(n18555), .IN2(n2708), .IN3(n16125), .IN4(n2673), .Q(
        n16285) );
  OA22X1 U32327 ( .IN1(n18543), .IN2(n2568), .IN3(n16130), .IN4(n2533), .Q(
        n16286) );
  OA22X1 U32328 ( .IN1(n18531), .IN2(n2358), .IN3(n16135), .IN4(n2323), .Q(
        n16287) );
  OA22X1 U32329 ( .IN1(n18555), .IN2(n2707), .IN3(n18552), .IN4(n2672), .Q(
        n16277) );
  OA22X1 U32330 ( .IN1(n18543), .IN2(n2567), .IN3(n16130), .IN4(n2532), .Q(
        n16278) );
  OA22X1 U32331 ( .IN1(n18531), .IN2(n2357), .IN3(n18528), .IN4(n2322), .Q(
        n16279) );
  OA22X1 U32332 ( .IN1(n18555), .IN2(n2706), .IN3(n18551), .IN4(n2671), .Q(
        n16269) );
  OA22X1 U32333 ( .IN1(n18543), .IN2(n2566), .IN3(n16130), .IN4(n2531), .Q(
        n16270) );
  OA22X1 U32334 ( .IN1(n18530), .IN2(n2356), .IN3(n18527), .IN4(n2321), .Q(
        n16271) );
  OA22X1 U32335 ( .IN1(n18556), .IN2(n2705), .IN3(n16125), .IN4(n2670), .Q(
        n16261) );
  OA22X1 U32336 ( .IN1(n18543), .IN2(n2565), .IN3(n16130), .IN4(n2530), .Q(
        n16262) );
  OA22X1 U32337 ( .IN1(n18530), .IN2(n2355), .IN3(n16135), .IN4(n2320), .Q(
        n16263) );
  OA22X1 U32338 ( .IN1(n18554), .IN2(n2704), .IN3(n18551), .IN4(n2669), .Q(
        n16253) );
  OA22X1 U32339 ( .IN1(n18543), .IN2(n2564), .IN3(n18539), .IN4(n2529), .Q(
        n16254) );
  OA22X1 U32340 ( .IN1(n18531), .IN2(n2354), .IN3(n18527), .IN4(n2319), .Q(
        n16255) );
  OA22X1 U32341 ( .IN1(n18554), .IN2(n2703), .IN3(n18551), .IN4(n2668), .Q(
        n16245) );
  OA22X1 U32342 ( .IN1(n18544), .IN2(n2563), .IN3(n18539), .IN4(n2528), .Q(
        n16246) );
  OA22X1 U32343 ( .IN1(n18531), .IN2(n2353), .IN3(n18527), .IN4(n2318), .Q(
        n16247) );
  OA22X1 U32344 ( .IN1(n18554), .IN2(n2702), .IN3(n16125), .IN4(n2667), .Q(
        n16237) );
  OA22X1 U32345 ( .IN1(n18543), .IN2(n2562), .IN3(n16130), .IN4(n2527), .Q(
        n16238) );
  OA22X1 U32346 ( .IN1(n18531), .IN2(n2352), .IN3(n18528), .IN4(n2317), .Q(
        n16239) );
  OA22X1 U32347 ( .IN1(n18556), .IN2(n2701), .IN3(n18551), .IN4(n2666), .Q(
        n16229) );
  OA22X1 U32348 ( .IN1(n18542), .IN2(n2561), .IN3(n16130), .IN4(n2526), .Q(
        n16230) );
  OA22X1 U32349 ( .IN1(n18531), .IN2(n2351), .IN3(n18527), .IN4(n2316), .Q(
        n16231) );
  OA22X1 U32350 ( .IN1(n18555), .IN2(n2700), .IN3(n16125), .IN4(n2665), .Q(
        n16221) );
  OA22X1 U32351 ( .IN1(n18544), .IN2(n2560), .IN3(n16130), .IN4(n2525), .Q(
        n16222) );
  OA22X1 U32352 ( .IN1(n18532), .IN2(n2350), .IN3(n16135), .IN4(n2315), .Q(
        n16223) );
  OA22X1 U32353 ( .IN1(n18556), .IN2(n2699), .IN3(n16125), .IN4(n2664), .Q(
        n16213) );
  OA22X1 U32354 ( .IN1(n18542), .IN2(n2559), .IN3(n18539), .IN4(n2524), .Q(
        n16214) );
  OA22X1 U32355 ( .IN1(n18531), .IN2(n2349), .IN3(n16135), .IN4(n2314), .Q(
        n16215) );
  OA22X1 U32356 ( .IN1(n18554), .IN2(n2698), .IN3(n16125), .IN4(n2663), .Q(
        n16197) );
  OA22X1 U32357 ( .IN1(n18544), .IN2(n2558), .IN3(n18540), .IN4(n2523), .Q(
        n16198) );
  OA22X1 U32358 ( .IN1(n18532), .IN2(n2348), .IN3(n16135), .IN4(n2313), .Q(
        n16199) );
  OA22X1 U32359 ( .IN1(n18555), .IN2(n2697), .IN3(n18552), .IN4(n2662), .Q(
        n16189) );
  OA22X1 U32360 ( .IN1(n18544), .IN2(n2557), .IN3(n18539), .IN4(n2522), .Q(
        n16190) );
  OA22X1 U32361 ( .IN1(n18532), .IN2(n2347), .IN3(n18528), .IN4(n2312), .Q(
        n16191) );
  OA22X1 U32362 ( .IN1(n18506), .IN2(n2728), .IN3(n18503), .IN4(n2693), .Q(
        n16686) );
  OA22X1 U32363 ( .IN1(n18494), .IN2(n2588), .IN3(n18491), .IN4(n2553), .Q(
        n16687) );
  OA22X1 U32364 ( .IN1(n18482), .IN2(n2378), .IN3(n18479), .IN4(n2343), .Q(
        n16688) );
  OA22X1 U32365 ( .IN1(n18508), .IN2(n2727), .IN3(n16430), .IN4(n2692), .Q(
        n16598) );
  OA22X1 U32366 ( .IN1(n18495), .IN2(n2587), .IN3(n18492), .IN4(n2552), .Q(
        n16599) );
  OA22X1 U32367 ( .IN1(n18483), .IN2(n2377), .IN3(n18480), .IN4(n2342), .Q(
        n16600) );
  OA22X1 U32368 ( .IN1(n18507), .IN2(n2726), .IN3(n18504), .IN4(n2691), .Q(
        n16510) );
  OA22X1 U32369 ( .IN1(n18495), .IN2(n2586), .IN3(n18493), .IN4(n2551), .Q(
        n16511) );
  OA22X1 U32370 ( .IN1(n18484), .IN2(n2376), .IN3(n16440), .IN4(n2341), .Q(
        n16512) );
  OA22X1 U32371 ( .IN1(n18506), .IN2(n2725), .IN3(n18504), .IN4(n2690), .Q(
        n16486) );
  OA22X1 U32372 ( .IN1(n18496), .IN2(n2585), .IN3(n18493), .IN4(n2550), .Q(
        n16487) );
  OA22X1 U32373 ( .IN1(n18482), .IN2(n2375), .IN3(n18480), .IN4(n2340), .Q(
        n16488) );
  OA22X1 U32374 ( .IN1(n18507), .IN2(n2724), .IN3(n18504), .IN4(n2689), .Q(
        n16478) );
  OA22X1 U32375 ( .IN1(n18494), .IN2(n2584), .IN3(n18493), .IN4(n2549), .Q(
        n16479) );
  OA22X1 U32376 ( .IN1(n18483), .IN2(n2374), .IN3(n18480), .IN4(n2339), .Q(
        n16480) );
  OA22X1 U32377 ( .IN1(n18508), .IN2(n2723), .IN3(n18504), .IN4(n2688), .Q(
        n16470) );
  OA22X1 U32378 ( .IN1(n18494), .IN2(n2583), .IN3(n18491), .IN4(n2548), .Q(
        n16471) );
  OA22X1 U32379 ( .IN1(n18484), .IN2(n2373), .IN3(n18480), .IN4(n2338), .Q(
        n16472) );
  OA22X1 U32380 ( .IN1(n18508), .IN2(n2722), .IN3(n18504), .IN4(n2687), .Q(
        n16462) );
  OA22X1 U32381 ( .IN1(n18496), .IN2(n2582), .IN3(n18493), .IN4(n2547), .Q(
        n16463) );
  OA22X1 U32382 ( .IN1(n18484), .IN2(n2372), .IN3(n18480), .IN4(n2337), .Q(
        n16464) );
  OA22X1 U32383 ( .IN1(n18508), .IN2(n2721), .IN3(n18504), .IN4(n2686), .Q(
        n16454) );
  OA22X1 U32384 ( .IN1(n18496), .IN2(n2581), .IN3(n18493), .IN4(n2546), .Q(
        n16455) );
  OA22X1 U32385 ( .IN1(n18484), .IN2(n2371), .IN3(n18480), .IN4(n2336), .Q(
        n16456) );
  OA22X1 U32386 ( .IN1(n18508), .IN2(n2720), .IN3(n18504), .IN4(n2685), .Q(
        n16446) );
  OA22X1 U32387 ( .IN1(n18496), .IN2(n2580), .IN3(n18493), .IN4(n2545), .Q(
        n16447) );
  OA22X1 U32388 ( .IN1(n18484), .IN2(n2370), .IN3(n18480), .IN4(n2335), .Q(
        n16448) );
  OA22X1 U32389 ( .IN1(n18508), .IN2(n2719), .IN3(n18504), .IN4(n2684), .Q(
        n16428) );
  OA22X1 U32390 ( .IN1(n18496), .IN2(n2579), .IN3(n18493), .IN4(n2544), .Q(
        n16433) );
  OA22X1 U32391 ( .IN1(n18484), .IN2(n2369), .IN3(n18480), .IN4(n2334), .Q(
        n16438) );
  OA22X1 U32392 ( .IN1(n18506), .IN2(n2718), .IN3(n18503), .IN4(n2683), .Q(
        n16678) );
  OA22X1 U32393 ( .IN1(n18494), .IN2(n2578), .IN3(n18491), .IN4(n2543), .Q(
        n16679) );
  OA22X1 U32394 ( .IN1(n18482), .IN2(n2368), .IN3(n18479), .IN4(n2333), .Q(
        n16680) );
  OA22X1 U32395 ( .IN1(n18506), .IN2(n2717), .IN3(n18503), .IN4(n2682), .Q(
        n16670) );
  OA22X1 U32396 ( .IN1(n18494), .IN2(n2577), .IN3(n18491), .IN4(n2542), .Q(
        n16671) );
  OA22X1 U32397 ( .IN1(n18482), .IN2(n2367), .IN3(n18479), .IN4(n2332), .Q(
        n16672) );
  OA22X1 U32398 ( .IN1(n18506), .IN2(n2716), .IN3(n18503), .IN4(n2681), .Q(
        n16662) );
  OA22X1 U32399 ( .IN1(n18494), .IN2(n2576), .IN3(n18491), .IN4(n2541), .Q(
        n16663) );
  OA22X1 U32400 ( .IN1(n18482), .IN2(n2366), .IN3(n18479), .IN4(n2331), .Q(
        n16664) );
  OA22X1 U32401 ( .IN1(n18506), .IN2(n2715), .IN3(n16430), .IN4(n2680), .Q(
        n16654) );
  OA22X1 U32402 ( .IN1(n18496), .IN2(n2575), .IN3(n18492), .IN4(n2540), .Q(
        n16655) );
  OA22X1 U32403 ( .IN1(n18482), .IN2(n2365), .IN3(n16440), .IN4(n2330), .Q(
        n16656) );
  OA22X1 U32404 ( .IN1(n18506), .IN2(n2714), .IN3(n16430), .IN4(n2679), .Q(
        n16646) );
  OA22X1 U32405 ( .IN1(n18494), .IN2(n2574), .IN3(n18492), .IN4(n2539), .Q(
        n16647) );
  OA22X1 U32406 ( .IN1(n18483), .IN2(n2364), .IN3(n16440), .IN4(n2329), .Q(
        n16648) );
  OA22X1 U32407 ( .IN1(n18508), .IN2(n2713), .IN3(n16430), .IN4(n2678), .Q(
        n16638) );
  OA22X1 U32408 ( .IN1(n18495), .IN2(n2573), .IN3(n18492), .IN4(n2538), .Q(
        n16639) );
  OA22X1 U32409 ( .IN1(n18484), .IN2(n2363), .IN3(n16440), .IN4(n2328), .Q(
        n16640) );
  OA22X1 U32410 ( .IN1(n18506), .IN2(n2712), .IN3(n16430), .IN4(n2677), .Q(
        n16630) );
  OA22X1 U32411 ( .IN1(n18496), .IN2(n2572), .IN3(n18492), .IN4(n2537), .Q(
        n16631) );
  OA22X1 U32412 ( .IN1(n18484), .IN2(n2362), .IN3(n16440), .IN4(n2327), .Q(
        n16632) );
  OA22X1 U32413 ( .IN1(n18506), .IN2(n2711), .IN3(n16430), .IN4(n2676), .Q(
        n16622) );
  OA22X1 U32414 ( .IN1(n18496), .IN2(n2571), .IN3(n18493), .IN4(n2536), .Q(
        n16623) );
  OA22X1 U32415 ( .IN1(n18483), .IN2(n2361), .IN3(n16440), .IN4(n2326), .Q(
        n16624) );
  OA22X1 U32416 ( .IN1(n18508), .IN2(n2710), .IN3(n16430), .IN4(n2675), .Q(
        n16614) );
  OA22X1 U32417 ( .IN1(n18494), .IN2(n2570), .IN3(n18491), .IN4(n2535), .Q(
        n16615) );
  OA22X1 U32418 ( .IN1(n18483), .IN2(n2360), .IN3(n16440), .IN4(n2325), .Q(
        n16616) );
  OA22X1 U32419 ( .IN1(n18506), .IN2(n2709), .IN3(n16430), .IN4(n2674), .Q(
        n16606) );
  OA22X1 U32420 ( .IN1(n18496), .IN2(n2569), .IN3(n18492), .IN4(n2534), .Q(
        n16607) );
  OA22X1 U32421 ( .IN1(n18483), .IN2(n2359), .IN3(n16440), .IN4(n2324), .Q(
        n16608) );
  OA22X1 U32422 ( .IN1(n18507), .IN2(n2708), .IN3(n18503), .IN4(n2673), .Q(
        n16590) );
  OA22X1 U32423 ( .IN1(n18496), .IN2(n2568), .IN3(n18491), .IN4(n2533), .Q(
        n16591) );
  OA22X1 U32424 ( .IN1(n18482), .IN2(n2358), .IN3(n18479), .IN4(n2323), .Q(
        n16592) );
  OA22X1 U32425 ( .IN1(n18507), .IN2(n2707), .IN3(n16430), .IN4(n2672), .Q(
        n16582) );
  OA22X1 U32426 ( .IN1(n18496), .IN2(n2567), .IN3(n18492), .IN4(n2532), .Q(
        n16583) );
  OA22X1 U32427 ( .IN1(n18482), .IN2(n2357), .IN3(n18480), .IN4(n2322), .Q(
        n16584) );
  OA22X1 U32428 ( .IN1(n18507), .IN2(n2706), .IN3(n18503), .IN4(n2671), .Q(
        n16574) );
  OA22X1 U32429 ( .IN1(n18494), .IN2(n2566), .IN3(n18493), .IN4(n2531), .Q(
        n16575) );
  OA22X1 U32430 ( .IN1(n18483), .IN2(n2356), .IN3(n18479), .IN4(n2321), .Q(
        n16576) );
  OA22X1 U32431 ( .IN1(n18507), .IN2(n2705), .IN3(n18503), .IN4(n2670), .Q(
        n16566) );
  OA22X1 U32432 ( .IN1(n18495), .IN2(n2565), .IN3(n18491), .IN4(n2530), .Q(
        n16567) );
  OA22X1 U32433 ( .IN1(n18483), .IN2(n2355), .IN3(n16440), .IN4(n2320), .Q(
        n16568) );
  OA22X1 U32434 ( .IN1(n18507), .IN2(n2704), .IN3(n18503), .IN4(n2669), .Q(
        n16558) );
  OA22X1 U32435 ( .IN1(n18495), .IN2(n2564), .IN3(n18491), .IN4(n2529), .Q(
        n16559) );
  OA22X1 U32436 ( .IN1(n18483), .IN2(n2354), .IN3(n18479), .IN4(n2319), .Q(
        n16560) );
  OA22X1 U32437 ( .IN1(n18508), .IN2(n2703), .IN3(n18503), .IN4(n2668), .Q(
        n16550) );
  OA22X1 U32438 ( .IN1(n18495), .IN2(n2563), .IN3(n18492), .IN4(n2528), .Q(
        n16551) );
  OA22X1 U32439 ( .IN1(n18484), .IN2(n2353), .IN3(n18479), .IN4(n2318), .Q(
        n16552) );
  OA22X1 U32440 ( .IN1(n18507), .IN2(n2702), .IN3(n16430), .IN4(n2667), .Q(
        n16542) );
  OA22X1 U32441 ( .IN1(n18495), .IN2(n2562), .IN3(n18493), .IN4(n2527), .Q(
        n16543) );
  OA22X1 U32442 ( .IN1(n18483), .IN2(n2352), .IN3(n16440), .IN4(n2317), .Q(
        n16544) );
  OA22X1 U32443 ( .IN1(n18508), .IN2(n2701), .IN3(n18503), .IN4(n2666), .Q(
        n16534) );
  OA22X1 U32444 ( .IN1(n18495), .IN2(n2561), .IN3(n18491), .IN4(n2526), .Q(
        n16535) );
  OA22X1 U32445 ( .IN1(n18482), .IN2(n2351), .IN3(n18479), .IN4(n2316), .Q(
        n16536) );
  OA22X1 U32446 ( .IN1(n18507), .IN2(n2700), .IN3(n18504), .IN4(n2665), .Q(
        n16526) );
  OA22X1 U32447 ( .IN1(n18495), .IN2(n2560), .IN3(n18491), .IN4(n2525), .Q(
        n16527) );
  OA22X1 U32448 ( .IN1(n18484), .IN2(n2350), .IN3(n16440), .IN4(n2315), .Q(
        n16528) );
  OA22X1 U32449 ( .IN1(n18507), .IN2(n2699), .IN3(n16430), .IN4(n2664), .Q(
        n16518) );
  OA22X1 U32450 ( .IN1(n18495), .IN2(n2559), .IN3(n18492), .IN4(n2524), .Q(
        n16519) );
  OA22X1 U32451 ( .IN1(n18482), .IN2(n2349), .IN3(n16440), .IN4(n2314), .Q(
        n16520) );
  OA22X1 U32452 ( .IN1(n18508), .IN2(n2698), .IN3(n18504), .IN4(n2663), .Q(
        n16502) );
  OA22X1 U32453 ( .IN1(n18495), .IN2(n2558), .IN3(n18493), .IN4(n2523), .Q(
        n16503) );
  OA22X1 U32454 ( .IN1(n18484), .IN2(n2348), .IN3(n16440), .IN4(n2313), .Q(
        n16504) );
  OA22X1 U32455 ( .IN1(n18507), .IN2(n2697), .IN3(n16430), .IN4(n2662), .Q(
        n16494) );
  OA22X1 U32456 ( .IN1(n18494), .IN2(n2557), .IN3(n18492), .IN4(n2522), .Q(
        n16495) );
  OA22X1 U32457 ( .IN1(n18482), .IN2(n2347), .IN3(n16440), .IN4(n2312), .Q(
        n16496) );
  OA22X1 U32458 ( .IN1(n18458), .IN2(n2728), .IN3(n18455), .IN4(n2693), .Q(
        n16991) );
  OA22X1 U32459 ( .IN1(n18446), .IN2(n2588), .IN3(n16740), .IN4(n2553), .Q(
        n16992) );
  OA22X1 U32460 ( .IN1(n18436), .IN2(n2378), .IN3(n18431), .IN4(n2343), .Q(
        n16993) );
  OA22X1 U32461 ( .IN1(n18460), .IN2(n2727), .IN3(n16735), .IN4(n2692), .Q(
        n16903) );
  OA22X1 U32462 ( .IN1(n18448), .IN2(n2587), .IN3(n18444), .IN4(n2552), .Q(
        n16904) );
  OA22X1 U32463 ( .IN1(n18434), .IN2(n2377), .IN3(n16745), .IN4(n2342), .Q(
        n16905) );
  OA22X1 U32464 ( .IN1(n18458), .IN2(n2726), .IN3(n18456), .IN4(n2691), .Q(
        n16815) );
  OA22X1 U32465 ( .IN1(n18446), .IN2(n2586), .IN3(n18444), .IN4(n2551), .Q(
        n16816) );
  OA22X1 U32466 ( .IN1(n18436), .IN2(n2376), .IN3(n18432), .IN4(n2341), .Q(
        n16817) );
  OA22X1 U32467 ( .IN1(n18459), .IN2(n2725), .IN3(n18456), .IN4(n2690), .Q(
        n16791) );
  OA22X1 U32468 ( .IN1(n18448), .IN2(n2585), .IN3(n18444), .IN4(n2550), .Q(
        n16792) );
  OA22X1 U32469 ( .IN1(n18435), .IN2(n2375), .IN3(n16745), .IN4(n2340), .Q(
        n16793) );
  OA22X1 U32470 ( .IN1(n18460), .IN2(n2724), .IN3(n18456), .IN4(n2689), .Q(
        n16783) );
  OA22X1 U32471 ( .IN1(n18446), .IN2(n2584), .IN3(n18443), .IN4(n2549), .Q(
        n16784) );
  OA22X1 U32472 ( .IN1(n18434), .IN2(n2374), .IN3(n18432), .IN4(n2339), .Q(
        n16785) );
  OA22X1 U32473 ( .IN1(n18458), .IN2(n2723), .IN3(n18456), .IN4(n2688), .Q(
        n16775) );
  OA22X1 U32474 ( .IN1(n18447), .IN2(n2583), .IN3(n16740), .IN4(n2548), .Q(
        n16776) );
  OA22X1 U32475 ( .IN1(n18434), .IN2(n2373), .IN3(n16745), .IN4(n2338), .Q(
        n16777) );
  OA22X1 U32476 ( .IN1(n18460), .IN2(n2722), .IN3(n18456), .IN4(n2687), .Q(
        n16767) );
  OA22X1 U32477 ( .IN1(n18448), .IN2(n2582), .IN3(n18444), .IN4(n2547), .Q(
        n16768) );
  OA22X1 U32478 ( .IN1(n18436), .IN2(n2372), .IN3(n18432), .IN4(n2337), .Q(
        n16769) );
  OA22X1 U32479 ( .IN1(n18458), .IN2(n2721), .IN3(n18456), .IN4(n2686), .Q(
        n16759) );
  OA22X1 U32480 ( .IN1(n18448), .IN2(n2581), .IN3(n18444), .IN4(n2546), .Q(
        n16760) );
  OA22X1 U32481 ( .IN1(n18436), .IN2(n2371), .IN3(n18432), .IN4(n2336), .Q(
        n16761) );
  OA22X1 U32482 ( .IN1(n18459), .IN2(n2720), .IN3(n18456), .IN4(n2685), .Q(
        n16751) );
  OA22X1 U32483 ( .IN1(n18448), .IN2(n2580), .IN3(n18444), .IN4(n2545), .Q(
        n16752) );
  OA22X1 U32484 ( .IN1(n18436), .IN2(n2370), .IN3(n18432), .IN4(n2335), .Q(
        n16753) );
  OA22X1 U32485 ( .IN1(n18460), .IN2(n2719), .IN3(n18456), .IN4(n2684), .Q(
        n16733) );
  OA22X1 U32486 ( .IN1(n18448), .IN2(n2579), .IN3(n18444), .IN4(n2544), .Q(
        n16738) );
  OA22X1 U32487 ( .IN1(n18436), .IN2(n2369), .IN3(n18432), .IN4(n2334), .Q(
        n16743) );
  OA22X1 U32488 ( .IN1(n18458), .IN2(n2718), .IN3(n18455), .IN4(n2683), .Q(
        n16983) );
  OA22X1 U32489 ( .IN1(n18447), .IN2(n2578), .IN3(n16740), .IN4(n2543), .Q(
        n16984) );
  OA22X1 U32490 ( .IN1(n18434), .IN2(n2368), .IN3(n18431), .IN4(n2333), .Q(
        n16985) );
  OA22X1 U32491 ( .IN1(n18458), .IN2(n2717), .IN3(n18455), .IN4(n2682), .Q(
        n16975) );
  OA22X1 U32492 ( .IN1(n18446), .IN2(n2577), .IN3(n16740), .IN4(n2542), .Q(
        n16976) );
  OA22X1 U32493 ( .IN1(n18435), .IN2(n2367), .IN3(n18431), .IN4(n2332), .Q(
        n16977) );
  OA22X1 U32494 ( .IN1(n18458), .IN2(n2716), .IN3(n18455), .IN4(n2681), .Q(
        n16967) );
  OA22X1 U32495 ( .IN1(n18447), .IN2(n2576), .IN3(n16740), .IN4(n2541), .Q(
        n16968) );
  OA22X1 U32496 ( .IN1(n18436), .IN2(n2366), .IN3(n18431), .IN4(n2331), .Q(
        n16969) );
  OA22X1 U32497 ( .IN1(n18459), .IN2(n2715), .IN3(n18455), .IN4(n2680), .Q(
        n16959) );
  OA22X1 U32498 ( .IN1(n18446), .IN2(n2575), .IN3(n18443), .IN4(n2540), .Q(
        n16960) );
  OA22X1 U32499 ( .IN1(n18434), .IN2(n2365), .IN3(n16745), .IN4(n2330), .Q(
        n16961) );
  OA22X1 U32500 ( .IN1(n18459), .IN2(n2714), .IN3(n18455), .IN4(n2679), .Q(
        n16951) );
  OA22X1 U32501 ( .IN1(n18446), .IN2(n2574), .IN3(n18443), .IN4(n2539), .Q(
        n16952) );
  OA22X1 U32502 ( .IN1(n18434), .IN2(n2364), .IN3(n16745), .IN4(n2329), .Q(
        n16953) );
  OA22X1 U32503 ( .IN1(n18459), .IN2(n2713), .IN3(n16735), .IN4(n2678), .Q(
        n16943) );
  OA22X1 U32504 ( .IN1(n18446), .IN2(n2573), .IN3(n18443), .IN4(n2538), .Q(
        n16944) );
  OA22X1 U32505 ( .IN1(n18434), .IN2(n2363), .IN3(n16745), .IN4(n2328), .Q(
        n16945) );
  OA22X1 U32506 ( .IN1(n18459), .IN2(n2712), .IN3(n16735), .IN4(n2677), .Q(
        n16935) );
  OA22X1 U32507 ( .IN1(n18446), .IN2(n2572), .IN3(n18443), .IN4(n2537), .Q(
        n16936) );
  OA22X1 U32508 ( .IN1(n18434), .IN2(n2362), .IN3(n16745), .IN4(n2327), .Q(
        n16937) );
  OA22X1 U32509 ( .IN1(n18460), .IN2(n2711), .IN3(n16735), .IN4(n2676), .Q(
        n16927) );
  OA22X1 U32510 ( .IN1(n18447), .IN2(n2571), .IN3(n18443), .IN4(n2536), .Q(
        n16928) );
  OA22X1 U32511 ( .IN1(n18435), .IN2(n2361), .IN3(n18431), .IN4(n2326), .Q(
        n16929) );
  OA22X1 U32512 ( .IN1(n18460), .IN2(n2710), .IN3(n16735), .IN4(n2675), .Q(
        n16919) );
  OA22X1 U32513 ( .IN1(n18447), .IN2(n2570), .IN3(n18444), .IN4(n2535), .Q(
        n16920) );
  OA22X1 U32514 ( .IN1(n18434), .IN2(n2360), .IN3(n16745), .IN4(n2325), .Q(
        n16921) );
  OA22X1 U32515 ( .IN1(n18460), .IN2(n2709), .IN3(n16735), .IN4(n2674), .Q(
        n16911) );
  OA22X1 U32516 ( .IN1(n18446), .IN2(n2569), .IN3(n18444), .IN4(n2534), .Q(
        n16912) );
  OA22X1 U32517 ( .IN1(n18435), .IN2(n2359), .IN3(n16745), .IN4(n2324), .Q(
        n16913) );
  OA22X1 U32518 ( .IN1(n18459), .IN2(n2708), .IN3(n16735), .IN4(n2673), .Q(
        n16895) );
  OA22X1 U32519 ( .IN1(n18447), .IN2(n2568), .IN3(n16740), .IN4(n2533), .Q(
        n16896) );
  OA22X1 U32520 ( .IN1(n18435), .IN2(n2358), .IN3(n16745), .IN4(n2323), .Q(
        n16897) );
  OA22X1 U32521 ( .IN1(n18459), .IN2(n2707), .IN3(n18456), .IN4(n2672), .Q(
        n16887) );
  OA22X1 U32522 ( .IN1(n18447), .IN2(n2567), .IN3(n16740), .IN4(n2532), .Q(
        n16888) );
  OA22X1 U32523 ( .IN1(n18435), .IN2(n2357), .IN3(n18432), .IN4(n2322), .Q(
        n16889) );
  OA22X1 U32524 ( .IN1(n18459), .IN2(n2706), .IN3(n18455), .IN4(n2671), .Q(
        n16879) );
  OA22X1 U32525 ( .IN1(n18447), .IN2(n2566), .IN3(n16740), .IN4(n2531), .Q(
        n16880) );
  OA22X1 U32526 ( .IN1(n18434), .IN2(n2356), .IN3(n18431), .IN4(n2321), .Q(
        n16881) );
  OA22X1 U32527 ( .IN1(n18460), .IN2(n2705), .IN3(n16735), .IN4(n2670), .Q(
        n16871) );
  OA22X1 U32528 ( .IN1(n18447), .IN2(n2565), .IN3(n16740), .IN4(n2530), .Q(
        n16872) );
  OA22X1 U32529 ( .IN1(n18434), .IN2(n2355), .IN3(n16745), .IN4(n2320), .Q(
        n16873) );
  OA22X1 U32530 ( .IN1(n18458), .IN2(n2704), .IN3(n18455), .IN4(n2669), .Q(
        n16863) );
  OA22X1 U32531 ( .IN1(n18447), .IN2(n2564), .IN3(n18443), .IN4(n2529), .Q(
        n16864) );
  OA22X1 U32532 ( .IN1(n18435), .IN2(n2354), .IN3(n18431), .IN4(n2319), .Q(
        n16865) );
  OA22X1 U32533 ( .IN1(n18458), .IN2(n2703), .IN3(n18455), .IN4(n2668), .Q(
        n16855) );
  OA22X1 U32534 ( .IN1(n18448), .IN2(n2563), .IN3(n18443), .IN4(n2528), .Q(
        n16856) );
  OA22X1 U32535 ( .IN1(n18435), .IN2(n2353), .IN3(n18431), .IN4(n2318), .Q(
        n16857) );
  OA22X1 U32536 ( .IN1(n18458), .IN2(n2702), .IN3(n16735), .IN4(n2667), .Q(
        n16847) );
  OA22X1 U32537 ( .IN1(n18447), .IN2(n2562), .IN3(n16740), .IN4(n2527), .Q(
        n16848) );
  OA22X1 U32538 ( .IN1(n18435), .IN2(n2352), .IN3(n18432), .IN4(n2317), .Q(
        n16849) );
  OA22X1 U32539 ( .IN1(n18460), .IN2(n2701), .IN3(n18455), .IN4(n2666), .Q(
        n16839) );
  OA22X1 U32540 ( .IN1(n18446), .IN2(n2561), .IN3(n16740), .IN4(n2526), .Q(
        n16840) );
  OA22X1 U32541 ( .IN1(n18435), .IN2(n2351), .IN3(n18431), .IN4(n2316), .Q(
        n16841) );
  OA22X1 U32542 ( .IN1(n18459), .IN2(n2700), .IN3(n16735), .IN4(n2665), .Q(
        n16831) );
  OA22X1 U32543 ( .IN1(n18448), .IN2(n2560), .IN3(n16740), .IN4(n2525), .Q(
        n16832) );
  OA22X1 U32544 ( .IN1(n18436), .IN2(n2350), .IN3(n16745), .IN4(n2315), .Q(
        n16833) );
  OA22X1 U32545 ( .IN1(n18460), .IN2(n2699), .IN3(n16735), .IN4(n2664), .Q(
        n16823) );
  OA22X1 U32546 ( .IN1(n18446), .IN2(n2559), .IN3(n18443), .IN4(n2524), .Q(
        n16824) );
  OA22X1 U32547 ( .IN1(n18435), .IN2(n2349), .IN3(n16745), .IN4(n2314), .Q(
        n16825) );
  OA22X1 U32548 ( .IN1(n18458), .IN2(n2698), .IN3(n16735), .IN4(n2663), .Q(
        n16807) );
  OA22X1 U32549 ( .IN1(n18448), .IN2(n2558), .IN3(n18444), .IN4(n2523), .Q(
        n16808) );
  OA22X1 U32550 ( .IN1(n18436), .IN2(n2348), .IN3(n16745), .IN4(n2313), .Q(
        n16809) );
  OA22X1 U32551 ( .IN1(n18459), .IN2(n2697), .IN3(n18456), .IN4(n2662), .Q(
        n16799) );
  OA22X1 U32552 ( .IN1(n18448), .IN2(n2557), .IN3(n18443), .IN4(n2522), .Q(
        n16800) );
  OA22X1 U32553 ( .IN1(n18436), .IN2(n2347), .IN3(n18432), .IN4(n2312), .Q(
        n16801) );
  OA22X1 U32554 ( .IN1(n5111), .IN2(n2591), .IN3(n5407), .IN4(n2556), .Q(
        n14494) );
  OA22X1 U32555 ( .IN1(n5703), .IN2(n2521), .IN3(n5999), .IN4(n2486), .Q(
        n14495) );
  OA22X1 U32556 ( .IN1(n7959), .IN2(n2766), .IN3(n8255), .IN4(n2731), .Q(
        n14499) );
  OA22X1 U32557 ( .IN1(n5111), .IN2(n2590), .IN3(n5407), .IN4(n2555), .Q(
        n14504) );
  OA22X1 U32558 ( .IN1(n5703), .IN2(n2520), .IN3(n5999), .IN4(n2485), .Q(
        n14505) );
  OA22X1 U32559 ( .IN1(n7959), .IN2(n2765), .IN3(n8255), .IN4(n2730), .Q(
        n14508) );
  OA22X1 U32560 ( .IN1(n5111), .IN2(n2589), .IN3(n5407), .IN4(n2554), .Q(
        n14817) );
  OA22X1 U32561 ( .IN1(n5703), .IN2(n2519), .IN3(n5999), .IN4(n2484), .Q(
        n14836) );
  OA22X1 U32562 ( .IN1(n7959), .IN2(n2764), .IN3(n8255), .IN4(n2729), .Q(
        n14862) );
  OA22X1 U32563 ( .IN1(n5112), .IN2(n2591), .IN3(n5408), .IN4(n2556), .Q(
        n14879) );
  OA22X1 U32564 ( .IN1(n5704), .IN2(n2521), .IN3(n6000), .IN4(n2486), .Q(
        n14880) );
  OA22X1 U32565 ( .IN1(n7960), .IN2(n2766), .IN3(n8256), .IN4(n2731), .Q(
        n14883) );
  OA22X1 U32566 ( .IN1(n5112), .IN2(n2590), .IN3(n5408), .IN4(n2555), .Q(
        n14888) );
  OA22X1 U32567 ( .IN1(n5704), .IN2(n2520), .IN3(n6000), .IN4(n2485), .Q(
        n14889) );
  OA22X1 U32568 ( .IN1(n7960), .IN2(n2765), .IN3(n8256), .IN4(n2730), .Q(
        n14891) );
  OA22X1 U32569 ( .IN1(n5112), .IN2(n2589), .IN3(n5408), .IN4(n2554), .Q(
        n15168) );
  OA22X1 U32570 ( .IN1(n5704), .IN2(n2519), .IN3(n6000), .IN4(n2484), .Q(
        n15175) );
  OA22X1 U32571 ( .IN1(n7960), .IN2(n2764), .IN3(n8256), .IN4(n2729), .Q(
        n15179) );
  OA22X1 U32572 ( .IN1(n5113), .IN2(n2591), .IN3(n5409), .IN4(n2556), .Q(
        n15184) );
  OA22X1 U32573 ( .IN1(n5705), .IN2(n2521), .IN3(n6001), .IN4(n2486), .Q(
        n15185) );
  OA22X1 U32574 ( .IN1(n7961), .IN2(n2766), .IN3(n8257), .IN4(n2731), .Q(
        n15188) );
  OA22X1 U32575 ( .IN1(n5113), .IN2(n2590), .IN3(n5409), .IN4(n2555), .Q(
        n15193) );
  OA22X1 U32576 ( .IN1(n5705), .IN2(n2520), .IN3(n6001), .IN4(n2485), .Q(
        n15194) );
  OA22X1 U32577 ( .IN1(n7961), .IN2(n2765), .IN3(n8257), .IN4(n2730), .Q(
        n15196) );
  OA22X1 U32578 ( .IN1(n5113), .IN2(n2589), .IN3(n5409), .IN4(n2554), .Q(
        n15473) );
  OA22X1 U32579 ( .IN1(n5705), .IN2(n2519), .IN3(n6001), .IN4(n2484), .Q(
        n15480) );
  OA22X1 U32580 ( .IN1(n7961), .IN2(n2764), .IN3(n8257), .IN4(n2729), .Q(
        n15484) );
  OA22X1 U32581 ( .IN1(n5114), .IN2(n2591), .IN3(n5410), .IN4(n2556), .Q(
        n15489) );
  OA22X1 U32582 ( .IN1(n5706), .IN2(n2521), .IN3(n6002), .IN4(n2486), .Q(
        n15490) );
  OA22X1 U32583 ( .IN1(n7962), .IN2(n2766), .IN3(n8258), .IN4(n2731), .Q(
        n15493) );
  OA22X1 U32584 ( .IN1(n5114), .IN2(n2590), .IN3(n5410), .IN4(n2555), .Q(
        n15498) );
  OA22X1 U32585 ( .IN1(n5706), .IN2(n2520), .IN3(n6002), .IN4(n2485), .Q(
        n15499) );
  OA22X1 U32586 ( .IN1(n7962), .IN2(n2765), .IN3(n8258), .IN4(n2730), .Q(
        n15501) );
  OA22X1 U32587 ( .IN1(n5114), .IN2(n2589), .IN3(n5410), .IN4(n2554), .Q(
        n15778) );
  OA22X1 U32588 ( .IN1(n5706), .IN2(n2519), .IN3(n6002), .IN4(n2484), .Q(
        n15785) );
  OA22X1 U32589 ( .IN1(n7962), .IN2(n2764), .IN3(n8258), .IN4(n2729), .Q(
        n15789) );
  OA22X1 U32590 ( .IN1(n5115), .IN2(n2591), .IN3(n5411), .IN4(n2556), .Q(
        n15794) );
  OA22X1 U32591 ( .IN1(n5707), .IN2(n2521), .IN3(n6003), .IN4(n2486), .Q(
        n15795) );
  OA22X1 U32592 ( .IN1(n7963), .IN2(n2766), .IN3(n8259), .IN4(n2731), .Q(
        n15798) );
  OA22X1 U32593 ( .IN1(n5115), .IN2(n2590), .IN3(n5411), .IN4(n2555), .Q(
        n15803) );
  OA22X1 U32594 ( .IN1(n5707), .IN2(n2520), .IN3(n6003), .IN4(n2485), .Q(
        n15804) );
  OA22X1 U32595 ( .IN1(n7963), .IN2(n2765), .IN3(n8259), .IN4(n2730), .Q(
        n15806) );
  OA22X1 U32596 ( .IN1(n5115), .IN2(n2589), .IN3(n5411), .IN4(n2554), .Q(
        n16083) );
  OA22X1 U32597 ( .IN1(n5707), .IN2(n2519), .IN3(n6003), .IN4(n2484), .Q(
        n16090) );
  OA22X1 U32598 ( .IN1(n7963), .IN2(n2764), .IN3(n8259), .IN4(n2729), .Q(
        n16094) );
  OA22X1 U32599 ( .IN1(n5116), .IN2(n2591), .IN3(n5412), .IN4(n2556), .Q(
        n16099) );
  OA22X1 U32600 ( .IN1(n5708), .IN2(n2521), .IN3(n6004), .IN4(n2486), .Q(
        n16100) );
  OA22X1 U32601 ( .IN1(n7964), .IN2(n2766), .IN3(n8260), .IN4(n2731), .Q(
        n16103) );
  OA22X1 U32602 ( .IN1(n5116), .IN2(n2590), .IN3(n5412), .IN4(n2555), .Q(
        n16108) );
  OA22X1 U32603 ( .IN1(n5708), .IN2(n2520), .IN3(n6004), .IN4(n2485), .Q(
        n16109) );
  OA22X1 U32604 ( .IN1(n7964), .IN2(n2765), .IN3(n8260), .IN4(n2730), .Q(
        n16111) );
  OA22X1 U32605 ( .IN1(n5116), .IN2(n2589), .IN3(n5412), .IN4(n2554), .Q(
        n16388) );
  OA22X1 U32606 ( .IN1(n5708), .IN2(n2519), .IN3(n6004), .IN4(n2484), .Q(
        n16395) );
  OA22X1 U32607 ( .IN1(n7964), .IN2(n2764), .IN3(n8260), .IN4(n2729), .Q(
        n16399) );
  OA22X1 U32608 ( .IN1(n5117), .IN2(n2591), .IN3(n5413), .IN4(n2556), .Q(
        n16404) );
  OA22X1 U32609 ( .IN1(n5709), .IN2(n2521), .IN3(n6005), .IN4(n2486), .Q(
        n16405) );
  OA22X1 U32610 ( .IN1(n7965), .IN2(n2766), .IN3(n8261), .IN4(n2731), .Q(
        n16408) );
  OA22X1 U32611 ( .IN1(n5117), .IN2(n2590), .IN3(n5413), .IN4(n2555), .Q(
        n16413) );
  OA22X1 U32612 ( .IN1(n5709), .IN2(n2520), .IN3(n6005), .IN4(n2485), .Q(
        n16414) );
  OA22X1 U32613 ( .IN1(n7965), .IN2(n2765), .IN3(n8261), .IN4(n2730), .Q(
        n16416) );
  OA22X1 U32614 ( .IN1(n5117), .IN2(n2589), .IN3(n5413), .IN4(n2554), .Q(
        n16693) );
  OA22X1 U32615 ( .IN1(n5709), .IN2(n2519), .IN3(n6005), .IN4(n2484), .Q(
        n16700) );
  OA22X1 U32616 ( .IN1(n7965), .IN2(n2764), .IN3(n8261), .IN4(n2729), .Q(
        n16704) );
  OA22X1 U32617 ( .IN1(n5118), .IN2(n2591), .IN3(n5414), .IN4(n2556), .Q(
        n16709) );
  OA22X1 U32618 ( .IN1(n5710), .IN2(n2521), .IN3(n6006), .IN4(n2486), .Q(
        n16710) );
  OA22X1 U32619 ( .IN1(n7966), .IN2(n2766), .IN3(n8262), .IN4(n2731), .Q(
        n16713) );
  OA22X1 U32620 ( .IN1(n5118), .IN2(n2590), .IN3(n5414), .IN4(n2555), .Q(
        n16718) );
  OA22X1 U32621 ( .IN1(n5710), .IN2(n2520), .IN3(n6006), .IN4(n2485), .Q(
        n16719) );
  OA22X1 U32622 ( .IN1(n7966), .IN2(n2765), .IN3(n8262), .IN4(n2730), .Q(
        n16721) );
  OA22X1 U32623 ( .IN1(n5118), .IN2(n2589), .IN3(n5414), .IN4(n2554), .Q(
        n16998) );
  OA22X1 U32624 ( .IN1(n5710), .IN2(n2519), .IN3(n6006), .IN4(n2484), .Q(
        n17033) );
  OA22X1 U32625 ( .IN1(n7966), .IN2(n2764), .IN3(n8262), .IN4(n2729), .Q(
        n17127) );
  INVX0 U32626 ( .IN(n14824), .QN(n3851) );
  INVX0 U32627 ( .IN(n14819), .QN(n3806) );
  INVX0 U32628 ( .IN(n14857), .QN(n4166) );
  INVX0 U32629 ( .IN(n14842), .QN(n3761) );
  INVX0 U32630 ( .IN(n14838), .QN(n3716) );
  INVX0 U32631 ( .IN(n14854), .QN(n4121) );
  INVX0 U32632 ( .IN(n14867), .QN(n4076) );
  INVX0 U32633 ( .IN(n14845), .QN(n3671) );
  INVX0 U32634 ( .IN(n14849), .QN(n3626) );
  INVX0 U32635 ( .IN(n14864), .QN(n4031) );
  INVX0 U32636 ( .IN(n14870), .QN(n3986) );
  INVX0 U32637 ( .IN(n14860), .QN(n3581) );
  INVX0 U32638 ( .IN(n14873), .QN(n3536) );
  INVX0 U32639 ( .IN(n14833), .QN(n3896) );
  INVX0 U32640 ( .IN(n14828), .QN(n3941) );
  INVX0 U32641 ( .IN(n14825), .QN(n3850) );
  INVX0 U32642 ( .IN(n14820), .QN(n3805) );
  INVX0 U32643 ( .IN(n14858), .QN(n4165) );
  INVX0 U32644 ( .IN(n14843), .QN(n3760) );
  INVX0 U32645 ( .IN(n14839), .QN(n3715) );
  INVX0 U32646 ( .IN(n14855), .QN(n4120) );
  INVX0 U32647 ( .IN(n14868), .QN(n4075) );
  INVX0 U32648 ( .IN(n14846), .QN(n3670) );
  INVX0 U32649 ( .IN(n14850), .QN(n3625) );
  INVX0 U32650 ( .IN(n14865), .QN(n4030) );
  INVX0 U32651 ( .IN(n14871), .QN(n3985) );
  INVX0 U32652 ( .IN(n14861), .QN(n3580) );
  INVX0 U32653 ( .IN(n14874), .QN(n3535) );
  INVX0 U32654 ( .IN(n14834), .QN(n3895) );
  INVX0 U32655 ( .IN(n14829), .QN(n3940) );
  INVX0 U32656 ( .IN(n14823), .QN(n3845) );
  INVX0 U32657 ( .IN(n14818), .QN(n3800) );
  INVX0 U32658 ( .IN(n14856), .QN(n4160) );
  INVX0 U32659 ( .IN(n14841), .QN(n3755) );
  INVX0 U32660 ( .IN(n14837), .QN(n3710) );
  INVX0 U32661 ( .IN(n14853), .QN(n4115) );
  INVX0 U32662 ( .IN(n14866), .QN(n4070) );
  INVX0 U32663 ( .IN(n14844), .QN(n3665) );
  INVX0 U32664 ( .IN(n14848), .QN(n3620) );
  INVX0 U32665 ( .IN(n14863), .QN(n4025) );
  INVX0 U32666 ( .IN(n14869), .QN(n3980) );
  INVX0 U32667 ( .IN(n14859), .QN(n3575) );
  INVX0 U32668 ( .IN(n14872), .QN(n3530) );
  INVX0 U32669 ( .IN(n14832), .QN(n3890) );
  INVX0 U32670 ( .IN(n14827), .QN(n3935) );
  INVX0 U32671 ( .IN(n13677), .QN(n3430) );
  INVX0 U32672 ( .IN(n13368), .QN(n3434) );
  INVX0 U32673 ( .IN(n11202), .QN(n3402) );
  INVX0 U32674 ( .IN(n13059), .QN(n3438) );
  INVX0 U32675 ( .IN(n12750), .QN(n3442) );
  INVX0 U32676 ( .IN(n10893), .QN(n3406) );
  INVX0 U32677 ( .IN(n10583), .QN(n3410) );
  INVX0 U32678 ( .IN(n12441), .QN(n3446) );
  INVX0 U32679 ( .IN(n12132), .QN(n3450) );
  INVX0 U32680 ( .IN(n10274), .QN(n3414) );
  INVX0 U32681 ( .IN(n9964), .QN(n3418) );
  INVX0 U32682 ( .IN(n11822), .QN(n3454) );
  INVX0 U32683 ( .IN(n11512), .QN(n3458) );
  INVX0 U32684 ( .IN(n9654), .QN(n3422) );
  INVX0 U32685 ( .IN(n9343), .QN(n3426) );
  OA21X1 U32686 ( .IN1(n13916), .IN2(n3146), .IN3(n13903), .Q(n13897) );
  OA21X1 U32687 ( .IN1(n13849), .IN2(n13835), .IN3(n13837), .Q(n13829) );
  OA21X1 U32688 ( .IN1(n13719), .IN2(n13675), .IN3(n13709), .Q(n13703) );
  OA21X1 U32689 ( .IN1(n13607), .IN2(n3152), .IN3(n13594), .Q(n13588) );
  OA21X1 U32690 ( .IN1(n13540), .IN2(n13526), .IN3(n13528), .Q(n13520) );
  OA21X1 U32691 ( .IN1(n13410), .IN2(n13366), .IN3(n13400), .Q(n13394) );
  OA21X1 U32692 ( .IN1(n11441), .IN2(n3104), .IN3(n11428), .Q(n11422) );
  OA21X1 U32693 ( .IN1(n11374), .IN2(n11360), .IN3(n11362), .Q(n11354) );
  OA21X1 U32694 ( .IN1(n11244), .IN2(n11200), .IN3(n11234), .Q(n11228) );
  OA21X1 U32695 ( .IN1(n13298), .IN2(n3158), .IN3(n13285), .Q(n13279) );
  OA21X1 U32696 ( .IN1(n13231), .IN2(n13217), .IN3(n13219), .Q(n13211) );
  OA21X1 U32697 ( .IN1(n13101), .IN2(n13057), .IN3(n13091), .Q(n13085) );
  OA21X1 U32698 ( .IN1(n12989), .IN2(n3164), .IN3(n12976), .Q(n12970) );
  OA21X1 U32699 ( .IN1(n12922), .IN2(n12908), .IN3(n12910), .Q(n12902) );
  OA21X1 U32700 ( .IN1(n12792), .IN2(n12748), .IN3(n12782), .Q(n12776) );
  OA21X1 U32701 ( .IN1(n11132), .IN2(n3110), .IN3(n11119), .Q(n11113) );
  OA21X1 U32702 ( .IN1(n11065), .IN2(n11051), .IN3(n11053), .Q(n11045) );
  OA21X1 U32703 ( .IN1(n10935), .IN2(n10891), .IN3(n10925), .Q(n10919) );
  OA21X1 U32704 ( .IN1(n10822), .IN2(n3116), .IN3(n10809), .Q(n10803) );
  OA21X1 U32705 ( .IN1(n10755), .IN2(n10741), .IN3(n10743), .Q(n10735) );
  OA21X1 U32706 ( .IN1(n10625), .IN2(n10581), .IN3(n10615), .Q(n10609) );
  OA21X1 U32707 ( .IN1(n12680), .IN2(n3170), .IN3(n12667), .Q(n12661) );
  OA21X1 U32708 ( .IN1(n12613), .IN2(n12599), .IN3(n12601), .Q(n12593) );
  OA21X1 U32709 ( .IN1(n12483), .IN2(n12439), .IN3(n12473), .Q(n12467) );
  OA21X1 U32710 ( .IN1(n12371), .IN2(n3176), .IN3(n12358), .Q(n12352) );
  OA21X1 U32711 ( .IN1(n12304), .IN2(n12290), .IN3(n12292), .Q(n12284) );
  OA21X1 U32712 ( .IN1(n12174), .IN2(n12130), .IN3(n12164), .Q(n12158) );
  OA21X1 U32713 ( .IN1(n10513), .IN2(n3122), .IN3(n10500), .Q(n10494) );
  OA21X1 U32714 ( .IN1(n10446), .IN2(n10432), .IN3(n10434), .Q(n10426) );
  OA21X1 U32715 ( .IN1(n10316), .IN2(n10272), .IN3(n10306), .Q(n10300) );
  OA21X1 U32716 ( .IN1(n10203), .IN2(n3128), .IN3(n10190), .Q(n10184) );
  OA21X1 U32717 ( .IN1(n10136), .IN2(n10122), .IN3(n10124), .Q(n10116) );
  OA21X1 U32718 ( .IN1(n10006), .IN2(n9962), .IN3(n9996), .Q(n9990) );
  OA21X1 U32719 ( .IN1(n12061), .IN2(n3182), .IN3(n12048), .Q(n12042) );
  OA21X1 U32720 ( .IN1(n11994), .IN2(n11980), .IN3(n11982), .Q(n11974) );
  OA21X1 U32721 ( .IN1(n11864), .IN2(n11820), .IN3(n11854), .Q(n11848) );
  OA21X1 U32722 ( .IN1(n11751), .IN2(n3188), .IN3(n11738), .Q(n11732) );
  OA21X1 U32723 ( .IN1(n11684), .IN2(n11670), .IN3(n11672), .Q(n11664) );
  OA21X1 U32724 ( .IN1(n11554), .IN2(n11510), .IN3(n11544), .Q(n11538) );
  OA21X1 U32725 ( .IN1(n9893), .IN2(n3134), .IN3(n9880), .Q(n9874) );
  OA21X1 U32726 ( .IN1(n9826), .IN2(n9812), .IN3(n9814), .Q(n9806) );
  OA21X1 U32727 ( .IN1(n9696), .IN2(n9652), .IN3(n9686), .Q(n9680) );
  OA21X1 U32728 ( .IN1(n9582), .IN2(n3140), .IN3(n9569), .Q(n9563) );
  OA21X1 U32729 ( .IN1(n9515), .IN2(n9501), .IN3(n9503), .Q(n9495) );
  OA21X1 U32730 ( .IN1(n9385), .IN2(n9341), .IN3(n9375), .Q(n9369) );
  OA21X1 U32731 ( .IN1(n13982), .IN2(n13968), .IN3(n13970), .Q(n13962) );
  OA21X1 U32732 ( .IN1(n14190), .IN2(n3094), .IN3(n14177), .Q(n14171) );
  OA21X1 U32733 ( .IN1(n14122), .IN2(n14108), .IN3(n14110), .Q(n14102) );
  OA21X1 U32734 ( .IN1(n13818), .IN2(n13846), .IN3(n13816), .Q(n13819) );
  OA21X1 U32735 ( .IN1(n13832), .IN2(n13829), .IN3(n13834), .Q(n13846) );
  OA21X1 U32736 ( .IN1(n13674), .IN2(n13717), .IN3(n13691), .Q(n13693) );
  OA21X1 U32737 ( .IN1(n13673), .IN2(n13703), .IN3(n13707), .Q(n13717) );
  OA21X1 U32738 ( .IN1(n13509), .IN2(n13537), .IN3(n13507), .Q(n13510) );
  OA21X1 U32739 ( .IN1(n13523), .IN2(n13520), .IN3(n13525), .Q(n13537) );
  OA21X1 U32740 ( .IN1(n13365), .IN2(n13408), .IN3(n13382), .Q(n13384) );
  OA21X1 U32741 ( .IN1(n13364), .IN2(n13394), .IN3(n13398), .Q(n13408) );
  OA21X1 U32742 ( .IN1(n11343), .IN2(n11371), .IN3(n11341), .Q(n11344) );
  OA21X1 U32743 ( .IN1(n11357), .IN2(n11354), .IN3(n11359), .Q(n11371) );
  OA21X1 U32744 ( .IN1(n11199), .IN2(n11242), .IN3(n11216), .Q(n11218) );
  OA21X1 U32745 ( .IN1(n11198), .IN2(n11228), .IN3(n11232), .Q(n11242) );
  OA21X1 U32746 ( .IN1(n13200), .IN2(n13228), .IN3(n13198), .Q(n13201) );
  OA21X1 U32747 ( .IN1(n13214), .IN2(n13211), .IN3(n13216), .Q(n13228) );
  OA21X1 U32748 ( .IN1(n13056), .IN2(n13099), .IN3(n13073), .Q(n13075) );
  OA21X1 U32749 ( .IN1(n13055), .IN2(n13085), .IN3(n13089), .Q(n13099) );
  OA21X1 U32750 ( .IN1(n12891), .IN2(n12919), .IN3(n12889), .Q(n12892) );
  OA21X1 U32751 ( .IN1(n12905), .IN2(n12902), .IN3(n12907), .Q(n12919) );
  OA21X1 U32752 ( .IN1(n12747), .IN2(n12790), .IN3(n12764), .Q(n12766) );
  OA21X1 U32753 ( .IN1(n12746), .IN2(n12776), .IN3(n12780), .Q(n12790) );
  OA21X1 U32754 ( .IN1(n11034), .IN2(n11062), .IN3(n11032), .Q(n11035) );
  OA21X1 U32755 ( .IN1(n11048), .IN2(n11045), .IN3(n11050), .Q(n11062) );
  OA21X1 U32756 ( .IN1(n10890), .IN2(n10933), .IN3(n10907), .Q(n10909) );
  OA21X1 U32757 ( .IN1(n10889), .IN2(n10919), .IN3(n10923), .Q(n10933) );
  OA21X1 U32758 ( .IN1(n10724), .IN2(n10752), .IN3(n10722), .Q(n10725) );
  OA21X1 U32759 ( .IN1(n10738), .IN2(n10735), .IN3(n10740), .Q(n10752) );
  OA21X1 U32760 ( .IN1(n10580), .IN2(n10623), .IN3(n10597), .Q(n10599) );
  OA21X1 U32761 ( .IN1(n10579), .IN2(n10609), .IN3(n10613), .Q(n10623) );
  OA21X1 U32762 ( .IN1(n12582), .IN2(n12610), .IN3(n12580), .Q(n12583) );
  OA21X1 U32763 ( .IN1(n12596), .IN2(n12593), .IN3(n12598), .Q(n12610) );
  OA21X1 U32764 ( .IN1(n12438), .IN2(n12481), .IN3(n12455), .Q(n12457) );
  OA21X1 U32765 ( .IN1(n12437), .IN2(n12467), .IN3(n12471), .Q(n12481) );
  OA21X1 U32766 ( .IN1(n12273), .IN2(n12301), .IN3(n12271), .Q(n12274) );
  OA21X1 U32767 ( .IN1(n12287), .IN2(n12284), .IN3(n12289), .Q(n12301) );
  OA21X1 U32768 ( .IN1(n12129), .IN2(n12172), .IN3(n12146), .Q(n12148) );
  OA21X1 U32769 ( .IN1(n12128), .IN2(n12158), .IN3(n12162), .Q(n12172) );
  OA21X1 U32770 ( .IN1(n10415), .IN2(n10443), .IN3(n10413), .Q(n10416) );
  OA21X1 U32771 ( .IN1(n10429), .IN2(n10426), .IN3(n10431), .Q(n10443) );
  OA21X1 U32772 ( .IN1(n10271), .IN2(n10314), .IN3(n10288), .Q(n10290) );
  OA21X1 U32773 ( .IN1(n10270), .IN2(n10300), .IN3(n10304), .Q(n10314) );
  OA21X1 U32774 ( .IN1(n10105), .IN2(n10133), .IN3(n10103), .Q(n10106) );
  OA21X1 U32775 ( .IN1(n10119), .IN2(n10116), .IN3(n10121), .Q(n10133) );
  OA21X1 U32776 ( .IN1(n9961), .IN2(n10004), .IN3(n9978), .Q(n9980) );
  OA21X1 U32777 ( .IN1(n9960), .IN2(n9990), .IN3(n9994), .Q(n10004) );
  OA21X1 U32778 ( .IN1(n11963), .IN2(n11991), .IN3(n11961), .Q(n11964) );
  OA21X1 U32779 ( .IN1(n11977), .IN2(n11974), .IN3(n11979), .Q(n11991) );
  OA21X1 U32780 ( .IN1(n11819), .IN2(n11862), .IN3(n11836), .Q(n11838) );
  OA21X1 U32781 ( .IN1(n11818), .IN2(n11848), .IN3(n11852), .Q(n11862) );
  OA21X1 U32782 ( .IN1(n11653), .IN2(n11681), .IN3(n11651), .Q(n11654) );
  OA21X1 U32783 ( .IN1(n11667), .IN2(n11664), .IN3(n11669), .Q(n11681) );
  OA21X1 U32784 ( .IN1(n11509), .IN2(n11552), .IN3(n11526), .Q(n11528) );
  OA21X1 U32785 ( .IN1(n11508), .IN2(n11538), .IN3(n11542), .Q(n11552) );
  OA21X1 U32786 ( .IN1(n9795), .IN2(n9823), .IN3(n9793), .Q(n9796) );
  OA21X1 U32787 ( .IN1(n9809), .IN2(n9806), .IN3(n9811), .Q(n9823) );
  OA21X1 U32788 ( .IN1(n9651), .IN2(n9694), .IN3(n9668), .Q(n9670) );
  OA21X1 U32789 ( .IN1(n9650), .IN2(n9680), .IN3(n9684), .Q(n9694) );
  OA21X1 U32790 ( .IN1(n9484), .IN2(n9512), .IN3(n9482), .Q(n9485) );
  OA21X1 U32791 ( .IN1(n9498), .IN2(n9495), .IN3(n9500), .Q(n9512) );
  OA21X1 U32792 ( .IN1(n9340), .IN2(n9383), .IN3(n9357), .Q(n9359) );
  OA21X1 U32793 ( .IN1(n9339), .IN2(n9369), .IN3(n9373), .Q(n9383) );
  OA21X1 U32794 ( .IN1(n13950), .IN2(n13979), .IN3(n13948), .Q(n13951) );
  OA21X1 U32795 ( .IN1(n13965), .IN2(n13962), .IN3(n13967), .Q(n13979) );
  OA21X1 U32796 ( .IN1(n14090), .IN2(n14119), .IN3(n14088), .Q(n14091) );
  OA21X1 U32797 ( .IN1(n14105), .IN2(n14102), .IN3(n14107), .Q(n14119) );
  NOR2X0 U32798 ( .IN1(n14101), .IN2(n14105), .QN(n14086) );
  NOR2X0 U32799 ( .IN1(n13702), .IN2(n13673), .QN(n13689) );
  NOR2X0 U32800 ( .IN1(n13393), .IN2(n13364), .QN(n13380) );
  NOR2X0 U32801 ( .IN1(n11227), .IN2(n11198), .QN(n11214) );
  NOR2X0 U32802 ( .IN1(n13084), .IN2(n13055), .QN(n13071) );
  NOR2X0 U32803 ( .IN1(n12775), .IN2(n12746), .QN(n12762) );
  NOR2X0 U32804 ( .IN1(n10918), .IN2(n10889), .QN(n10905) );
  NOR2X0 U32805 ( .IN1(n10608), .IN2(n10579), .QN(n10595) );
  NOR2X0 U32806 ( .IN1(n12466), .IN2(n12437), .QN(n12453) );
  NOR2X0 U32807 ( .IN1(n12157), .IN2(n12128), .QN(n12144) );
  NOR2X0 U32808 ( .IN1(n10299), .IN2(n10270), .QN(n10286) );
  NOR2X0 U32809 ( .IN1(n9989), .IN2(n9960), .QN(n9976) );
  NOR2X0 U32810 ( .IN1(n11847), .IN2(n11818), .QN(n11834) );
  NOR2X0 U32811 ( .IN1(n11537), .IN2(n11508), .QN(n11524) );
  NOR2X0 U32812 ( .IN1(n9679), .IN2(n9650), .QN(n9666) );
  NOR2X0 U32813 ( .IN1(n9368), .IN2(n9339), .QN(n9355) );
  NOR2X0 U32814 ( .IN1(n13961), .IN2(n13965), .QN(n13946) );
  NOR2X0 U32815 ( .IN1(n13765), .IN2(n13769), .QN(n13756) );
  NOR2X0 U32816 ( .IN1(n13456), .IN2(n13460), .QN(n13447) );
  NOR2X0 U32817 ( .IN1(n11290), .IN2(n11294), .QN(n11281) );
  NOR2X0 U32818 ( .IN1(n13147), .IN2(n13151), .QN(n13138) );
  NOR2X0 U32819 ( .IN1(n12838), .IN2(n12842), .QN(n12829) );
  NOR2X0 U32820 ( .IN1(n10981), .IN2(n10985), .QN(n10972) );
  NOR2X0 U32821 ( .IN1(n10671), .IN2(n10675), .QN(n10662) );
  NOR2X0 U32822 ( .IN1(n12529), .IN2(n12533), .QN(n12520) );
  NOR2X0 U32823 ( .IN1(n12220), .IN2(n12224), .QN(n12211) );
  NOR2X0 U32824 ( .IN1(n10362), .IN2(n10366), .QN(n10353) );
  NOR2X0 U32825 ( .IN1(n10052), .IN2(n10056), .QN(n10043) );
  NOR2X0 U32826 ( .IN1(n11910), .IN2(n11914), .QN(n11901) );
  NOR2X0 U32827 ( .IN1(n11600), .IN2(n11604), .QN(n11591) );
  NOR2X0 U32828 ( .IN1(n9742), .IN2(n9746), .QN(n9733) );
  NOR2X0 U32829 ( .IN1(n9431), .IN2(n9435), .QN(n9422) );
  NOR2X0 U32830 ( .IN1(n14029), .IN2(n14033), .QN(n14020) );
  NOR2X0 U32831 ( .IN1(n13828), .IN2(n13832), .QN(n13814) );
  NOR2X0 U32832 ( .IN1(n13519), .IN2(n13523), .QN(n13505) );
  NOR2X0 U32833 ( .IN1(n11353), .IN2(n11357), .QN(n11339) );
  NOR2X0 U32834 ( .IN1(n13210), .IN2(n13214), .QN(n13196) );
  NOR2X0 U32835 ( .IN1(n12901), .IN2(n12905), .QN(n12887) );
  NOR2X0 U32836 ( .IN1(n11044), .IN2(n11048), .QN(n11030) );
  NOR2X0 U32837 ( .IN1(n10734), .IN2(n10738), .QN(n10720) );
  NOR2X0 U32838 ( .IN1(n12592), .IN2(n12596), .QN(n12578) );
  NOR2X0 U32839 ( .IN1(n12283), .IN2(n12287), .QN(n12269) );
  NOR2X0 U32840 ( .IN1(n10425), .IN2(n10429), .QN(n10411) );
  NOR2X0 U32841 ( .IN1(n10115), .IN2(n10119), .QN(n10101) );
  NOR2X0 U32842 ( .IN1(n11973), .IN2(n11977), .QN(n11959) );
  NOR2X0 U32843 ( .IN1(n11663), .IN2(n11667), .QN(n11649) );
  NOR2X0 U32844 ( .IN1(n9805), .IN2(n9809), .QN(n9791) );
  NOR2X0 U32845 ( .IN1(n9494), .IN2(n9498), .QN(n9480) );
  AND3X1 U32846 ( .IN1(n13815), .IN2(n13816), .IN3(n13809), .Q(n13810) );
  OR2X1 U32847 ( .IN1(n13817), .IN2(n13818), .Q(n13815) );
  AND3X1 U32848 ( .IN1(n13690), .IN2(n13691), .IN3(n13684), .Q(n13685) );
  OR2X1 U32849 ( .IN1(n13692), .IN2(n13674), .Q(n13690) );
  AND3X1 U32850 ( .IN1(n13506), .IN2(n13507), .IN3(n13500), .Q(n13501) );
  OR2X1 U32851 ( .IN1(n13508), .IN2(n13509), .Q(n13506) );
  AND3X1 U32852 ( .IN1(n13381), .IN2(n13382), .IN3(n13375), .Q(n13376) );
  OR2X1 U32853 ( .IN1(n13383), .IN2(n13365), .Q(n13381) );
  AND3X1 U32854 ( .IN1(n11340), .IN2(n11341), .IN3(n11334), .Q(n11335) );
  OR2X1 U32855 ( .IN1(n11342), .IN2(n11343), .Q(n11340) );
  AND3X1 U32856 ( .IN1(n11215), .IN2(n11216), .IN3(n11209), .Q(n11210) );
  OR2X1 U32857 ( .IN1(n11217), .IN2(n11199), .Q(n11215) );
  AND3X1 U32858 ( .IN1(n13072), .IN2(n13073), .IN3(n13066), .Q(n13067) );
  OR2X1 U32859 ( .IN1(n13074), .IN2(n13056), .Q(n13072) );
  AND3X1 U32860 ( .IN1(n12763), .IN2(n12764), .IN3(n12757), .Q(n12758) );
  OR2X1 U32861 ( .IN1(n12765), .IN2(n12747), .Q(n12763) );
  AND3X1 U32862 ( .IN1(n10906), .IN2(n10907), .IN3(n10900), .Q(n10901) );
  OR2X1 U32863 ( .IN1(n10908), .IN2(n10890), .Q(n10906) );
  AND3X1 U32864 ( .IN1(n10596), .IN2(n10597), .IN3(n10590), .Q(n10591) );
  OR2X1 U32865 ( .IN1(n10598), .IN2(n10580), .Q(n10596) );
  AND3X1 U32866 ( .IN1(n12579), .IN2(n12580), .IN3(n12573), .Q(n12574) );
  OR2X1 U32867 ( .IN1(n12581), .IN2(n12582), .Q(n12579) );
  AND3X1 U32868 ( .IN1(n12454), .IN2(n12455), .IN3(n12448), .Q(n12449) );
  OR2X1 U32869 ( .IN1(n12456), .IN2(n12438), .Q(n12454) );
  AND3X1 U32870 ( .IN1(n12270), .IN2(n12271), .IN3(n12264), .Q(n12265) );
  OR2X1 U32871 ( .IN1(n12272), .IN2(n12273), .Q(n12270) );
  AND3X1 U32872 ( .IN1(n12145), .IN2(n12146), .IN3(n12139), .Q(n12140) );
  OR2X1 U32873 ( .IN1(n12147), .IN2(n12129), .Q(n12145) );
  AND3X1 U32874 ( .IN1(n10287), .IN2(n10288), .IN3(n10281), .Q(n10282) );
  OR2X1 U32875 ( .IN1(n10289), .IN2(n10271), .Q(n10287) );
  AND3X1 U32876 ( .IN1(n9977), .IN2(n9978), .IN3(n9971), .Q(n9972) );
  OR2X1 U32877 ( .IN1(n9979), .IN2(n9961), .Q(n9977) );
  AND3X1 U32878 ( .IN1(n11835), .IN2(n11836), .IN3(n11829), .Q(n11830) );
  OR2X1 U32879 ( .IN1(n11837), .IN2(n11819), .Q(n11835) );
  AND3X1 U32880 ( .IN1(n11525), .IN2(n11526), .IN3(n11519), .Q(n11520) );
  OR2X1 U32881 ( .IN1(n11527), .IN2(n11509), .Q(n11525) );
  AND3X1 U32882 ( .IN1(n9792), .IN2(n9793), .IN3(n9786), .Q(n9787) );
  OR2X1 U32883 ( .IN1(n9794), .IN2(n9795), .Q(n9792) );
  AND3X1 U32884 ( .IN1(n9667), .IN2(n9668), .IN3(n9661), .Q(n9662) );
  OR2X1 U32885 ( .IN1(n9669), .IN2(n9651), .Q(n9667) );
  AND3X1 U32886 ( .IN1(n9481), .IN2(n9482), .IN3(n9475), .Q(n9476) );
  OR2X1 U32887 ( .IN1(n9483), .IN2(n9484), .Q(n9481) );
  AND3X1 U32888 ( .IN1(n9356), .IN2(n9357), .IN3(n9350), .Q(n9351) );
  OR2X1 U32889 ( .IN1(n9358), .IN2(n9340), .Q(n9356) );
  AND3X1 U32890 ( .IN1(n13947), .IN2(n13948), .IN3(n13940), .Q(n13941) );
  OR2X1 U32891 ( .IN1(n13949), .IN2(n13950), .Q(n13947) );
  AND3X1 U32892 ( .IN1(n14087), .IN2(n14088), .IN3(n14081), .Q(n14082) );
  OR2X1 U32893 ( .IN1(n14089), .IN2(n14090), .Q(n14087) );
  AND3X1 U32894 ( .IN1(n13884), .IN2(n13885), .IN3(n13875), .Q(n13882) );
  OR2X1 U32895 ( .IN1(n13886), .IN2(n3323), .Q(n13884) );
  AND3X1 U32896 ( .IN1(n13575), .IN2(n13576), .IN3(n13566), .Q(n13573) );
  OR2X1 U32897 ( .IN1(n13577), .IN2(n3331), .Q(n13575) );
  AND3X1 U32898 ( .IN1(n11409), .IN2(n11410), .IN3(n11400), .Q(n11407) );
  OR2X1 U32899 ( .IN1(n11411), .IN2(n3267), .Q(n11409) );
  AND3X1 U32900 ( .IN1(n13266), .IN2(n13267), .IN3(n13257), .Q(n13264) );
  OR2X1 U32901 ( .IN1(n13268), .IN2(n3339), .Q(n13266) );
  AND3X1 U32902 ( .IN1(n12957), .IN2(n12958), .IN3(n12948), .Q(n12955) );
  OR2X1 U32903 ( .IN1(n12959), .IN2(n3347), .Q(n12957) );
  AND3X1 U32904 ( .IN1(n11100), .IN2(n11101), .IN3(n11091), .Q(n11098) );
  OR2X1 U32905 ( .IN1(n11102), .IN2(n3275), .Q(n11100) );
  AND3X1 U32906 ( .IN1(n10967), .IN2(n10968), .IN3(n10960), .Q(n10966) );
  OR2X1 U32907 ( .IN1(n10969), .IN2(n10970), .Q(n10967) );
  AND3X1 U32908 ( .IN1(n10790), .IN2(n10791), .IN3(n10781), .Q(n10788) );
  OR2X1 U32909 ( .IN1(n10792), .IN2(n3283), .Q(n10790) );
  AND3X1 U32910 ( .IN1(n12648), .IN2(n12649), .IN3(n12639), .Q(n12646) );
  OR2X1 U32911 ( .IN1(n12650), .IN2(n3355), .Q(n12648) );
  AND3X1 U32912 ( .IN1(n12339), .IN2(n12340), .IN3(n12330), .Q(n12337) );
  OR2X1 U32913 ( .IN1(n12341), .IN2(n3363), .Q(n12339) );
  AND3X1 U32914 ( .IN1(n10481), .IN2(n10482), .IN3(n10472), .Q(n10479) );
  OR2X1 U32915 ( .IN1(n10483), .IN2(n3291), .Q(n10481) );
  AND3X1 U32916 ( .IN1(n10348), .IN2(n10349), .IN3(n10341), .Q(n10347) );
  OR2X1 U32917 ( .IN1(n10350), .IN2(n10351), .Q(n10348) );
  AND3X1 U32918 ( .IN1(n10171), .IN2(n10172), .IN3(n10162), .Q(n10169) );
  OR2X1 U32919 ( .IN1(n10173), .IN2(n3299), .Q(n10171) );
  AND3X1 U32920 ( .IN1(n12029), .IN2(n12030), .IN3(n12020), .Q(n12027) );
  OR2X1 U32921 ( .IN1(n12031), .IN2(n3371), .Q(n12029) );
  AND3X1 U32922 ( .IN1(n11719), .IN2(n11720), .IN3(n11710), .Q(n11717) );
  OR2X1 U32923 ( .IN1(n11721), .IN2(n3379), .Q(n11719) );
  AND3X1 U32924 ( .IN1(n9861), .IN2(n9862), .IN3(n9852), .Q(n9859) );
  OR2X1 U32925 ( .IN1(n9863), .IN2(n3307), .Q(n9861) );
  AND3X1 U32926 ( .IN1(n9728), .IN2(n9729), .IN3(n9721), .Q(n9727) );
  OR2X1 U32927 ( .IN1(n9730), .IN2(n9731), .Q(n9728) );
  AND3X1 U32928 ( .IN1(n9550), .IN2(n9551), .IN3(n9541), .Q(n9548) );
  OR2X1 U32929 ( .IN1(n9552), .IN2(n3315), .Q(n9550) );
  AND3X1 U32930 ( .IN1(n14158), .IN2(n14159), .IN3(n14149), .Q(n14156) );
  OR2X1 U32931 ( .IN1(n14160), .IN2(n3255), .Q(n14158) );
  AND3X1 U32932 ( .IN1(n13751), .IN2(n13752), .IN3(n13744), .Q(n13750) );
  OR2X1 U32933 ( .IN1(n13753), .IN2(n13754), .Q(n13751) );
  AND3X1 U32934 ( .IN1(n11276), .IN2(n11277), .IN3(n11269), .Q(n11275) );
  OR2X1 U32935 ( .IN1(n11278), .IN2(n11279), .Q(n11276) );
  AND3X1 U32936 ( .IN1(n13133), .IN2(n13134), .IN3(n13126), .Q(n13132) );
  OR2X1 U32937 ( .IN1(n13135), .IN2(n13136), .Q(n13133) );
  AND3X1 U32938 ( .IN1(n12824), .IN2(n12825), .IN3(n12817), .Q(n12823) );
  OR2X1 U32939 ( .IN1(n12826), .IN2(n12827), .Q(n12824) );
  AND3X1 U32940 ( .IN1(n10657), .IN2(n10658), .IN3(n10650), .Q(n10656) );
  OR2X1 U32941 ( .IN1(n10659), .IN2(n10660), .Q(n10657) );
  AND3X1 U32942 ( .IN1(n12515), .IN2(n12516), .IN3(n12508), .Q(n12514) );
  OR2X1 U32943 ( .IN1(n12517), .IN2(n12518), .Q(n12515) );
  AND3X1 U32944 ( .IN1(n12206), .IN2(n12207), .IN3(n12199), .Q(n12205) );
  OR2X1 U32945 ( .IN1(n12208), .IN2(n12209), .Q(n12206) );
  AND3X1 U32946 ( .IN1(n10038), .IN2(n10039), .IN3(n10031), .Q(n10037) );
  OR2X1 U32947 ( .IN1(n10040), .IN2(n10041), .Q(n10038) );
  AND3X1 U32948 ( .IN1(n11896), .IN2(n11897), .IN3(n11889), .Q(n11895) );
  OR2X1 U32949 ( .IN1(n11898), .IN2(n11899), .Q(n11896) );
  AND3X1 U32950 ( .IN1(n11586), .IN2(n11587), .IN3(n11579), .Q(n11585) );
  OR2X1 U32951 ( .IN1(n11588), .IN2(n11589), .Q(n11586) );
  AND3X1 U32952 ( .IN1(n9417), .IN2(n9418), .IN3(n9410), .Q(n9416) );
  OR2X1 U32953 ( .IN1(n9419), .IN2(n9420), .Q(n9417) );
  AND3X1 U32954 ( .IN1(n14015), .IN2(n14016), .IN3(n14008), .Q(n14014) );
  OR2X1 U32955 ( .IN1(n14017), .IN2(n14018), .Q(n14015) );
  OA21X1 U32956 ( .IN1(n3224), .IN2(n13900), .IN3(n13901), .Q(n13886) );
  OA21X1 U32957 ( .IN1(n3146), .IN2(n13902), .IN3(n13903), .Q(n13900) );
  OA21X1 U32958 ( .IN1(n13832), .IN2(n13833), .IN3(n13834), .Q(n13817) );
  OA21X1 U32959 ( .IN1(n13835), .IN2(n13836), .IN3(n13837), .Q(n13833) );
  OA21X1 U32960 ( .IN1(n13769), .IN2(n13770), .IN3(n13771), .Q(n13753) );
  OA21X1 U32961 ( .IN1(n13772), .IN2(n13773), .IN3(n13774), .Q(n13770) );
  OA21X1 U32962 ( .IN1(n13673), .IN2(n13706), .IN3(n13707), .Q(n13692) );
  OA21X1 U32963 ( .IN1(n13675), .IN2(n13708), .IN3(n13709), .Q(n13706) );
  OA21X1 U32964 ( .IN1(n3228), .IN2(n13591), .IN3(n13592), .Q(n13577) );
  OA21X1 U32965 ( .IN1(n3152), .IN2(n13593), .IN3(n13594), .Q(n13591) );
  OA21X1 U32966 ( .IN1(n13523), .IN2(n13524), .IN3(n13525), .Q(n13508) );
  OA21X1 U32967 ( .IN1(n13526), .IN2(n13527), .IN3(n13528), .Q(n13524) );
  OA21X1 U32968 ( .IN1(n13460), .IN2(n13461), .IN3(n13462), .Q(n13444) );
  OA21X1 U32969 ( .IN1(n13463), .IN2(n13464), .IN3(n13465), .Q(n13461) );
  OA21X1 U32970 ( .IN1(n13364), .IN2(n13397), .IN3(n13398), .Q(n13383) );
  OA21X1 U32971 ( .IN1(n13366), .IN2(n13399), .IN3(n13400), .Q(n13397) );
  OA21X1 U32972 ( .IN1(n3196), .IN2(n11425), .IN3(n11426), .Q(n11411) );
  OA21X1 U32973 ( .IN1(n3104), .IN2(n11427), .IN3(n11428), .Q(n11425) );
  OA21X1 U32974 ( .IN1(n11357), .IN2(n11358), .IN3(n11359), .Q(n11342) );
  OA21X1 U32975 ( .IN1(n11360), .IN2(n11361), .IN3(n11362), .Q(n11358) );
  OA21X1 U32976 ( .IN1(n11294), .IN2(n11295), .IN3(n11296), .Q(n11278) );
  OA21X1 U32977 ( .IN1(n11297), .IN2(n11298), .IN3(n11299), .Q(n11295) );
  OA21X1 U32978 ( .IN1(n11198), .IN2(n11231), .IN3(n11232), .Q(n11217) );
  OA21X1 U32979 ( .IN1(n11200), .IN2(n11233), .IN3(n11234), .Q(n11231) );
  OA21X1 U32980 ( .IN1(n3232), .IN2(n13282), .IN3(n13283), .Q(n13268) );
  OA21X1 U32981 ( .IN1(n3158), .IN2(n13284), .IN3(n13285), .Q(n13282) );
  OA21X1 U32982 ( .IN1(n13214), .IN2(n13215), .IN3(n13216), .Q(n13199) );
  OA21X1 U32983 ( .IN1(n13217), .IN2(n13218), .IN3(n13219), .Q(n13215) );
  OA21X1 U32984 ( .IN1(n13151), .IN2(n13152), .IN3(n13153), .Q(n13135) );
  OA21X1 U32985 ( .IN1(n13154), .IN2(n13155), .IN3(n13156), .Q(n13152) );
  OA21X1 U32986 ( .IN1(n13055), .IN2(n13088), .IN3(n13089), .Q(n13074) );
  OA21X1 U32987 ( .IN1(n13057), .IN2(n13090), .IN3(n13091), .Q(n13088) );
  OA21X1 U32988 ( .IN1(n3236), .IN2(n12973), .IN3(n12974), .Q(n12959) );
  OA21X1 U32989 ( .IN1(n3164), .IN2(n12975), .IN3(n12976), .Q(n12973) );
  OA21X1 U32990 ( .IN1(n12905), .IN2(n12906), .IN3(n12907), .Q(n12890) );
  OA21X1 U32991 ( .IN1(n12908), .IN2(n12909), .IN3(n12910), .Q(n12906) );
  OA21X1 U32992 ( .IN1(n12842), .IN2(n12843), .IN3(n12844), .Q(n12826) );
  OA21X1 U32993 ( .IN1(n12845), .IN2(n12846), .IN3(n12847), .Q(n12843) );
  OA21X1 U32994 ( .IN1(n12746), .IN2(n12779), .IN3(n12780), .Q(n12765) );
  OA21X1 U32995 ( .IN1(n12748), .IN2(n12781), .IN3(n12782), .Q(n12779) );
  OA21X1 U32996 ( .IN1(n3200), .IN2(n11116), .IN3(n11117), .Q(n11102) );
  OA21X1 U32997 ( .IN1(n3110), .IN2(n11118), .IN3(n11119), .Q(n11116) );
  OA21X1 U32998 ( .IN1(n11048), .IN2(n11049), .IN3(n11050), .Q(n11033) );
  OA21X1 U32999 ( .IN1(n11051), .IN2(n11052), .IN3(n11053), .Q(n11049) );
  OA21X1 U33000 ( .IN1(n10985), .IN2(n10986), .IN3(n10987), .Q(n10969) );
  OA21X1 U33001 ( .IN1(n10988), .IN2(n10989), .IN3(n10990), .Q(n10986) );
  OA21X1 U33002 ( .IN1(n10889), .IN2(n10922), .IN3(n10923), .Q(n10908) );
  OA21X1 U33003 ( .IN1(n10891), .IN2(n10924), .IN3(n10925), .Q(n10922) );
  OA21X1 U33004 ( .IN1(n3204), .IN2(n10806), .IN3(n10807), .Q(n10792) );
  OA21X1 U33005 ( .IN1(n3116), .IN2(n10808), .IN3(n10809), .Q(n10806) );
  OA21X1 U33006 ( .IN1(n10738), .IN2(n10739), .IN3(n10740), .Q(n10723) );
  OA21X1 U33007 ( .IN1(n10741), .IN2(n10742), .IN3(n10743), .Q(n10739) );
  OA21X1 U33008 ( .IN1(n10675), .IN2(n10676), .IN3(n10677), .Q(n10659) );
  OA21X1 U33009 ( .IN1(n10678), .IN2(n10679), .IN3(n10680), .Q(n10676) );
  OA21X1 U33010 ( .IN1(n10579), .IN2(n10612), .IN3(n10613), .Q(n10598) );
  OA21X1 U33011 ( .IN1(n10581), .IN2(n10614), .IN3(n10615), .Q(n10612) );
  OA21X1 U33012 ( .IN1(n3240), .IN2(n12664), .IN3(n12665), .Q(n12650) );
  OA21X1 U33013 ( .IN1(n3170), .IN2(n12666), .IN3(n12667), .Q(n12664) );
  OA21X1 U33014 ( .IN1(n12596), .IN2(n12597), .IN3(n12598), .Q(n12581) );
  OA21X1 U33015 ( .IN1(n12599), .IN2(n12600), .IN3(n12601), .Q(n12597) );
  OA21X1 U33016 ( .IN1(n12533), .IN2(n12534), .IN3(n12535), .Q(n12517) );
  OA21X1 U33017 ( .IN1(n12536), .IN2(n12537), .IN3(n12538), .Q(n12534) );
  OA21X1 U33018 ( .IN1(n12437), .IN2(n12470), .IN3(n12471), .Q(n12456) );
  OA21X1 U33019 ( .IN1(n12439), .IN2(n12472), .IN3(n12473), .Q(n12470) );
  OA21X1 U33020 ( .IN1(n3244), .IN2(n12355), .IN3(n12356), .Q(n12341) );
  OA21X1 U33021 ( .IN1(n3176), .IN2(n12357), .IN3(n12358), .Q(n12355) );
  OA21X1 U33022 ( .IN1(n12287), .IN2(n12288), .IN3(n12289), .Q(n12272) );
  OA21X1 U33023 ( .IN1(n12290), .IN2(n12291), .IN3(n12292), .Q(n12288) );
  OA21X1 U33024 ( .IN1(n12224), .IN2(n12225), .IN3(n12226), .Q(n12208) );
  OA21X1 U33025 ( .IN1(n12227), .IN2(n12228), .IN3(n12229), .Q(n12225) );
  OA21X1 U33026 ( .IN1(n12128), .IN2(n12161), .IN3(n12162), .Q(n12147) );
  OA21X1 U33027 ( .IN1(n12130), .IN2(n12163), .IN3(n12164), .Q(n12161) );
  OA21X1 U33028 ( .IN1(n3208), .IN2(n10497), .IN3(n10498), .Q(n10483) );
  OA21X1 U33029 ( .IN1(n3122), .IN2(n10499), .IN3(n10500), .Q(n10497) );
  OA21X1 U33030 ( .IN1(n10429), .IN2(n10430), .IN3(n10431), .Q(n10414) );
  OA21X1 U33031 ( .IN1(n10432), .IN2(n10433), .IN3(n10434), .Q(n10430) );
  OA21X1 U33032 ( .IN1(n10366), .IN2(n10367), .IN3(n10368), .Q(n10350) );
  OA21X1 U33033 ( .IN1(n10369), .IN2(n10370), .IN3(n10371), .Q(n10367) );
  OA21X1 U33034 ( .IN1(n10270), .IN2(n10303), .IN3(n10304), .Q(n10289) );
  OA21X1 U33035 ( .IN1(n10272), .IN2(n10305), .IN3(n10306), .Q(n10303) );
  OA21X1 U33036 ( .IN1(n3212), .IN2(n10187), .IN3(n10188), .Q(n10173) );
  OA21X1 U33037 ( .IN1(n3128), .IN2(n10189), .IN3(n10190), .Q(n10187) );
  OA21X1 U33038 ( .IN1(n10119), .IN2(n10120), .IN3(n10121), .Q(n10104) );
  OA21X1 U33039 ( .IN1(n10122), .IN2(n10123), .IN3(n10124), .Q(n10120) );
  OA21X1 U33040 ( .IN1(n10056), .IN2(n10057), .IN3(n10058), .Q(n10040) );
  OA21X1 U33041 ( .IN1(n10059), .IN2(n10060), .IN3(n10061), .Q(n10057) );
  OA21X1 U33042 ( .IN1(n9960), .IN2(n9993), .IN3(n9994), .Q(n9979) );
  OA21X1 U33043 ( .IN1(n9962), .IN2(n9995), .IN3(n9996), .Q(n9993) );
  OA21X1 U33044 ( .IN1(n3248), .IN2(n12045), .IN3(n12046), .Q(n12031) );
  OA21X1 U33045 ( .IN1(n3182), .IN2(n12047), .IN3(n12048), .Q(n12045) );
  OA21X1 U33046 ( .IN1(n11977), .IN2(n11978), .IN3(n11979), .Q(n11962) );
  OA21X1 U33047 ( .IN1(n11980), .IN2(n11981), .IN3(n11982), .Q(n11978) );
  OA21X1 U33048 ( .IN1(n11914), .IN2(n11915), .IN3(n11916), .Q(n11898) );
  OA21X1 U33049 ( .IN1(n11917), .IN2(n11918), .IN3(n11919), .Q(n11915) );
  OA21X1 U33050 ( .IN1(n11818), .IN2(n11851), .IN3(n11852), .Q(n11837) );
  OA21X1 U33051 ( .IN1(n11820), .IN2(n11853), .IN3(n11854), .Q(n11851) );
  OA21X1 U33052 ( .IN1(n3252), .IN2(n11735), .IN3(n11736), .Q(n11721) );
  OA21X1 U33053 ( .IN1(n3188), .IN2(n11737), .IN3(n11738), .Q(n11735) );
  OA21X1 U33054 ( .IN1(n11667), .IN2(n11668), .IN3(n11669), .Q(n11652) );
  OA21X1 U33055 ( .IN1(n11670), .IN2(n11671), .IN3(n11672), .Q(n11668) );
  OA21X1 U33056 ( .IN1(n11604), .IN2(n11605), .IN3(n11606), .Q(n11588) );
  OA21X1 U33057 ( .IN1(n11607), .IN2(n11608), .IN3(n11609), .Q(n11605) );
  OA21X1 U33058 ( .IN1(n11508), .IN2(n11541), .IN3(n11542), .Q(n11527) );
  OA21X1 U33059 ( .IN1(n11510), .IN2(n11543), .IN3(n11544), .Q(n11541) );
  OA21X1 U33060 ( .IN1(n3216), .IN2(n9877), .IN3(n9878), .Q(n9863) );
  OA21X1 U33061 ( .IN1(n3134), .IN2(n9879), .IN3(n9880), .Q(n9877) );
  OA21X1 U33062 ( .IN1(n9809), .IN2(n9810), .IN3(n9811), .Q(n9794) );
  OA21X1 U33063 ( .IN1(n9812), .IN2(n9813), .IN3(n9814), .Q(n9810) );
  OA21X1 U33064 ( .IN1(n9746), .IN2(n9747), .IN3(n9748), .Q(n9730) );
  OA21X1 U33065 ( .IN1(n9749), .IN2(n9750), .IN3(n9751), .Q(n9747) );
  OA21X1 U33066 ( .IN1(n9650), .IN2(n9683), .IN3(n9684), .Q(n9669) );
  OA21X1 U33067 ( .IN1(n9652), .IN2(n9685), .IN3(n9686), .Q(n9683) );
  OA21X1 U33068 ( .IN1(n3220), .IN2(n9566), .IN3(n9567), .Q(n9552) );
  OA21X1 U33069 ( .IN1(n3140), .IN2(n9568), .IN3(n9569), .Q(n9566) );
  OA21X1 U33070 ( .IN1(n9498), .IN2(n9499), .IN3(n9500), .Q(n9483) );
  OA21X1 U33071 ( .IN1(n9501), .IN2(n9502), .IN3(n9503), .Q(n9499) );
  OA21X1 U33072 ( .IN1(n9435), .IN2(n9436), .IN3(n9437), .Q(n9419) );
  OA21X1 U33073 ( .IN1(n9438), .IN2(n9439), .IN3(n9440), .Q(n9436) );
  OA21X1 U33074 ( .IN1(n9339), .IN2(n9372), .IN3(n9373), .Q(n9358) );
  OA21X1 U33075 ( .IN1(n9341), .IN2(n9374), .IN3(n9375), .Q(n9372) );
  OA21X1 U33076 ( .IN1(n13965), .IN2(n13966), .IN3(n13967), .Q(n13949) );
  OA21X1 U33077 ( .IN1(n13968), .IN2(n13969), .IN3(n13970), .Q(n13966) );
  OA21X1 U33078 ( .IN1(n3190), .IN2(n14174), .IN3(n14175), .Q(n14160) );
  OA21X1 U33079 ( .IN1(n3094), .IN2(n14176), .IN3(n14177), .Q(n14174) );
  OA21X1 U33080 ( .IN1(n14105), .IN2(n14106), .IN3(n14107), .Q(n14089) );
  OA21X1 U33081 ( .IN1(n14108), .IN2(n14109), .IN3(n14110), .Q(n14106) );
  OA21X1 U33082 ( .IN1(n14033), .IN2(n14034), .IN3(n14035), .Q(n14017) );
  OA21X1 U33083 ( .IN1(n14036), .IN2(n14037), .IN3(n14038), .Q(n14034) );
  OA21X1 U33084 ( .IN1(n3323), .IN2(n13914), .IN3(n13885), .Q(n13881) );
  OA21X1 U33085 ( .IN1(n3224), .IN2(n13897), .IN3(n13901), .Q(n13914) );
  OA21X1 U33086 ( .IN1(n3331), .IN2(n13605), .IN3(n13576), .Q(n13572) );
  OA21X1 U33087 ( .IN1(n3228), .IN2(n13588), .IN3(n13592), .Q(n13605) );
  OA21X1 U33088 ( .IN1(n3267), .IN2(n11439), .IN3(n11410), .Q(n11406) );
  OA21X1 U33089 ( .IN1(n3196), .IN2(n11422), .IN3(n11426), .Q(n11439) );
  OA21X1 U33090 ( .IN1(n3339), .IN2(n13296), .IN3(n13267), .Q(n13263) );
  OA21X1 U33091 ( .IN1(n3232), .IN2(n13279), .IN3(n13283), .Q(n13296) );
  OA21X1 U33092 ( .IN1(n3347), .IN2(n12987), .IN3(n12958), .Q(n12954) );
  OA21X1 U33093 ( .IN1(n3236), .IN2(n12970), .IN3(n12974), .Q(n12987) );
  OA21X1 U33094 ( .IN1(n3275), .IN2(n11130), .IN3(n11101), .Q(n11097) );
  OA21X1 U33095 ( .IN1(n3200), .IN2(n11113), .IN3(n11117), .Q(n11130) );
  OA21X1 U33096 ( .IN1(n3283), .IN2(n10820), .IN3(n10791), .Q(n10787) );
  OA21X1 U33097 ( .IN1(n3204), .IN2(n10803), .IN3(n10807), .Q(n10820) );
  OA21X1 U33098 ( .IN1(n3355), .IN2(n12678), .IN3(n12649), .Q(n12645) );
  OA21X1 U33099 ( .IN1(n3240), .IN2(n12661), .IN3(n12665), .Q(n12678) );
  OA21X1 U33100 ( .IN1(n3363), .IN2(n12369), .IN3(n12340), .Q(n12336) );
  OA21X1 U33101 ( .IN1(n3244), .IN2(n12352), .IN3(n12356), .Q(n12369) );
  OA21X1 U33102 ( .IN1(n3291), .IN2(n10511), .IN3(n10482), .Q(n10478) );
  OA21X1 U33103 ( .IN1(n3208), .IN2(n10494), .IN3(n10498), .Q(n10511) );
  OA21X1 U33104 ( .IN1(n3299), .IN2(n10201), .IN3(n10172), .Q(n10168) );
  OA21X1 U33105 ( .IN1(n3212), .IN2(n10184), .IN3(n10188), .Q(n10201) );
  OA21X1 U33106 ( .IN1(n3371), .IN2(n12059), .IN3(n12030), .Q(n12026) );
  OA21X1 U33107 ( .IN1(n3248), .IN2(n12042), .IN3(n12046), .Q(n12059) );
  OA21X1 U33108 ( .IN1(n3379), .IN2(n11749), .IN3(n11720), .Q(n11716) );
  OA21X1 U33109 ( .IN1(n3252), .IN2(n11732), .IN3(n11736), .Q(n11749) );
  OA21X1 U33110 ( .IN1(n3307), .IN2(n9891), .IN3(n9862), .Q(n9858) );
  OA21X1 U33111 ( .IN1(n3216), .IN2(n9874), .IN3(n9878), .Q(n9891) );
  OA21X1 U33112 ( .IN1(n3315), .IN2(n9580), .IN3(n9551), .Q(n9547) );
  OA21X1 U33113 ( .IN1(n3220), .IN2(n9563), .IN3(n9567), .Q(n9580) );
  OA21X1 U33114 ( .IN1(n3255), .IN2(n14188), .IN3(n14159), .Q(n14155) );
  OA21X1 U33115 ( .IN1(n3190), .IN2(n14171), .IN3(n14175), .Q(n14188) );
  OA21X1 U33116 ( .IN1(n13927), .IN2(n2979), .IN3(n13902), .Q(n13916) );
  OA21X1 U33117 ( .IN1(n13862), .IN2(n13847), .IN3(n13836), .Q(n13849) );
  OA21X1 U33118 ( .IN1(n13731), .IN2(n13676), .IN3(n13708), .Q(n13719) );
  OA21X1 U33119 ( .IN1(n13618), .IN2(n2995), .IN3(n13593), .Q(n13607) );
  OA21X1 U33120 ( .IN1(n13553), .IN2(n13538), .IN3(n13527), .Q(n13540) );
  OA21X1 U33121 ( .IN1(n13422), .IN2(n13367), .IN3(n13399), .Q(n13410) );
  OA21X1 U33122 ( .IN1(n11452), .IN2(n2867), .IN3(n11427), .Q(n11441) );
  OA21X1 U33123 ( .IN1(n11387), .IN2(n11372), .IN3(n11361), .Q(n11374) );
  OA21X1 U33124 ( .IN1(n11256), .IN2(n11201), .IN3(n11233), .Q(n11244) );
  OA21X1 U33125 ( .IN1(n13309), .IN2(n3011), .IN3(n13284), .Q(n13298) );
  OA21X1 U33126 ( .IN1(n13244), .IN2(n13229), .IN3(n13218), .Q(n13231) );
  OA21X1 U33127 ( .IN1(n13113), .IN2(n13058), .IN3(n13090), .Q(n13101) );
  OA21X1 U33128 ( .IN1(n13000), .IN2(n3027), .IN3(n12975), .Q(n12989) );
  OA21X1 U33129 ( .IN1(n12935), .IN2(n12920), .IN3(n12909), .Q(n12922) );
  OA21X1 U33130 ( .IN1(n12804), .IN2(n12749), .IN3(n12781), .Q(n12792) );
  OA21X1 U33131 ( .IN1(n11143), .IN2(n2883), .IN3(n11118), .Q(n11132) );
  OA21X1 U33132 ( .IN1(n11078), .IN2(n11063), .IN3(n11052), .Q(n11065) );
  OA21X1 U33133 ( .IN1(n10947), .IN2(n10892), .IN3(n10924), .Q(n10935) );
  OA21X1 U33134 ( .IN1(n10833), .IN2(n2899), .IN3(n10808), .Q(n10822) );
  OA21X1 U33135 ( .IN1(n10768), .IN2(n10753), .IN3(n10742), .Q(n10755) );
  OA21X1 U33136 ( .IN1(n10637), .IN2(n10582), .IN3(n10614), .Q(n10625) );
  OA21X1 U33137 ( .IN1(n12691), .IN2(n3043), .IN3(n12666), .Q(n12680) );
  OA21X1 U33138 ( .IN1(n12626), .IN2(n12611), .IN3(n12600), .Q(n12613) );
  OA21X1 U33139 ( .IN1(n12495), .IN2(n12440), .IN3(n12472), .Q(n12483) );
  OA21X1 U33140 ( .IN1(n12382), .IN2(n3059), .IN3(n12357), .Q(n12371) );
  OA21X1 U33141 ( .IN1(n12317), .IN2(n12302), .IN3(n12291), .Q(n12304) );
  OA21X1 U33142 ( .IN1(n12186), .IN2(n12131), .IN3(n12163), .Q(n12174) );
  OA21X1 U33143 ( .IN1(n10524), .IN2(n2915), .IN3(n10499), .Q(n10513) );
  OA21X1 U33144 ( .IN1(n10459), .IN2(n10444), .IN3(n10433), .Q(n10446) );
  OA21X1 U33145 ( .IN1(n10328), .IN2(n10273), .IN3(n10305), .Q(n10316) );
  OA21X1 U33146 ( .IN1(n10214), .IN2(n2931), .IN3(n10189), .Q(n10203) );
  OA21X1 U33147 ( .IN1(n10149), .IN2(n10134), .IN3(n10123), .Q(n10136) );
  OA21X1 U33148 ( .IN1(n10018), .IN2(n9963), .IN3(n9995), .Q(n10006) );
  OA21X1 U33149 ( .IN1(n12072), .IN2(n3075), .IN3(n12047), .Q(n12061) );
  OA21X1 U33150 ( .IN1(n12007), .IN2(n11992), .IN3(n11981), .Q(n11994) );
  OA21X1 U33151 ( .IN1(n11876), .IN2(n11821), .IN3(n11853), .Q(n11864) );
  OA21X1 U33152 ( .IN1(n11762), .IN2(n3091), .IN3(n11737), .Q(n11751) );
  OA21X1 U33153 ( .IN1(n11697), .IN2(n11682), .IN3(n11671), .Q(n11684) );
  OA21X1 U33154 ( .IN1(n11566), .IN2(n11511), .IN3(n11543), .Q(n11554) );
  OA21X1 U33155 ( .IN1(n9904), .IN2(n2947), .IN3(n9879), .Q(n9893) );
  OA21X1 U33156 ( .IN1(n9839), .IN2(n9824), .IN3(n9813), .Q(n9826) );
  OA21X1 U33157 ( .IN1(n9708), .IN2(n9653), .IN3(n9685), .Q(n9696) );
  OA21X1 U33158 ( .IN1(n9593), .IN2(n2963), .IN3(n9568), .Q(n9582) );
  OA21X1 U33159 ( .IN1(n9528), .IN2(n9513), .IN3(n9502), .Q(n9515) );
  OA21X1 U33160 ( .IN1(n9397), .IN2(n9342), .IN3(n9374), .Q(n9385) );
  OA21X1 U33161 ( .IN1(n13995), .IN2(n13980), .IN3(n13969), .Q(n13982) );
  OA21X1 U33162 ( .IN1(n14201), .IN2(n2842), .IN3(n14176), .Q(n14190) );
  OA21X1 U33163 ( .IN1(n14135), .IN2(n14120), .IN3(n14109), .Q(n14122) );
  NAND2X0 U33164 ( .IN1(n13928), .IN2(n13907), .QN(n13896) );
  NAND2X0 U33165 ( .IN1(n13619), .IN2(n13598), .QN(n13587) );
  NAND2X0 U33166 ( .IN1(n11453), .IN2(n11432), .QN(n11421) );
  NAND2X0 U33167 ( .IN1(n13310), .IN2(n13289), .QN(n13278) );
  NAND2X0 U33168 ( .IN1(n13001), .IN2(n12980), .QN(n12969) );
  NAND2X0 U33169 ( .IN1(n11144), .IN2(n11123), .QN(n11112) );
  NAND2X0 U33170 ( .IN1(n10834), .IN2(n10813), .QN(n10802) );
  NAND2X0 U33171 ( .IN1(n12692), .IN2(n12671), .QN(n12660) );
  NAND2X0 U33172 ( .IN1(n12383), .IN2(n12362), .QN(n12351) );
  NAND2X0 U33173 ( .IN1(n10525), .IN2(n10504), .QN(n10493) );
  NAND2X0 U33174 ( .IN1(n10215), .IN2(n10194), .QN(n10183) );
  NAND2X0 U33175 ( .IN1(n12073), .IN2(n12052), .QN(n12041) );
  NAND2X0 U33176 ( .IN1(n11763), .IN2(n11742), .QN(n11731) );
  NAND2X0 U33177 ( .IN1(n9905), .IN2(n9884), .QN(n9873) );
  NAND2X0 U33178 ( .IN1(n9594), .IN2(n9573), .QN(n9562) );
  NAND2X0 U33179 ( .IN1(n14202), .IN2(n14181), .QN(n14170) );
  NAND2X0 U33180 ( .IN1(n13757), .IN2(n13758), .QN(n13755) );
  NAND2X0 U33181 ( .IN1(n13448), .IN2(n13449), .QN(n13446) );
  NAND2X0 U33182 ( .IN1(n11282), .IN2(n11283), .QN(n11280) );
  NAND2X0 U33183 ( .IN1(n13139), .IN2(n13140), .QN(n13137) );
  NAND2X0 U33184 ( .IN1(n12830), .IN2(n12831), .QN(n12828) );
  NAND2X0 U33185 ( .IN1(n10973), .IN2(n10974), .QN(n10971) );
  NAND2X0 U33186 ( .IN1(n10663), .IN2(n10664), .QN(n10661) );
  NAND2X0 U33187 ( .IN1(n12521), .IN2(n12522), .QN(n12519) );
  NAND2X0 U33188 ( .IN1(n12212), .IN2(n12213), .QN(n12210) );
  NAND2X0 U33189 ( .IN1(n10354), .IN2(n10355), .QN(n10352) );
  NAND2X0 U33190 ( .IN1(n10044), .IN2(n10045), .QN(n10042) );
  NAND2X0 U33191 ( .IN1(n11902), .IN2(n11903), .QN(n11900) );
  NAND2X0 U33192 ( .IN1(n11592), .IN2(n11593), .QN(n11590) );
  NAND2X0 U33193 ( .IN1(n9734), .IN2(n9735), .QN(n9732) );
  NAND2X0 U33194 ( .IN1(n9423), .IN2(n9424), .QN(n9421) );
  NAND2X0 U33195 ( .IN1(n14021), .IN2(n14022), .QN(n14019) );
  AND3X1 U33196 ( .IN1(n13442), .IN2(n13443), .IN3(n13435), .Q(n13441) );
  OR2X1 U33197 ( .IN1(n13444), .IN2(n13445), .Q(n13442) );
  AND3X1 U33198 ( .IN1(n13197), .IN2(n13198), .IN3(n13191), .Q(n13192) );
  OR2X1 U33199 ( .IN1(n13199), .IN2(n13200), .Q(n13197) );
  AND3X1 U33200 ( .IN1(n12888), .IN2(n12889), .IN3(n12882), .Q(n12883) );
  OR2X1 U33201 ( .IN1(n12890), .IN2(n12891), .Q(n12888) );
  AND3X1 U33202 ( .IN1(n11031), .IN2(n11032), .IN3(n11025), .Q(n11026) );
  OR2X1 U33203 ( .IN1(n11033), .IN2(n11034), .Q(n11031) );
  AND3X1 U33204 ( .IN1(n10721), .IN2(n10722), .IN3(n10715), .Q(n10716) );
  OR2X1 U33205 ( .IN1(n10723), .IN2(n10724), .Q(n10721) );
  AND3X1 U33206 ( .IN1(n10412), .IN2(n10413), .IN3(n10406), .Q(n10407) );
  OR2X1 U33207 ( .IN1(n10414), .IN2(n10415), .Q(n10412) );
  AND3X1 U33208 ( .IN1(n10102), .IN2(n10103), .IN3(n10096), .Q(n10097) );
  OR2X1 U33209 ( .IN1(n10104), .IN2(n10105), .Q(n10102) );
  AND3X1 U33210 ( .IN1(n11960), .IN2(n11961), .IN3(n11954), .Q(n11955) );
  OR2X1 U33211 ( .IN1(n11962), .IN2(n11963), .Q(n11960) );
  AND3X1 U33212 ( .IN1(n11650), .IN2(n11651), .IN3(n11644), .Q(n11645) );
  OR2X1 U33213 ( .IN1(n11652), .IN2(n11653), .Q(n11650) );
  NAND2X0 U33214 ( .IN1(n18189), .IN2(n18036), .QN(n14069) );
  NAND2X0 U33215 ( .IN1(n18190), .IN2(n18035), .QN(n14068) );
  NAND2X0 U33216 ( .IN1(n18191), .IN2(n18032), .QN(n13657) );
  NAND2X0 U33217 ( .IN1(n18037), .IN2(n18201), .QN(n13348) );
  NAND2X0 U33218 ( .IN1(n18038), .IN2(n18202), .QN(n11182) );
  NAND2X0 U33219 ( .IN1(n18192), .IN2(n18033), .QN(n12421) );
  NAND2X0 U33220 ( .IN1(n18039), .IN2(n18203), .QN(n12112) );
  NAND2X0 U33221 ( .IN1(n18193), .IN2(n18034), .QN(n9634) );
  NAND2X0 U33222 ( .IN1(n18040), .IN2(n18204), .QN(n9323) );
  NAND2X0 U33223 ( .IN1(n18194), .IN2(n18029), .QN(n13660) );
  NAND2X0 U33224 ( .IN1(n18041), .IN2(n18197), .QN(n13351) );
  NAND2X0 U33225 ( .IN1(n18042), .IN2(n18198), .QN(n11185) );
  NAND2X0 U33226 ( .IN1(n18195), .IN2(n18030), .QN(n12424) );
  NAND2X0 U33227 ( .IN1(n18043), .IN2(n18199), .QN(n12115) );
  NAND2X0 U33228 ( .IN1(n18196), .IN2(n18031), .QN(n9637) );
  NAND2X0 U33229 ( .IN1(n18044), .IN2(n18200), .QN(n9326) );
  NAND2X0 U33230 ( .IN1(n18205), .IN2(n18049), .QN(n13039) );
  NAND2X0 U33231 ( .IN1(n18206), .IN2(n18050), .QN(n10873) );
  NAND2X0 U33232 ( .IN1(n18207), .IN2(n18051), .QN(n10254) );
  NAND2X0 U33233 ( .IN1(n18208), .IN2(n18052), .QN(n11802) );
  NAND2X0 U33234 ( .IN1(n18209), .IN2(n18045), .QN(n13042) );
  NAND2X0 U33235 ( .IN1(n18210), .IN2(n18046), .QN(n10876) );
  NAND2X0 U33236 ( .IN1(n18211), .IN2(n18047), .QN(n10257) );
  NAND2X0 U33237 ( .IN1(n18212), .IN2(n18048), .QN(n11805) );
  NAND2X0 U33238 ( .IN1(n18053), .IN2(n18217), .QN(n12730) );
  NAND2X0 U33239 ( .IN1(n18054), .IN2(n18218), .QN(n10563) );
  NAND2X0 U33240 ( .IN1(n18055), .IN2(n18219), .QN(n9944) );
  NAND2X0 U33241 ( .IN1(n18056), .IN2(n18220), .QN(n11492) );
  NAND2X0 U33242 ( .IN1(n18057), .IN2(n18213), .QN(n12733) );
  NAND2X0 U33243 ( .IN1(n18058), .IN2(n18214), .QN(n10566) );
  NAND2X0 U33244 ( .IN1(n18059), .IN2(n18215), .QN(n9947) );
  NAND2X0 U33245 ( .IN1(n18060), .IN2(n18216), .QN(n11495) );
  INVX0 U33246 ( .IN(n13838), .QN(n3432) );
  INVX0 U33247 ( .IN(n13529), .QN(n3436) );
  INVX0 U33248 ( .IN(n11363), .QN(n3404) );
  INVX0 U33249 ( .IN(n13220), .QN(n3440) );
  INVX0 U33250 ( .IN(n12911), .QN(n3444) );
  INVX0 U33251 ( .IN(n11054), .QN(n3408) );
  INVX0 U33252 ( .IN(n10744), .QN(n3412) );
  INVX0 U33253 ( .IN(n12602), .QN(n3448) );
  INVX0 U33254 ( .IN(n12293), .QN(n3452) );
  INVX0 U33255 ( .IN(n10435), .QN(n3416) );
  INVX0 U33256 ( .IN(n10125), .QN(n3420) );
  INVX0 U33257 ( .IN(n11983), .QN(n3456) );
  INVX0 U33258 ( .IN(n11673), .QN(n3460) );
  INVX0 U33259 ( .IN(n9815), .QN(n3424) );
  INVX0 U33260 ( .IN(n9504), .QN(n3428) );
  INVX0 U33261 ( .IN(n13971), .QN(n3400) );
  INVX0 U33262 ( .IN(n14111), .QN(n3401) );
  INVX0 U33263 ( .IN(n13883), .QN(n3433) );
  INVX0 U33264 ( .IN(n13574), .QN(n3437) );
  INVX0 U33265 ( .IN(n11408), .QN(n3405) );
  INVX0 U33266 ( .IN(n13265), .QN(n3441) );
  INVX0 U33267 ( .IN(n12956), .QN(n3445) );
  INVX0 U33268 ( .IN(n11099), .QN(n3409) );
  INVX0 U33269 ( .IN(n10789), .QN(n3413) );
  INVX0 U33270 ( .IN(n12647), .QN(n3449) );
  INVX0 U33271 ( .IN(n12338), .QN(n3453) );
  INVX0 U33272 ( .IN(n10480), .QN(n3417) );
  INVX0 U33273 ( .IN(n10170), .QN(n3421) );
  INVX0 U33274 ( .IN(n12028), .QN(n3457) );
  INVX0 U33275 ( .IN(n11718), .QN(n3461) );
  INVX0 U33276 ( .IN(n9860), .QN(n3425) );
  INVX0 U33277 ( .IN(n9549), .QN(n3429) );
  INVX0 U33278 ( .IN(n14157), .QN(n3399) );
  INVX0 U33279 ( .IN(n13894), .QN(n3224) );
  INVX0 U33280 ( .IN(n13585), .QN(n3228) );
  INVX0 U33281 ( .IN(n11419), .QN(n3196) );
  INVX0 U33282 ( .IN(n13276), .QN(n3232) );
  INVX0 U33283 ( .IN(n12967), .QN(n3236) );
  INVX0 U33284 ( .IN(n11110), .QN(n3200) );
  INVX0 U33285 ( .IN(n10800), .QN(n3204) );
  INVX0 U33286 ( .IN(n12658), .QN(n3240) );
  INVX0 U33287 ( .IN(n12349), .QN(n3244) );
  INVX0 U33288 ( .IN(n10491), .QN(n3208) );
  INVX0 U33289 ( .IN(n10181), .QN(n3212) );
  INVX0 U33290 ( .IN(n12039), .QN(n3248) );
  INVX0 U33291 ( .IN(n11729), .QN(n3252) );
  INVX0 U33292 ( .IN(n9871), .QN(n3216) );
  INVX0 U33293 ( .IN(n9560), .QN(n3220) );
  INVX0 U33294 ( .IN(n14168), .QN(n3190) );
  INVX0 U33295 ( .IN(n13888), .QN(n3323) );
  INVX0 U33296 ( .IN(n13579), .QN(n3331) );
  INVX0 U33297 ( .IN(n11413), .QN(n3267) );
  INVX0 U33298 ( .IN(n13270), .QN(n3339) );
  INVX0 U33299 ( .IN(n12961), .QN(n3347) );
  INVX0 U33300 ( .IN(n11104), .QN(n3275) );
  INVX0 U33301 ( .IN(n10794), .QN(n3283) );
  INVX0 U33302 ( .IN(n12652), .QN(n3355) );
  INVX0 U33303 ( .IN(n12343), .QN(n3363) );
  INVX0 U33304 ( .IN(n10485), .QN(n3291) );
  INVX0 U33305 ( .IN(n10175), .QN(n3299) );
  INVX0 U33306 ( .IN(n12033), .QN(n3371) );
  INVX0 U33307 ( .IN(n11723), .QN(n3379) );
  INVX0 U33308 ( .IN(n9865), .QN(n3307) );
  INVX0 U33309 ( .IN(n9554), .QN(n3315) );
  INVX0 U33310 ( .IN(n14162), .QN(n3255) );
  INVX0 U33311 ( .IN(n13775), .QN(n3431) );
  INVX0 U33312 ( .IN(n13466), .QN(n3435) );
  INVX0 U33313 ( .IN(n11300), .QN(n3403) );
  INVX0 U33314 ( .IN(n13157), .QN(n3439) );
  INVX0 U33315 ( .IN(n12848), .QN(n3443) );
  INVX0 U33316 ( .IN(n10991), .QN(n3407) );
  INVX0 U33317 ( .IN(n10681), .QN(n3411) );
  INVX0 U33318 ( .IN(n12539), .QN(n3447) );
  INVX0 U33319 ( .IN(n12230), .QN(n3451) );
  INVX0 U33320 ( .IN(n10372), .QN(n3415) );
  INVX0 U33321 ( .IN(n10062), .QN(n3419) );
  INVX0 U33322 ( .IN(n11920), .QN(n3455) );
  INVX0 U33323 ( .IN(n11610), .QN(n3459) );
  INVX0 U33324 ( .IN(n9752), .QN(n3423) );
  INVX0 U33325 ( .IN(n9441), .QN(n3427) );
  INVX0 U33326 ( .IN(n14039), .QN(n3398) );
  INVX0 U33327 ( .IN(n13907), .QN(n3146) );
  INVX0 U33328 ( .IN(n13598), .QN(n3152) );
  INVX0 U33329 ( .IN(n11432), .QN(n3104) );
  INVX0 U33330 ( .IN(n13289), .QN(n3158) );
  INVX0 U33331 ( .IN(n12980), .QN(n3164) );
  INVX0 U33332 ( .IN(n11123), .QN(n3110) );
  INVX0 U33333 ( .IN(n10813), .QN(n3116) );
  INVX0 U33334 ( .IN(n12671), .QN(n3170) );
  INVX0 U33335 ( .IN(n12362), .QN(n3176) );
  INVX0 U33336 ( .IN(n10504), .QN(n3122) );
  INVX0 U33337 ( .IN(n10194), .QN(n3128) );
  INVX0 U33338 ( .IN(n12052), .QN(n3182) );
  INVX0 U33339 ( .IN(n11742), .QN(n3188) );
  INVX0 U33340 ( .IN(n9884), .QN(n3134) );
  INVX0 U33341 ( .IN(n9573), .QN(n3140) );
  INVX0 U33342 ( .IN(n14181), .QN(n3094) );
  INVX0 U33343 ( .IN(n13818), .QN(n3322) );
  INVX0 U33344 ( .IN(n13509), .QN(n3330) );
  INVX0 U33345 ( .IN(n11343), .QN(n3266) );
  INVX0 U33346 ( .IN(n13200), .QN(n3338) );
  INVX0 U33347 ( .IN(n12891), .QN(n3346) );
  INVX0 U33348 ( .IN(n11034), .QN(n3274) );
  INVX0 U33349 ( .IN(n10724), .QN(n3282) );
  INVX0 U33350 ( .IN(n12582), .QN(n3354) );
  INVX0 U33351 ( .IN(n12273), .QN(n3362) );
  INVX0 U33352 ( .IN(n10415), .QN(n3290) );
  INVX0 U33353 ( .IN(n10105), .QN(n3298) );
  INVX0 U33354 ( .IN(n11963), .QN(n3370) );
  INVX0 U33355 ( .IN(n11653), .QN(n3378) );
  INVX0 U33356 ( .IN(n9795), .QN(n3306) );
  INVX0 U33357 ( .IN(n9484), .QN(n3314) );
  INVX0 U33358 ( .IN(n13950), .QN(n3258) );
  INVX0 U33359 ( .IN(n13835), .QN(n3144) );
  INVX0 U33360 ( .IN(n13526), .QN(n3150) );
  INVX0 U33361 ( .IN(n11360), .QN(n3102) );
  INVX0 U33362 ( .IN(n13217), .QN(n3156) );
  INVX0 U33363 ( .IN(n12908), .QN(n3162) );
  INVX0 U33364 ( .IN(n11051), .QN(n3108) );
  INVX0 U33365 ( .IN(n10741), .QN(n3114) );
  INVX0 U33366 ( .IN(n12599), .QN(n3168) );
  INVX0 U33367 ( .IN(n12290), .QN(n3174) );
  INVX0 U33368 ( .IN(n10432), .QN(n3120) );
  INVX0 U33369 ( .IN(n10122), .QN(n3126) );
  INVX0 U33370 ( .IN(n11980), .QN(n3180) );
  INVX0 U33371 ( .IN(n11670), .QN(n3186) );
  INVX0 U33372 ( .IN(n9812), .QN(n3132) );
  INVX0 U33373 ( .IN(n9501), .QN(n3138) );
  INVX0 U33374 ( .IN(n13968), .QN(n3095) );
  INVX0 U33375 ( .IN(n13445), .QN(n3328) );
  INVX0 U33376 ( .IN(n10970), .QN(n3272) );
  INVX0 U33377 ( .IN(n10351), .QN(n3288) );
  INVX0 U33378 ( .IN(n9731), .QN(n3304) );
  INVX0 U33379 ( .IN(n13832), .QN(n3223) );
  INVX0 U33380 ( .IN(n13523), .QN(n3227) );
  INVX0 U33381 ( .IN(n11357), .QN(n3195) );
  INVX0 U33382 ( .IN(n13214), .QN(n3231) );
  INVX0 U33383 ( .IN(n12905), .QN(n3235) );
  INVX0 U33384 ( .IN(n11048), .QN(n3199) );
  INVX0 U33385 ( .IN(n10738), .QN(n3203) );
  INVX0 U33386 ( .IN(n12596), .QN(n3239) );
  INVX0 U33387 ( .IN(n12287), .QN(n3243) );
  INVX0 U33388 ( .IN(n10429), .QN(n3207) );
  INVX0 U33389 ( .IN(n10119), .QN(n3211) );
  INVX0 U33390 ( .IN(n11977), .QN(n3247) );
  INVX0 U33391 ( .IN(n11667), .QN(n3251) );
  INVX0 U33392 ( .IN(n9809), .QN(n3215) );
  INVX0 U33393 ( .IN(n9498), .QN(n3219) );
  INVX0 U33394 ( .IN(n13965), .QN(n3191) );
  INVX0 U33395 ( .IN(n13674), .QN(n3318) );
  INVX0 U33396 ( .IN(n13365), .QN(n3326) );
  INVX0 U33397 ( .IN(n11199), .QN(n3262) );
  INVX0 U33398 ( .IN(n13056), .QN(n3334) );
  INVX0 U33399 ( .IN(n12747), .QN(n3342) );
  INVX0 U33400 ( .IN(n10890), .QN(n3270) );
  INVX0 U33401 ( .IN(n10580), .QN(n3278) );
  INVX0 U33402 ( .IN(n12438), .QN(n3350) );
  INVX0 U33403 ( .IN(n12129), .QN(n3358) );
  INVX0 U33404 ( .IN(n10271), .QN(n3286) );
  INVX0 U33405 ( .IN(n9961), .QN(n3294) );
  INVX0 U33406 ( .IN(n11819), .QN(n3366) );
  INVX0 U33407 ( .IN(n11509), .QN(n3374) );
  INVX0 U33408 ( .IN(n9651), .QN(n3302) );
  INVX0 U33409 ( .IN(n9340), .QN(n3310) );
  INVX0 U33410 ( .IN(n14090), .QN(n3260) );
  INVX0 U33411 ( .IN(n13448), .QN(n3809) );
  INVX0 U33412 ( .IN(n10973), .QN(n4124) );
  INVX0 U33413 ( .IN(n10354), .QN(n4034) );
  INVX0 U33414 ( .IN(n9734), .QN(n3944) );
  INVX0 U33415 ( .IN(n13757), .QN(n3854) );
  INVX0 U33416 ( .IN(n11282), .QN(n4169) );
  INVX0 U33417 ( .IN(n13139), .QN(n3764) );
  INVX0 U33418 ( .IN(n12830), .QN(n3719) );
  INVX0 U33419 ( .IN(n10663), .QN(n4079) );
  INVX0 U33420 ( .IN(n12521), .QN(n3674) );
  INVX0 U33421 ( .IN(n12212), .QN(n3629) );
  INVX0 U33422 ( .IN(n10044), .QN(n3989) );
  INVX0 U33423 ( .IN(n11902), .QN(n3584) );
  INVX0 U33424 ( .IN(n11592), .QN(n3539) );
  INVX0 U33425 ( .IN(n9423), .QN(n3899) );
  INVX0 U33426 ( .IN(n14021), .QN(n4214) );
  INVX0 U33427 ( .IN(n13675), .QN(n3141) );
  INVX0 U33428 ( .IN(n13366), .QN(n3147) );
  INVX0 U33429 ( .IN(n11200), .QN(n3099) );
  INVX0 U33430 ( .IN(n13057), .QN(n3153) );
  INVX0 U33431 ( .IN(n12748), .QN(n3159) );
  INVX0 U33432 ( .IN(n10891), .QN(n3105) );
  INVX0 U33433 ( .IN(n10581), .QN(n3111) );
  INVX0 U33434 ( .IN(n12439), .QN(n3165) );
  INVX0 U33435 ( .IN(n12130), .QN(n3171) );
  INVX0 U33436 ( .IN(n10272), .QN(n3117) );
  INVX0 U33437 ( .IN(n9962), .QN(n3123) );
  INVX0 U33438 ( .IN(n11820), .QN(n3177) );
  INVX0 U33439 ( .IN(n11510), .QN(n3183) );
  INVX0 U33440 ( .IN(n9652), .QN(n3129) );
  INVX0 U33441 ( .IN(n9341), .QN(n3135) );
  INVX0 U33442 ( .IN(n14108), .QN(n3097) );
  INVX0 U33443 ( .IN(n11279), .QN(n3264) );
  INVX0 U33444 ( .IN(n10660), .QN(n3280) );
  INVX0 U33445 ( .IN(n10041), .QN(n3296) );
  INVX0 U33446 ( .IN(n9420), .QN(n3312) );
  INVX0 U33447 ( .IN(n13754), .QN(n3320) );
  INVX0 U33448 ( .IN(n13136), .QN(n3336) );
  INVX0 U33449 ( .IN(n12827), .QN(n3344) );
  INVX0 U33450 ( .IN(n12518), .QN(n3352) );
  INVX0 U33451 ( .IN(n12209), .QN(n3360) );
  INVX0 U33452 ( .IN(n11899), .QN(n3368) );
  INVX0 U33453 ( .IN(n11589), .QN(n3376) );
  INVX0 U33454 ( .IN(n14018), .QN(n3254) );
  INVX0 U33455 ( .IN(n13673), .QN(n3221) );
  INVX0 U33456 ( .IN(n13364), .QN(n3225) );
  INVX0 U33457 ( .IN(n11198), .QN(n3193) );
  INVX0 U33458 ( .IN(n13055), .QN(n3229) );
  INVX0 U33459 ( .IN(n12746), .QN(n3233) );
  INVX0 U33460 ( .IN(n10889), .QN(n3197) );
  INVX0 U33461 ( .IN(n10579), .QN(n3201) );
  INVX0 U33462 ( .IN(n12437), .QN(n3237) );
  INVX0 U33463 ( .IN(n12128), .QN(n3241) );
  INVX0 U33464 ( .IN(n10270), .QN(n3205) );
  INVX0 U33465 ( .IN(n9960), .QN(n3209) );
  INVX0 U33466 ( .IN(n11818), .QN(n3245) );
  INVX0 U33467 ( .IN(n11508), .QN(n3249) );
  INVX0 U33468 ( .IN(n9650), .QN(n3213) );
  INVX0 U33469 ( .IN(n9339), .QN(n3217) );
  INVX0 U33470 ( .IN(n14105), .QN(n3192) );
  INVX0 U33471 ( .IN(n13463), .QN(n3149) );
  INVX0 U33472 ( .IN(n10988), .QN(n3107) );
  INVX0 U33473 ( .IN(n10369), .QN(n3119) );
  INVX0 U33474 ( .IN(n9749), .QN(n3131) );
  INVX0 U33475 ( .IN(n13772), .QN(n3143) );
  INVX0 U33476 ( .IN(n11297), .QN(n3101) );
  INVX0 U33477 ( .IN(n13154), .QN(n3155) );
  INVX0 U33478 ( .IN(n12845), .QN(n3161) );
  INVX0 U33479 ( .IN(n10678), .QN(n3113) );
  INVX0 U33480 ( .IN(n12536), .QN(n3167) );
  INVX0 U33481 ( .IN(n12227), .QN(n3173) );
  INVX0 U33482 ( .IN(n10059), .QN(n3125) );
  INVX0 U33483 ( .IN(n11917), .QN(n3179) );
  INVX0 U33484 ( .IN(n11607), .QN(n3185) );
  INVX0 U33485 ( .IN(n9438), .QN(n3137) );
  INVX0 U33486 ( .IN(n14036), .QN(n3093) );
  INVX0 U33487 ( .IN(n13758), .QN(n3858) );
  INVX0 U33488 ( .IN(n13449), .QN(n3813) );
  INVX0 U33489 ( .IN(n11283), .QN(n4173) );
  INVX0 U33490 ( .IN(n13140), .QN(n3768) );
  INVX0 U33491 ( .IN(n12831), .QN(n3723) );
  INVX0 U33492 ( .IN(n10974), .QN(n4128) );
  INVX0 U33493 ( .IN(n10664), .QN(n4083) );
  INVX0 U33494 ( .IN(n12522), .QN(n3678) );
  INVX0 U33495 ( .IN(n12213), .QN(n3633) );
  INVX0 U33496 ( .IN(n10355), .QN(n4038) );
  INVX0 U33497 ( .IN(n10045), .QN(n3993) );
  INVX0 U33498 ( .IN(n11903), .QN(n3588) );
  INVX0 U33499 ( .IN(n11593), .QN(n3543) );
  INVX0 U33500 ( .IN(n9735), .QN(n3948) );
  INVX0 U33501 ( .IN(n9424), .QN(n3903) );
  INVX0 U33502 ( .IN(n14022), .QN(n4218) );
  INVX0 U33503 ( .IN(n13876), .QN(n3497) );
  INVX0 U33504 ( .IN(n13567), .QN(n3501) );
  INVX0 U33505 ( .IN(n11401), .QN(n3469) );
  INVX0 U33506 ( .IN(n13258), .QN(n3505) );
  INVX0 U33507 ( .IN(n12949), .QN(n3509) );
  INVX0 U33508 ( .IN(n11092), .QN(n3473) );
  INVX0 U33509 ( .IN(n10782), .QN(n3477) );
  INVX0 U33510 ( .IN(n12640), .QN(n3513) );
  INVX0 U33511 ( .IN(n12331), .QN(n3517) );
  INVX0 U33512 ( .IN(n10473), .QN(n3481) );
  INVX0 U33513 ( .IN(n10163), .QN(n3485) );
  INVX0 U33514 ( .IN(n12021), .QN(n3521) );
  INVX0 U33515 ( .IN(n11711), .QN(n3525) );
  INVX0 U33516 ( .IN(n9853), .QN(n3489) );
  INVX0 U33517 ( .IN(n9542), .QN(n3493) );
  INVX0 U33518 ( .IN(n14150), .QN(n3463) );
  INVX0 U33519 ( .IN(n13473), .QN(n3812) );
  INVX0 U33520 ( .IN(n10998), .QN(n4127) );
  INVX0 U33521 ( .IN(n10379), .QN(n4037) );
  INVX0 U33522 ( .IN(n9759), .QN(n3947) );
  INVX0 U33523 ( .IN(n13782), .QN(n3857) );
  INVX0 U33524 ( .IN(n11307), .QN(n4172) );
  INVX0 U33525 ( .IN(n13164), .QN(n3767) );
  INVX0 U33526 ( .IN(n12855), .QN(n3722) );
  INVX0 U33527 ( .IN(n10688), .QN(n4082) );
  INVX0 U33528 ( .IN(n12546), .QN(n3677) );
  INVX0 U33529 ( .IN(n12237), .QN(n3632) );
  INVX0 U33530 ( .IN(n10069), .QN(n3992) );
  INVX0 U33531 ( .IN(n11927), .QN(n3587) );
  INVX0 U33532 ( .IN(n11617), .QN(n3542) );
  INVX0 U33533 ( .IN(n9448), .QN(n3902) );
  INVX0 U33534 ( .IN(n14046), .QN(n4217) );
  INVX0 U33535 ( .IN(n13911), .QN(n3881) );
  INVX0 U33536 ( .IN(n13602), .QN(n3836) );
  INVX0 U33537 ( .IN(n11436), .QN(n4196) );
  INVX0 U33538 ( .IN(n13293), .QN(n3791) );
  INVX0 U33539 ( .IN(n12984), .QN(n3746) );
  INVX0 U33540 ( .IN(n11127), .QN(n4151) );
  INVX0 U33541 ( .IN(n10817), .QN(n4106) );
  INVX0 U33542 ( .IN(n12675), .QN(n3701) );
  INVX0 U33543 ( .IN(n12366), .QN(n3656) );
  INVX0 U33544 ( .IN(n10508), .QN(n4061) );
  INVX0 U33545 ( .IN(n10198), .QN(n4016) );
  INVX0 U33546 ( .IN(n12056), .QN(n3611) );
  INVX0 U33547 ( .IN(n11746), .QN(n3566) );
  INVX0 U33548 ( .IN(n9888), .QN(n3971) );
  INVX0 U33549 ( .IN(n9577), .QN(n3926) );
  INVX0 U33550 ( .IN(n14185), .QN(n4241) );
  INVX0 U33551 ( .IN(n13844), .QN(n3865) );
  INVX0 U33552 ( .IN(n13715), .QN(n3873) );
  INVX0 U33553 ( .IN(n13535), .QN(n3820) );
  INVX0 U33554 ( .IN(n13406), .QN(n3828) );
  INVX0 U33555 ( .IN(n11369), .QN(n4180) );
  INVX0 U33556 ( .IN(n11240), .QN(n4188) );
  INVX0 U33557 ( .IN(n13226), .QN(n3775) );
  INVX0 U33558 ( .IN(n13097), .QN(n3783) );
  INVX0 U33559 ( .IN(n12917), .QN(n3730) );
  INVX0 U33560 ( .IN(n12788), .QN(n3738) );
  INVX0 U33561 ( .IN(n11060), .QN(n4135) );
  INVX0 U33562 ( .IN(n10931), .QN(n4143) );
  INVX0 U33563 ( .IN(n10750), .QN(n4090) );
  INVX0 U33564 ( .IN(n10621), .QN(n4098) );
  INVX0 U33565 ( .IN(n12608), .QN(n3685) );
  INVX0 U33566 ( .IN(n12479), .QN(n3693) );
  INVX0 U33567 ( .IN(n12299), .QN(n3640) );
  INVX0 U33568 ( .IN(n12170), .QN(n3648) );
  INVX0 U33569 ( .IN(n10441), .QN(n4045) );
  INVX0 U33570 ( .IN(n10312), .QN(n4053) );
  INVX0 U33571 ( .IN(n10131), .QN(n4000) );
  INVX0 U33572 ( .IN(n10002), .QN(n4008) );
  INVX0 U33573 ( .IN(n11989), .QN(n3595) );
  INVX0 U33574 ( .IN(n11860), .QN(n3603) );
  INVX0 U33575 ( .IN(n11679), .QN(n3550) );
  INVX0 U33576 ( .IN(n11550), .QN(n3558) );
  INVX0 U33577 ( .IN(n9821), .QN(n3955) );
  INVX0 U33578 ( .IN(n9692), .QN(n3963) );
  INVX0 U33579 ( .IN(n9510), .QN(n3910) );
  INVX0 U33580 ( .IN(n9381), .QN(n3918) );
  INVX0 U33581 ( .IN(n13977), .QN(n4225) );
  INVX0 U33582 ( .IN(n14117), .QN(n4233) );
  INVX0 U33583 ( .IN(n13769), .QN(n3222) );
  INVX0 U33584 ( .IN(n13460), .QN(n3226) );
  INVX0 U33585 ( .IN(n11294), .QN(n3194) );
  INVX0 U33586 ( .IN(n13151), .QN(n3230) );
  INVX0 U33587 ( .IN(n12842), .QN(n3234) );
  INVX0 U33588 ( .IN(n10985), .QN(n3198) );
  INVX0 U33589 ( .IN(n10675), .QN(n3202) );
  INVX0 U33590 ( .IN(n12533), .QN(n3238) );
  INVX0 U33591 ( .IN(n12224), .QN(n3242) );
  INVX0 U33592 ( .IN(n10366), .QN(n3206) );
  INVX0 U33593 ( .IN(n10056), .QN(n3210) );
  INVX0 U33594 ( .IN(n11914), .QN(n3246) );
  INVX0 U33595 ( .IN(n11604), .QN(n3250) );
  INVX0 U33596 ( .IN(n9746), .QN(n3214) );
  INVX0 U33597 ( .IN(n9435), .QN(n3218) );
  INVX0 U33598 ( .IN(n14033), .QN(n3189) );
  INVX0 U33599 ( .IN(n13863), .QN(n3862) );
  INVX0 U33600 ( .IN(n13732), .QN(n3870) );
  INVX0 U33601 ( .IN(n13554), .QN(n3817) );
  INVX0 U33602 ( .IN(n13423), .QN(n3825) );
  INVX0 U33603 ( .IN(n11388), .QN(n4177) );
  INVX0 U33604 ( .IN(n11257), .QN(n4185) );
  INVX0 U33605 ( .IN(n13245), .QN(n3772) );
  INVX0 U33606 ( .IN(n13114), .QN(n3780) );
  INVX0 U33607 ( .IN(n12936), .QN(n3727) );
  INVX0 U33608 ( .IN(n12805), .QN(n3735) );
  INVX0 U33609 ( .IN(n11079), .QN(n4132) );
  INVX0 U33610 ( .IN(n10948), .QN(n4140) );
  INVX0 U33611 ( .IN(n10769), .QN(n4087) );
  INVX0 U33612 ( .IN(n10638), .QN(n4095) );
  INVX0 U33613 ( .IN(n12627), .QN(n3682) );
  INVX0 U33614 ( .IN(n12496), .QN(n3690) );
  INVX0 U33615 ( .IN(n12318), .QN(n3637) );
  INVX0 U33616 ( .IN(n12187), .QN(n3645) );
  INVX0 U33617 ( .IN(n10460), .QN(n4042) );
  INVX0 U33618 ( .IN(n10329), .QN(n4050) );
  INVX0 U33619 ( .IN(n10150), .QN(n3997) );
  INVX0 U33620 ( .IN(n10019), .QN(n4005) );
  INVX0 U33621 ( .IN(n12008), .QN(n3592) );
  INVX0 U33622 ( .IN(n11877), .QN(n3600) );
  INVX0 U33623 ( .IN(n11698), .QN(n3547) );
  INVX0 U33624 ( .IN(n11567), .QN(n3555) );
  INVX0 U33625 ( .IN(n9840), .QN(n3952) );
  INVX0 U33626 ( .IN(n9709), .QN(n3960) );
  INVX0 U33627 ( .IN(n9529), .QN(n3907) );
  INVX0 U33628 ( .IN(n9398), .QN(n3915) );
  INVX0 U33629 ( .IN(n13996), .QN(n4222) );
  INVX0 U33630 ( .IN(n14136), .QN(n4230) );
  INVX0 U33631 ( .IN(n11277), .QN(n4170) );
  INVX0 U33632 ( .IN(n10658), .QN(n4080) );
  INVX0 U33633 ( .IN(n10039), .QN(n3990) );
  INVX0 U33634 ( .IN(n9418), .QN(n3900) );
  INVX0 U33635 ( .IN(n13885), .QN(n3879) );
  INVX0 U33636 ( .IN(n13576), .QN(n3834) );
  INVX0 U33637 ( .IN(n11410), .QN(n4194) );
  INVX0 U33638 ( .IN(n13267), .QN(n3789) );
  INVX0 U33639 ( .IN(n12958), .QN(n3744) );
  INVX0 U33640 ( .IN(n11101), .QN(n4149) );
  INVX0 U33641 ( .IN(n10791), .QN(n4104) );
  INVX0 U33642 ( .IN(n12649), .QN(n3699) );
  INVX0 U33643 ( .IN(n12340), .QN(n3654) );
  INVX0 U33644 ( .IN(n10482), .QN(n4059) );
  INVX0 U33645 ( .IN(n10172), .QN(n4014) );
  INVX0 U33646 ( .IN(n12030), .QN(n3609) );
  INVX0 U33647 ( .IN(n11720), .QN(n3564) );
  INVX0 U33648 ( .IN(n9862), .QN(n3969) );
  INVX0 U33649 ( .IN(n9551), .QN(n3924) );
  INVX0 U33650 ( .IN(n14159), .QN(n4239) );
  INVX0 U33651 ( .IN(n13752), .QN(n3855) );
  INVX0 U33652 ( .IN(n13134), .QN(n3765) );
  INVX0 U33653 ( .IN(n12825), .QN(n3720) );
  INVX0 U33654 ( .IN(n12516), .QN(n3675) );
  INVX0 U33655 ( .IN(n12207), .QN(n3630) );
  INVX0 U33656 ( .IN(n11897), .QN(n3585) );
  INVX0 U33657 ( .IN(n11587), .QN(n3540) );
  INVX0 U33658 ( .IN(n14016), .QN(n4215) );
  INVX0 U33659 ( .IN(n13443), .QN(n3810) );
  INVX0 U33660 ( .IN(n10968), .QN(n4125) );
  INVX0 U33661 ( .IN(n10349), .QN(n4035) );
  INVX0 U33662 ( .IN(n9729), .QN(n3945) );
  INVX0 U33663 ( .IN(n13929), .QN(n3878) );
  INVX0 U33664 ( .IN(n13620), .QN(n3833) );
  INVX0 U33665 ( .IN(n11454), .QN(n4193) );
  INVX0 U33666 ( .IN(n13311), .QN(n3788) );
  INVX0 U33667 ( .IN(n13002), .QN(n3743) );
  INVX0 U33668 ( .IN(n11145), .QN(n4148) );
  INVX0 U33669 ( .IN(n10835), .QN(n4103) );
  INVX0 U33670 ( .IN(n12693), .QN(n3698) );
  INVX0 U33671 ( .IN(n12384), .QN(n3653) );
  INVX0 U33672 ( .IN(n10526), .QN(n4058) );
  INVX0 U33673 ( .IN(n10216), .QN(n4013) );
  INVX0 U33674 ( .IN(n12074), .QN(n3608) );
  INVX0 U33675 ( .IN(n11764), .QN(n3563) );
  INVX0 U33676 ( .IN(n9906), .QN(n3968) );
  INVX0 U33677 ( .IN(n9595), .QN(n3923) );
  INVX0 U33678 ( .IN(n14203), .QN(n4238) );
  INVX0 U33679 ( .IN(n13948), .QN(n4223) );
  INVX0 U33680 ( .IN(n14088), .QN(n4231) );
  INVX0 U33681 ( .IN(n13928), .QN(n2979) );
  INVX0 U33682 ( .IN(n13619), .QN(n2995) );
  INVX0 U33683 ( .IN(n11453), .QN(n2867) );
  INVX0 U33684 ( .IN(n13310), .QN(n3011) );
  INVX0 U33685 ( .IN(n13001), .QN(n3027) );
  INVX0 U33686 ( .IN(n11144), .QN(n2883) );
  INVX0 U33687 ( .IN(n10834), .QN(n2899) );
  INVX0 U33688 ( .IN(n12692), .QN(n3043) );
  INVX0 U33689 ( .IN(n12383), .QN(n3059) );
  INVX0 U33690 ( .IN(n10525), .QN(n2915) );
  INVX0 U33691 ( .IN(n10215), .QN(n2931) );
  INVX0 U33692 ( .IN(n12073), .QN(n3075) );
  INVX0 U33693 ( .IN(n11763), .QN(n3091) );
  INVX0 U33694 ( .IN(n9905), .QN(n2947) );
  INVX0 U33695 ( .IN(n9594), .QN(n2963) );
  INVX0 U33696 ( .IN(n14202), .QN(n2842) );
  INVX0 U33697 ( .IN(n13816), .QN(n3863) );
  INVX0 U33698 ( .IN(n13691), .QN(n3871) );
  INVX0 U33699 ( .IN(n13507), .QN(n3818) );
  INVX0 U33700 ( .IN(n13382), .QN(n3826) );
  INVX0 U33701 ( .IN(n11341), .QN(n4178) );
  INVX0 U33702 ( .IN(n11216), .QN(n4186) );
  INVX0 U33703 ( .IN(n13198), .QN(n3773) );
  INVX0 U33704 ( .IN(n13073), .QN(n3781) );
  INVX0 U33705 ( .IN(n12889), .QN(n3728) );
  INVX0 U33706 ( .IN(n12764), .QN(n3736) );
  INVX0 U33707 ( .IN(n11032), .QN(n4133) );
  INVX0 U33708 ( .IN(n10907), .QN(n4141) );
  INVX0 U33709 ( .IN(n10722), .QN(n4088) );
  INVX0 U33710 ( .IN(n10597), .QN(n4096) );
  INVX0 U33711 ( .IN(n12580), .QN(n3683) );
  INVX0 U33712 ( .IN(n12455), .QN(n3691) );
  INVX0 U33713 ( .IN(n12271), .QN(n3638) );
  INVX0 U33714 ( .IN(n12146), .QN(n3646) );
  INVX0 U33715 ( .IN(n10413), .QN(n4043) );
  INVX0 U33716 ( .IN(n10288), .QN(n4051) );
  INVX0 U33717 ( .IN(n10103), .QN(n3998) );
  INVX0 U33718 ( .IN(n9978), .QN(n4006) );
  INVX0 U33719 ( .IN(n11961), .QN(n3593) );
  INVX0 U33720 ( .IN(n11836), .QN(n3601) );
  INVX0 U33721 ( .IN(n11651), .QN(n3548) );
  INVX0 U33722 ( .IN(n11526), .QN(n3556) );
  INVX0 U33723 ( .IN(n9793), .QN(n3953) );
  INVX0 U33724 ( .IN(n9668), .QN(n3961) );
  INVX0 U33725 ( .IN(n9482), .QN(n3908) );
  INVX0 U33726 ( .IN(n9357), .QN(n3916) );
  INVX0 U33727 ( .IN(n13847), .QN(n2974) );
  INVX0 U33728 ( .IN(n13538), .QN(n2990) );
  INVX0 U33729 ( .IN(n11372), .QN(n2862) );
  INVX0 U33730 ( .IN(n13229), .QN(n3006) );
  INVX0 U33731 ( .IN(n12920), .QN(n3022) );
  INVX0 U33732 ( .IN(n11063), .QN(n2878) );
  INVX0 U33733 ( .IN(n10753), .QN(n2894) );
  INVX0 U33734 ( .IN(n12611), .QN(n3038) );
  INVX0 U33735 ( .IN(n12302), .QN(n3054) );
  INVX0 U33736 ( .IN(n10444), .QN(n2910) );
  INVX0 U33737 ( .IN(n10134), .QN(n2926) );
  INVX0 U33738 ( .IN(n11992), .QN(n3070) );
  INVX0 U33739 ( .IN(n11682), .QN(n3086) );
  INVX0 U33740 ( .IN(n9824), .QN(n2942) );
  INVX0 U33741 ( .IN(n9513), .QN(n2958) );
  INVX0 U33742 ( .IN(n13980), .QN(n2844) );
  INVX0 U33743 ( .IN(n13850), .QN(n3866) );
  INVX0 U33744 ( .IN(n13720), .QN(n3874) );
  INVX0 U33745 ( .IN(n13541), .QN(n3821) );
  INVX0 U33746 ( .IN(n13411), .QN(n3829) );
  INVX0 U33747 ( .IN(n11375), .QN(n4181) );
  INVX0 U33748 ( .IN(n11245), .QN(n4189) );
  INVX0 U33749 ( .IN(n13232), .QN(n3776) );
  INVX0 U33750 ( .IN(n13102), .QN(n3784) );
  INVX0 U33751 ( .IN(n12923), .QN(n3731) );
  INVX0 U33752 ( .IN(n12793), .QN(n3739) );
  INVX0 U33753 ( .IN(n11066), .QN(n4136) );
  INVX0 U33754 ( .IN(n10936), .QN(n4144) );
  INVX0 U33755 ( .IN(n10756), .QN(n4091) );
  INVX0 U33756 ( .IN(n10626), .QN(n4099) );
  INVX0 U33757 ( .IN(n12614), .QN(n3686) );
  INVX0 U33758 ( .IN(n12484), .QN(n3694) );
  INVX0 U33759 ( .IN(n12305), .QN(n3641) );
  INVX0 U33760 ( .IN(n12175), .QN(n3649) );
  INVX0 U33761 ( .IN(n10447), .QN(n4046) );
  INVX0 U33762 ( .IN(n10317), .QN(n4054) );
  INVX0 U33763 ( .IN(n10137), .QN(n4001) );
  INVX0 U33764 ( .IN(n10007), .QN(n4009) );
  INVX0 U33765 ( .IN(n11995), .QN(n3596) );
  INVX0 U33766 ( .IN(n11865), .QN(n3604) );
  INVX0 U33767 ( .IN(n11685), .QN(n3551) );
  INVX0 U33768 ( .IN(n11555), .QN(n3559) );
  INVX0 U33769 ( .IN(n9827), .QN(n3956) );
  INVX0 U33770 ( .IN(n9697), .QN(n3964) );
  INVX0 U33771 ( .IN(n9516), .QN(n3911) );
  INVX0 U33772 ( .IN(n9386), .QN(n3919) );
  INVX0 U33773 ( .IN(n13983), .QN(n4226) );
  INVX0 U33774 ( .IN(n14123), .QN(n4234) );
  INVX0 U33775 ( .IN(n13917), .QN(n3882) );
  INVX0 U33776 ( .IN(n13608), .QN(n3837) );
  INVX0 U33777 ( .IN(n11442), .QN(n4197) );
  INVX0 U33778 ( .IN(n13299), .QN(n3792) );
  INVX0 U33779 ( .IN(n12990), .QN(n3747) );
  INVX0 U33780 ( .IN(n11133), .QN(n4152) );
  INVX0 U33781 ( .IN(n10823), .QN(n4107) );
  INVX0 U33782 ( .IN(n12681), .QN(n3702) );
  INVX0 U33783 ( .IN(n12372), .QN(n3657) );
  INVX0 U33784 ( .IN(n10514), .QN(n4062) );
  INVX0 U33785 ( .IN(n10204), .QN(n4017) );
  INVX0 U33786 ( .IN(n12062), .QN(n3612) );
  INVX0 U33787 ( .IN(n11752), .QN(n3567) );
  INVX0 U33788 ( .IN(n9894), .QN(n3972) );
  INVX0 U33789 ( .IN(n9583), .QN(n3927) );
  INVX0 U33790 ( .IN(n14191), .QN(n4242) );
  INVX0 U33791 ( .IN(n13987), .QN(n3464) );
  INVX0 U33792 ( .IN(n14120), .QN(n2849) );
  INVX0 U33793 ( .IN(n13854), .QN(n3496) );
  INVX0 U33794 ( .IN(n13545), .QN(n3500) );
  INVX0 U33795 ( .IN(n11379), .QN(n3468) );
  INVX0 U33796 ( .IN(n13236), .QN(n3504) );
  INVX0 U33797 ( .IN(n12927), .QN(n3508) );
  INVX0 U33798 ( .IN(n11070), .QN(n3472) );
  INVX0 U33799 ( .IN(n10760), .QN(n3476) );
  INVX0 U33800 ( .IN(n12618), .QN(n3512) );
  INVX0 U33801 ( .IN(n12309), .QN(n3516) );
  INVX0 U33802 ( .IN(n10451), .QN(n3480) );
  INVX0 U33803 ( .IN(n10141), .QN(n3484) );
  INVX0 U33804 ( .IN(n11999), .QN(n3520) );
  INVX0 U33805 ( .IN(n11689), .QN(n3524) );
  INVX0 U33806 ( .IN(n9831), .QN(n3488) );
  INVX0 U33807 ( .IN(n9520), .QN(n3492) );
  INVX0 U33808 ( .IN(n13676), .QN(n2966) );
  INVX0 U33809 ( .IN(n13367), .QN(n2982) );
  INVX0 U33810 ( .IN(n11201), .QN(n2854) );
  INVX0 U33811 ( .IN(n13058), .QN(n2998) );
  INVX0 U33812 ( .IN(n12749), .QN(n3014) );
  INVX0 U33813 ( .IN(n10892), .QN(n2870) );
  INVX0 U33814 ( .IN(n10582), .QN(n2886) );
  INVX0 U33815 ( .IN(n12440), .QN(n3030) );
  INVX0 U33816 ( .IN(n12131), .QN(n3046) );
  INVX0 U33817 ( .IN(n10273), .QN(n2902) );
  INVX0 U33818 ( .IN(n9963), .QN(n2918) );
  INVX0 U33819 ( .IN(n11821), .QN(n3062) );
  INVX0 U33820 ( .IN(n11511), .QN(n3078) );
  INVX0 U33821 ( .IN(n9653), .QN(n2934) );
  INVX0 U33822 ( .IN(n9342), .QN(n2950) );
  INVX0 U33823 ( .IN(n13678), .QN(n3494) );
  INVX0 U33824 ( .IN(n13369), .QN(n3498) );
  INVX0 U33825 ( .IN(n11203), .QN(n3466) );
  INVX0 U33826 ( .IN(n13060), .QN(n3502) );
  INVX0 U33827 ( .IN(n12751), .QN(n3506) );
  INVX0 U33828 ( .IN(n10894), .QN(n3470) );
  INVX0 U33829 ( .IN(n10584), .QN(n3474) );
  INVX0 U33830 ( .IN(n12442), .QN(n3510) );
  INVX0 U33831 ( .IN(n12133), .QN(n3514) );
  INVX0 U33832 ( .IN(n10275), .QN(n3478) );
  INVX0 U33833 ( .IN(n9965), .QN(n3482) );
  INVX0 U33834 ( .IN(n11823), .QN(n3518) );
  INVX0 U33835 ( .IN(n11513), .QN(n3522) );
  INVX0 U33836 ( .IN(n9655), .QN(n3486) );
  INVX0 U33837 ( .IN(n9344), .QN(n3490) );
  INVX0 U33838 ( .IN(n14127), .QN(n3465) );
  INVX0 U33839 ( .IN(n13786), .QN(n2971) );
  INVX0 U33840 ( .IN(n13477), .QN(n2987) );
  INVX0 U33841 ( .IN(n11311), .QN(n2859) );
  INVX0 U33842 ( .IN(n13168), .QN(n3003) );
  INVX0 U33843 ( .IN(n12859), .QN(n3019) );
  INVX0 U33844 ( .IN(n11002), .QN(n2875) );
  INVX0 U33845 ( .IN(n10692), .QN(n2891) );
  INVX0 U33846 ( .IN(n12550), .QN(n3035) );
  INVX0 U33847 ( .IN(n12241), .QN(n3051) );
  INVX0 U33848 ( .IN(n10383), .QN(n2907) );
  INVX0 U33849 ( .IN(n10073), .QN(n2923) );
  INVX0 U33850 ( .IN(n11931), .QN(n3067) );
  INVX0 U33851 ( .IN(n11621), .QN(n3083) );
  INVX0 U33852 ( .IN(n9763), .QN(n2939) );
  INVX0 U33853 ( .IN(n9452), .QN(n2955) );
  INVX0 U33854 ( .IN(n14050), .QN(n2838) );
  INVX0 U33855 ( .IN(n13791), .QN(n3495) );
  INVX0 U33856 ( .IN(n13482), .QN(n3499) );
  INVX0 U33857 ( .IN(n11316), .QN(n3467) );
  INVX0 U33858 ( .IN(n13173), .QN(n3503) );
  INVX0 U33859 ( .IN(n12864), .QN(n3507) );
  INVX0 U33860 ( .IN(n11007), .QN(n3471) );
  INVX0 U33861 ( .IN(n10697), .QN(n3475) );
  INVX0 U33862 ( .IN(n12555), .QN(n3511) );
  INVX0 U33863 ( .IN(n12246), .QN(n3515) );
  INVX0 U33864 ( .IN(n10388), .QN(n3479) );
  INVX0 U33865 ( .IN(n10078), .QN(n3483) );
  INVX0 U33866 ( .IN(n11936), .QN(n3519) );
  INVX0 U33867 ( .IN(n11626), .QN(n3523) );
  INVX0 U33868 ( .IN(n9768), .QN(n3487) );
  INVX0 U33869 ( .IN(n9457), .QN(n3491) );
  INVX0 U33870 ( .IN(n14055), .QN(n3462) );
  AO22X1 U33871 ( .IN1(test_so67), .IN2(n13737), .IN3(n2970), .IN4(n13776), 
        .Q(n17583) );
  NAND3X0 U33872 ( .IN1(n13760), .IN2(n13777), .IN3(n13778), .QN(n13776) );
  OR2X1 U33873 ( .IN1(n3859), .IN2(n13743), .Q(n13777) );
  AO22X1 U33874 ( .IN1(s6_msel_gnt_p0[0]), .IN2(n13428), .IN3(n2986), .IN4(
        n13467), .Q(n17553) );
  NAND3X0 U33875 ( .IN1(n13451), .IN2(n13468), .IN3(n13469), .QN(n13467) );
  OR2X1 U33876 ( .IN1(n3814), .IN2(n13434), .Q(n13468) );
  OA221X1 U33877 ( .IN1(n3149), .IN2(n13470), .IN3(n13471), .IN4(n13472), 
        .IN5(n13431), .Q(n13469) );
  AO22X1 U33878 ( .IN1(s14_msel_gnt_p0_0_), .IN2(n11262), .IN3(n2858), .IN4(
        n11301), .Q(n17343) );
  NAND3X0 U33879 ( .IN1(n11285), .IN2(n11302), .IN3(n11303), .QN(n11301) );
  OR2X1 U33880 ( .IN1(n4174), .IN2(n11268), .Q(n11302) );
  AO22X1 U33881 ( .IN1(s5_msel_gnt_p0[0]), .IN2(n13119), .IN3(n3002), .IN4(
        n13158), .Q(n17523) );
  NAND3X0 U33882 ( .IN1(n13142), .IN2(n13159), .IN3(n13160), .QN(n13158) );
  OR2X1 U33883 ( .IN1(n3769), .IN2(n13125), .Q(n13159) );
  AO22X1 U33884 ( .IN1(s4_msel_gnt_p0[0]), .IN2(n12810), .IN3(n3018), .IN4(
        n12849), .Q(n17493) );
  NAND3X0 U33885 ( .IN1(n12833), .IN2(n12850), .IN3(n12851), .QN(n12849) );
  OR2X1 U33886 ( .IN1(n3724), .IN2(n12816), .Q(n12850) );
  AO22X1 U33887 ( .IN1(test_so90), .IN2(n10953), .IN3(n2874), .IN4(n10992), 
        .Q(n17313) );
  NAND3X0 U33888 ( .IN1(n10976), .IN2(n10993), .IN3(n10994), .QN(n10992) );
  OR2X1 U33889 ( .IN1(n4129), .IN2(n10959), .Q(n10993) );
  OA221X1 U33890 ( .IN1(n3107), .IN2(n10995), .IN3(n10996), .IN4(n10997), 
        .IN5(n10956), .Q(n10994) );
  AO22X1 U33891 ( .IN1(s12_msel_gnt_p0[0]), .IN2(n10643), .IN3(n2890), .IN4(
        n10682), .Q(n17283) );
  NAND3X0 U33892 ( .IN1(n10666), .IN2(n10683), .IN3(n10684), .QN(n10682) );
  OR2X1 U33893 ( .IN1(n4084), .IN2(n10649), .Q(n10683) );
  AO22X1 U33894 ( .IN1(s3_msel_gnt_p0_0_), .IN2(n12501), .IN3(n3034), .IN4(
        n12540), .Q(n17463) );
  NAND3X0 U33895 ( .IN1(n12524), .IN2(n12541), .IN3(n12542), .QN(n12540) );
  OR2X1 U33896 ( .IN1(n3679), .IN2(n12507), .Q(n12541) );
  AO22X1 U33897 ( .IN1(s2_msel_gnt_p0_0_), .IN2(n12192), .IN3(n3050), .IN4(
        n12231), .Q(n17433) );
  NAND3X0 U33898 ( .IN1(n12215), .IN2(n12232), .IN3(n12233), .QN(n12231) );
  OR2X1 U33899 ( .IN1(n3634), .IN2(n12198), .Q(n12232) );
  AO22X1 U33900 ( .IN1(s11_msel_gnt_p0[0]), .IN2(n10334), .IN3(n2906), .IN4(
        n10373), .Q(n17253) );
  NAND3X0 U33901 ( .IN1(n10357), .IN2(n10374), .IN3(n10375), .QN(n10373) );
  OR2X1 U33902 ( .IN1(n4039), .IN2(n10340), .Q(n10374) );
  OA221X1 U33903 ( .IN1(n3119), .IN2(n10376), .IN3(n10377), .IN4(n10378), 
        .IN5(n10337), .Q(n10375) );
  AO22X1 U33904 ( .IN1(s10_msel_gnt_p0[0]), .IN2(n10024), .IN3(n2922), .IN4(
        n10063), .Q(n17223) );
  NAND3X0 U33905 ( .IN1(n10047), .IN2(n10064), .IN3(n10065), .QN(n10063) );
  OR2X1 U33906 ( .IN1(n3994), .IN2(n10030), .Q(n10064) );
  AO22X1 U33907 ( .IN1(test_so44), .IN2(n11882), .IN3(n3066), .IN4(n11921), 
        .Q(n17403) );
  NAND3X0 U33908 ( .IN1(n11905), .IN2(n11922), .IN3(n11923), .QN(n11921) );
  OR2X1 U33909 ( .IN1(n3589), .IN2(n11888), .Q(n11922) );
  AO22X1 U33910 ( .IN1(s0_msel_gnt_p0[0]), .IN2(n11572), .IN3(n3082), .IN4(
        n11611), .Q(n17373) );
  NAND3X0 U33911 ( .IN1(n11595), .IN2(n11612), .IN3(n11613), .QN(n11611) );
  OR2X1 U33912 ( .IN1(n3544), .IN2(n11578), .Q(n11612) );
  AO22X1 U33913 ( .IN1(s9_msel_gnt_p0_0_), .IN2(n9714), .IN3(n2938), .IN4(
        n9753), .Q(n17193) );
  NAND3X0 U33914 ( .IN1(n9737), .IN2(n9754), .IN3(n9755), .QN(n9753) );
  OR2X1 U33915 ( .IN1(n3949), .IN2(n9720), .Q(n9754) );
  OA221X1 U33916 ( .IN1(n3131), .IN2(n9756), .IN3(n9757), .IN4(n9758), .IN5(
        n9717), .Q(n9755) );
  AO22X1 U33917 ( .IN1(s8_msel_gnt_p0_0_), .IN2(n9403), .IN3(n2954), .IN4(
        n9442), .Q(n17163) );
  NAND3X0 U33918 ( .IN1(n9426), .IN2(n9443), .IN3(n9444), .QN(n9442) );
  OR2X1 U33919 ( .IN1(n3904), .IN2(n9409), .Q(n9443) );
  OA221X1 U33920 ( .IN1(n13743), .IN2(n3861), .IN3(n13744), .IN4(n3495), .IN5(
        n13745), .Q(n13742) );
  ISOLANDX1 U33921 ( .D(n13746), .ISO(n13747), .Q(n13745) );
  OA221X1 U33922 ( .IN1(n13434), .IN2(n3816), .IN3(n13435), .IN4(n3499), .IN5(
        n13436), .Q(n13433) );
  ISOLANDX1 U33923 ( .D(n13437), .ISO(n13438), .Q(n13436) );
  OA221X1 U33924 ( .IN1(n11268), .IN2(n4176), .IN3(n11269), .IN4(n3467), .IN5(
        n11270), .Q(n11267) );
  ISOLANDX1 U33925 ( .D(n11271), .ISO(n11272), .Q(n11270) );
  OA221X1 U33926 ( .IN1(n13125), .IN2(n3771), .IN3(n13126), .IN4(n3503), .IN5(
        n13127), .Q(n13124) );
  ISOLANDX1 U33927 ( .D(n13128), .ISO(n13129), .Q(n13127) );
  OA221X1 U33928 ( .IN1(n12816), .IN2(n3726), .IN3(n12817), .IN4(n3507), .IN5(
        n12818), .Q(n12815) );
  ISOLANDX1 U33929 ( .D(n12819), .ISO(n12820), .Q(n12818) );
  OA221X1 U33930 ( .IN1(n10959), .IN2(n4131), .IN3(n10960), .IN4(n3471), .IN5(
        n10961), .Q(n10958) );
  ISOLANDX1 U33931 ( .D(n10962), .ISO(n10963), .Q(n10961) );
  OA221X1 U33932 ( .IN1(n10649), .IN2(n4086), .IN3(n10650), .IN4(n3475), .IN5(
        n10651), .Q(n10648) );
  ISOLANDX1 U33933 ( .D(n10652), .ISO(n10653), .Q(n10651) );
  OA221X1 U33934 ( .IN1(n12507), .IN2(n3681), .IN3(n12508), .IN4(n3511), .IN5(
        n12509), .Q(n12506) );
  ISOLANDX1 U33935 ( .D(n12510), .ISO(n12511), .Q(n12509) );
  OA221X1 U33936 ( .IN1(n12198), .IN2(n3636), .IN3(n12199), .IN4(n3515), .IN5(
        n12200), .Q(n12197) );
  ISOLANDX1 U33937 ( .D(n12201), .ISO(n12202), .Q(n12200) );
  OA221X1 U33938 ( .IN1(n10340), .IN2(n4041), .IN3(n10341), .IN4(n3479), .IN5(
        n10342), .Q(n10339) );
  ISOLANDX1 U33939 ( .D(n10343), .ISO(n10344), .Q(n10342) );
  OA221X1 U33940 ( .IN1(n10030), .IN2(n3996), .IN3(n10031), .IN4(n3483), .IN5(
        n10032), .Q(n10029) );
  ISOLANDX1 U33941 ( .D(n10033), .ISO(n10034), .Q(n10032) );
  OA221X1 U33942 ( .IN1(n11888), .IN2(n3591), .IN3(n11889), .IN4(n3519), .IN5(
        n11890), .Q(n11887) );
  ISOLANDX1 U33943 ( .D(n11891), .ISO(n11892), .Q(n11890) );
  OA221X1 U33944 ( .IN1(n11578), .IN2(n3546), .IN3(n11579), .IN4(n3523), .IN5(
        n11580), .Q(n11577) );
  ISOLANDX1 U33945 ( .D(n11581), .ISO(n11582), .Q(n11580) );
  OA221X1 U33946 ( .IN1(n9720), .IN2(n3951), .IN3(n9721), .IN4(n3487), .IN5(
        n9722), .Q(n9719) );
  ISOLANDX1 U33947 ( .D(n9723), .ISO(n9724), .Q(n9722) );
  OA221X1 U33948 ( .IN1(n9409), .IN2(n3906), .IN3(n9410), .IN4(n3491), .IN5(
        n9411), .Q(n9408) );
  ISOLANDX1 U33949 ( .D(n9412), .ISO(n9413), .Q(n9411) );
  OA221X1 U33950 ( .IN1(n14007), .IN2(n4221), .IN3(n14008), .IN4(n3462), .IN5(
        n14009), .Q(n14006) );
  ISOLANDX1 U33951 ( .D(n14010), .ISO(n14011), .Q(n14009) );
  AO22X1 U33952 ( .IN1(s7_msel_gnt_p0_1_), .IN2(n13737), .IN3(n2970), .IN4(
        n13759), .Q(n17582) );
  NAND3X0 U33953 ( .IN1(n13760), .IN2(n13746), .IN3(n13761), .QN(n13759) );
  OA222X1 U33954 ( .IN1(n13743), .IN2(n3860), .IN3(n13762), .IN4(n3431), .IN5(
        n13763), .IN6(n3222), .Q(n13761) );
  OA21X1 U33955 ( .IN1(n13764), .IN2(n13765), .IN3(n13766), .Q(n13763) );
  AO22X1 U33956 ( .IN1(s7_msel_gnt_p0_2_), .IN2(n13737), .IN3(n2970), .IN4(
        n13738), .Q(n17581) );
  NAND4X0 U33957 ( .IN1(n13739), .IN2(n13740), .IN3(n13741), .IN4(n13742), 
        .QN(n13738) );
  NAND3X0 U33958 ( .IN1(n13755), .IN2(n3320), .IN3(n13756), .QN(n13739) );
  AO22X1 U33959 ( .IN1(s6_msel_gnt_p0[1]), .IN2(n13428), .IN3(n2986), .IN4(
        n13450), .Q(n17552) );
  NAND3X0 U33960 ( .IN1(n13451), .IN2(n13437), .IN3(n13452), .QN(n13450) );
  OA222X1 U33961 ( .IN1(n13434), .IN2(n3815), .IN3(n13453), .IN4(n3435), .IN5(
        n13454), .IN6(n3226), .Q(n13452) );
  OA21X1 U33962 ( .IN1(n13444), .IN2(n13458), .IN3(n13459), .Q(n13453) );
  AO22X1 U33963 ( .IN1(s6_msel_gnt_p0[2]), .IN2(n13428), .IN3(n2986), .IN4(
        n13429), .Q(n17551) );
  NAND4X0 U33964 ( .IN1(n13430), .IN2(n13431), .IN3(n13432), .IN4(n13433), 
        .QN(n13429) );
  NAND3X0 U33965 ( .IN1(n13446), .IN2(n3328), .IN3(n13447), .QN(n13430) );
  OA22X1 U33966 ( .IN1(n13439), .IN2(n13440), .IN3(n13441), .IN4(n3435), .Q(
        n13432) );
  AO22X1 U33967 ( .IN1(test_so94), .IN2(n11262), .IN3(n2858), .IN4(n11284), 
        .Q(n17342) );
  NAND3X0 U33968 ( .IN1(n11285), .IN2(n11271), .IN3(n11286), .QN(n11284) );
  OA222X1 U33969 ( .IN1(n11268), .IN2(n4175), .IN3(n11287), .IN4(n3403), .IN5(
        n11288), .IN6(n3194), .Q(n11286) );
  OA21X1 U33970 ( .IN1(n11289), .IN2(n11290), .IN3(n11291), .Q(n11288) );
  AO22X1 U33971 ( .IN1(s14_msel_gnt_p0_2_), .IN2(n11262), .IN3(n2858), .IN4(
        n11263), .Q(n17341) );
  NAND4X0 U33972 ( .IN1(n11264), .IN2(n11265), .IN3(n11266), .IN4(n11267), 
        .QN(n11263) );
  NAND3X0 U33973 ( .IN1(n11280), .IN2(n3264), .IN3(n11281), .QN(n11264) );
  AO22X1 U33974 ( .IN1(s5_msel_gnt_p0[1]), .IN2(n13119), .IN3(n3002), .IN4(
        n13141), .Q(n17522) );
  NAND3X0 U33975 ( .IN1(n13142), .IN2(n13128), .IN3(n13143), .QN(n13141) );
  OA222X1 U33976 ( .IN1(n13125), .IN2(n3770), .IN3(n13144), .IN4(n3439), .IN5(
        n13145), .IN6(n3230), .Q(n13143) );
  OA21X1 U33977 ( .IN1(n13146), .IN2(n13147), .IN3(n13148), .Q(n13145) );
  AO22X1 U33978 ( .IN1(s5_msel_gnt_p0[2]), .IN2(n13119), .IN3(n3002), .IN4(
        n13120), .Q(n17521) );
  NAND4X0 U33979 ( .IN1(n13121), .IN2(n13122), .IN3(n13123), .IN4(n13124), 
        .QN(n13120) );
  NAND3X0 U33980 ( .IN1(n13137), .IN2(n3336), .IN3(n13138), .QN(n13121) );
  AO22X1 U33981 ( .IN1(s4_msel_gnt_p0[1]), .IN2(n12810), .IN3(n3018), .IN4(
        n12832), .Q(n17492) );
  NAND3X0 U33982 ( .IN1(n12833), .IN2(n12819), .IN3(n12834), .QN(n12832) );
  OA222X1 U33983 ( .IN1(n12816), .IN2(n3725), .IN3(n12835), .IN4(n3443), .IN5(
        n12836), .IN6(n3234), .Q(n12834) );
  OA21X1 U33984 ( .IN1(n12837), .IN2(n12838), .IN3(n12839), .Q(n12836) );
  AO22X1 U33985 ( .IN1(s4_msel_gnt_p0[2]), .IN2(n12810), .IN3(n3018), .IN4(
        n12811), .Q(n17491) );
  NAND4X0 U33986 ( .IN1(n12812), .IN2(n12813), .IN3(n12814), .IN4(n12815), 
        .QN(n12811) );
  NAND3X0 U33987 ( .IN1(n12828), .IN2(n3344), .IN3(n12829), .QN(n12812) );
  AO22X1 U33988 ( .IN1(s13_msel_gnt_p0_1_), .IN2(n10953), .IN3(n2874), .IN4(
        n10975), .Q(n17312) );
  NAND3X0 U33989 ( .IN1(n10976), .IN2(n10962), .IN3(n10977), .QN(n10975) );
  OA222X1 U33990 ( .IN1(n10959), .IN2(n4130), .IN3(n10978), .IN4(n3407), .IN5(
        n10979), .IN6(n3198), .Q(n10977) );
  OA21X1 U33991 ( .IN1(n10969), .IN2(n10983), .IN3(n10984), .Q(n10978) );
  AO22X1 U33992 ( .IN1(s13_msel_gnt_p0_2_), .IN2(n10953), .IN3(n2874), .IN4(
        n10954), .Q(n17311) );
  NAND4X0 U33993 ( .IN1(n10955), .IN2(n10956), .IN3(n10957), .IN4(n10958), 
        .QN(n10954) );
  NAND3X0 U33994 ( .IN1(n10971), .IN2(n3272), .IN3(n10972), .QN(n10955) );
  OA22X1 U33995 ( .IN1(n10964), .IN2(n10965), .IN3(n10966), .IN4(n3407), .Q(
        n10957) );
  AO22X1 U33996 ( .IN1(s12_msel_gnt_p0[1]), .IN2(n10643), .IN3(n2890), .IN4(
        n10665), .Q(n17282) );
  NAND3X0 U33997 ( .IN1(n10666), .IN2(n10652), .IN3(n10667), .QN(n10665) );
  OA222X1 U33998 ( .IN1(n10649), .IN2(n4085), .IN3(n10668), .IN4(n3411), .IN5(
        n10669), .IN6(n3202), .Q(n10667) );
  OA21X1 U33999 ( .IN1(n10670), .IN2(n10671), .IN3(n10672), .Q(n10669) );
  AO22X1 U34000 ( .IN1(s12_msel_gnt_p0[2]), .IN2(n10643), .IN3(n2890), .IN4(
        n10644), .Q(n17281) );
  NAND4X0 U34001 ( .IN1(n10645), .IN2(n10646), .IN3(n10647), .IN4(n10648), 
        .QN(n10644) );
  NAND3X0 U34002 ( .IN1(n10661), .IN2(n3280), .IN3(n10662), .QN(n10645) );
  AO22X1 U34003 ( .IN1(s3_msel_gnt_p0_1_), .IN2(n12501), .IN3(n3034), .IN4(
        n12523), .Q(n17462) );
  NAND3X0 U34004 ( .IN1(n12524), .IN2(n12510), .IN3(n12525), .QN(n12523) );
  OA222X1 U34005 ( .IN1(n12507), .IN2(n3680), .IN3(n12526), .IN4(n3447), .IN5(
        n12527), .IN6(n3238), .Q(n12525) );
  OA21X1 U34006 ( .IN1(n12528), .IN2(n12529), .IN3(n12530), .Q(n12527) );
  AO22X1 U34007 ( .IN1(test_so52), .IN2(n12501), .IN3(n3034), .IN4(n12502), 
        .Q(n17461) );
  NAND4X0 U34008 ( .IN1(n12503), .IN2(n12504), .IN3(n12505), .IN4(n12506), 
        .QN(n12502) );
  NAND3X0 U34009 ( .IN1(n12519), .IN2(n3352), .IN3(n12520), .QN(n12503) );
  AO22X1 U34010 ( .IN1(test_so48), .IN2(n12192), .IN3(n3050), .IN4(n12214), 
        .Q(n17432) );
  NAND3X0 U34011 ( .IN1(n12215), .IN2(n12201), .IN3(n12216), .QN(n12214) );
  OA222X1 U34012 ( .IN1(n12198), .IN2(n3635), .IN3(n12217), .IN4(n3451), .IN5(
        n12218), .IN6(n3242), .Q(n12216) );
  OA21X1 U34013 ( .IN1(n12219), .IN2(n12220), .IN3(n12221), .Q(n12218) );
  AO22X1 U34014 ( .IN1(s2_msel_gnt_p0_2_), .IN2(n12192), .IN3(n3050), .IN4(
        n12193), .Q(n17431) );
  NAND4X0 U34015 ( .IN1(n12194), .IN2(n12195), .IN3(n12196), .IN4(n12197), 
        .QN(n12193) );
  NAND3X0 U34016 ( .IN1(n12210), .IN2(n3360), .IN3(n12211), .QN(n12194) );
  AO22X1 U34017 ( .IN1(s11_msel_gnt_p0[1]), .IN2(n10334), .IN3(n2906), .IN4(
        n10356), .Q(n17252) );
  NAND3X0 U34018 ( .IN1(n10357), .IN2(n10343), .IN3(n10358), .QN(n10356) );
  OA222X1 U34019 ( .IN1(n10340), .IN2(n4040), .IN3(n10359), .IN4(n3415), .IN5(
        n10360), .IN6(n3206), .Q(n10358) );
  OA21X1 U34020 ( .IN1(n10350), .IN2(n10364), .IN3(n10365), .Q(n10359) );
  AO22X1 U34021 ( .IN1(s11_msel_gnt_p0[2]), .IN2(n10334), .IN3(n2906), .IN4(
        n10335), .Q(n17251) );
  NAND4X0 U34022 ( .IN1(n10336), .IN2(n10337), .IN3(n10338), .IN4(n10339), 
        .QN(n10335) );
  NAND3X0 U34023 ( .IN1(n10352), .IN2(n3288), .IN3(n10353), .QN(n10336) );
  OA22X1 U34024 ( .IN1(n10345), .IN2(n10346), .IN3(n10347), .IN4(n3415), .Q(
        n10338) );
  AO22X1 U34025 ( .IN1(s10_msel_gnt_p0[1]), .IN2(n10024), .IN3(n2922), .IN4(
        n10046), .Q(n17222) );
  NAND3X0 U34026 ( .IN1(n10047), .IN2(n10033), .IN3(n10048), .QN(n10046) );
  OA222X1 U34027 ( .IN1(n10030), .IN2(n3995), .IN3(n10049), .IN4(n3419), .IN5(
        n10050), .IN6(n3210), .Q(n10048) );
  OA21X1 U34028 ( .IN1(n10051), .IN2(n10052), .IN3(n10053), .Q(n10050) );
  AO22X1 U34029 ( .IN1(s10_msel_gnt_p0[2]), .IN2(n10024), .IN3(n2922), .IN4(
        n10025), .Q(n17221) );
  NAND4X0 U34030 ( .IN1(n10026), .IN2(n10027), .IN3(n10028), .IN4(n10029), 
        .QN(n10025) );
  NAND3X0 U34031 ( .IN1(n10042), .IN2(n3296), .IN3(n10043), .QN(n10026) );
  AO22X1 U34032 ( .IN1(s1_msel_gnt_p0_1_), .IN2(n11882), .IN3(n3066), .IN4(
        n11904), .Q(n17402) );
  NAND3X0 U34033 ( .IN1(n11905), .IN2(n11891), .IN3(n11906), .QN(n11904) );
  OA222X1 U34034 ( .IN1(n11888), .IN2(n3590), .IN3(n11907), .IN4(n3455), .IN5(
        n11908), .IN6(n3246), .Q(n11906) );
  OA21X1 U34035 ( .IN1(n11909), .IN2(n11910), .IN3(n11911), .Q(n11908) );
  AO22X1 U34036 ( .IN1(s1_msel_gnt_p0_2_), .IN2(n11882), .IN3(n3066), .IN4(
        n11883), .Q(n17401) );
  NAND4X0 U34037 ( .IN1(n11884), .IN2(n11885), .IN3(n11886), .IN4(n11887), 
        .QN(n11883) );
  NAND3X0 U34038 ( .IN1(n11900), .IN2(n3368), .IN3(n11901), .QN(n11884) );
  AO22X1 U34039 ( .IN1(s0_msel_gnt_p0[1]), .IN2(n11572), .IN3(n3082), .IN4(
        n11594), .Q(n17372) );
  NAND3X0 U34040 ( .IN1(n11595), .IN2(n11581), .IN3(n11596), .QN(n11594) );
  OA222X1 U34041 ( .IN1(n11578), .IN2(n3545), .IN3(n11597), .IN4(n3459), .IN5(
        n11598), .IN6(n3250), .Q(n11596) );
  OA21X1 U34042 ( .IN1(n11599), .IN2(n11600), .IN3(n11601), .Q(n11598) );
  AO22X1 U34043 ( .IN1(s0_msel_gnt_p0[2]), .IN2(n11572), .IN3(n3082), .IN4(
        n11573), .Q(n17371) );
  NAND4X0 U34044 ( .IN1(n11574), .IN2(n11575), .IN3(n11576), .IN4(n11577), 
        .QN(n11573) );
  NAND3X0 U34045 ( .IN1(n11590), .IN2(n3376), .IN3(n11591), .QN(n11574) );
  AO22X1 U34046 ( .IN1(s9_msel_gnt_p0_1_), .IN2(n9714), .IN3(n2938), .IN4(
        n9736), .Q(n17192) );
  NAND3X0 U34047 ( .IN1(n9737), .IN2(n9723), .IN3(n9738), .QN(n9736) );
  OA222X1 U34048 ( .IN1(n9720), .IN2(n3950), .IN3(n9739), .IN4(n3423), .IN5(
        n9740), .IN6(n3214), .Q(n9738) );
  OA21X1 U34049 ( .IN1(n9730), .IN2(n9744), .IN3(n9745), .Q(n9739) );
  AO22X1 U34050 ( .IN1(test_so75), .IN2(n9714), .IN3(n2938), .IN4(n9715), .Q(
        n17191) );
  NAND4X0 U34051 ( .IN1(n9716), .IN2(n9717), .IN3(n9718), .IN4(n9719), .QN(
        n9715) );
  NAND3X0 U34052 ( .IN1(n9732), .IN2(n3304), .IN3(n9733), .QN(n9716) );
  OA22X1 U34053 ( .IN1(n9725), .IN2(n9726), .IN3(n9727), .IN4(n3423), .Q(n9718) );
  AO22X1 U34054 ( .IN1(test_so71), .IN2(n9403), .IN3(n2954), .IN4(n9425), .Q(
        n17162) );
  NAND3X0 U34055 ( .IN1(n9426), .IN2(n9412), .IN3(n9427), .QN(n9425) );
  OA222X1 U34056 ( .IN1(n9409), .IN2(n3905), .IN3(n9428), .IN4(n3427), .IN5(
        n9429), .IN6(n3218), .Q(n9427) );
  OA21X1 U34057 ( .IN1(n9430), .IN2(n9431), .IN3(n9432), .Q(n9429) );
  AO22X1 U34058 ( .IN1(s8_msel_gnt_p0_2_), .IN2(n9403), .IN3(n2954), .IN4(
        n9404), .Q(n17161) );
  NAND4X0 U34059 ( .IN1(n9405), .IN2(n9406), .IN3(n9407), .IN4(n9408), .QN(
        n9404) );
  NAND3X0 U34060 ( .IN1(n9421), .IN2(n3312), .IN3(n9422), .QN(n9405) );
  AO22X1 U34061 ( .IN1(s7_msel_gnt_p1[1]), .IN2(n13804), .IN3(n2973), .IN4(
        n13822), .Q(n17585) );
  NAND3X0 U34062 ( .IN1(n13823), .IN2(n13806), .IN3(n13824), .QN(n13822) );
  OA222X1 U34063 ( .IN1(n13820), .IN2(n3868), .IN3(n13825), .IN4(n3432), .IN5(
        n13826), .IN6(n3223), .Q(n13824) );
  OA21X1 U34064 ( .IN1(n13817), .IN2(n13830), .IN3(n13831), .Q(n13825) );
  AO22X1 U34065 ( .IN1(s7_msel_gnt_p1[0]), .IN2(n13804), .IN3(n2973), .IN4(
        n13839), .Q(n17586) );
  NAND3X0 U34066 ( .IN1(n13823), .IN2(n13840), .IN3(n13841), .QN(n13839) );
  OR2X1 U34067 ( .IN1(n3867), .IN2(n13820), .Q(n13840) );
  OA221X1 U34068 ( .IN1(n3144), .IN2(n13842), .IN3(n18163), .IN4(n13843), 
        .IN5(n13813), .Q(n13841) );
  AO22X1 U34069 ( .IN1(s7_msel_gnt_p1[2]), .IN2(n13804), .IN3(n2973), .IN4(
        n13805), .Q(n17584) );
  NAND4X0 U34070 ( .IN1(n3145), .IN2(n13806), .IN3(n13807), .IN4(n13808), .QN(
        n13805) );
  OA22X1 U34071 ( .IN1(n13819), .IN2(n18163), .IN3(n13820), .IN4(n3869), .Q(
        n13807) );
  OA221X1 U34072 ( .IN1(n13809), .IN2(n3496), .IN3(n13810), .IN4(n3432), .IN5(
        n13811), .Q(n13808) );
  AO22X1 U34073 ( .IN1(s7_msel_gnt_p2_1_), .IN2(n13679), .IN3(n2965), .IN4(
        n13696), .Q(n17579) );
  NAND3X0 U34074 ( .IN1(n13697), .IN2(n13681), .IN3(n13698), .QN(n13696) );
  OA222X1 U34075 ( .IN1(n13694), .IN2(n3876), .IN3(n13699), .IN4(n3430), .IN5(
        n13700), .IN6(n3221), .Q(n13698) );
  OA21X1 U34076 ( .IN1(n13692), .IN2(n13704), .IN3(n13705), .Q(n13699) );
  AO22X1 U34077 ( .IN1(test_so68), .IN2(n13679), .IN3(n2965), .IN4(n13710), 
        .Q(n17580) );
  NAND3X0 U34078 ( .IN1(n13697), .IN2(n13711), .IN3(n13712), .QN(n13710) );
  OR2X1 U34079 ( .IN1(n3875), .IN2(n13694), .Q(n13711) );
  OA221X1 U34080 ( .IN1(n3141), .IN2(n13713), .IN3(n18164), .IN4(n13714), 
        .IN5(n13688), .Q(n13712) );
  AO22X1 U34081 ( .IN1(s7_msel_gnt_p2_2_), .IN2(n13679), .IN3(n2965), .IN4(
        n13680), .Q(n17578) );
  NAND4X0 U34082 ( .IN1(n3142), .IN2(n13681), .IN3(n13682), .IN4(n13683), .QN(
        n13680) );
  OA22X1 U34083 ( .IN1(n13693), .IN2(n18164), .IN3(n13694), .IN4(n3877), .Q(
        n13682) );
  OA221X1 U34084 ( .IN1(n13684), .IN2(n3494), .IN3(n13685), .IN4(n3430), .IN5(
        n13686), .Q(n13683) );
  AO22X1 U34085 ( .IN1(s6_msel_gnt_p1_1_), .IN2(n13495), .IN3(n2989), .IN4(
        n13513), .Q(n17555) );
  NAND3X0 U34086 ( .IN1(n13514), .IN2(n13497), .IN3(n13515), .QN(n13513) );
  OA222X1 U34087 ( .IN1(n13511), .IN2(n3823), .IN3(n13516), .IN4(n3436), .IN5(
        n13517), .IN6(n3227), .Q(n13515) );
  OA21X1 U34088 ( .IN1(n13508), .IN2(n13521), .IN3(n13522), .Q(n13516) );
  AO22X1 U34089 ( .IN1(s6_msel_gnt_p1_0_), .IN2(n13495), .IN3(n2989), .IN4(
        n13530), .Q(n17556) );
  NAND3X0 U34090 ( .IN1(n13514), .IN2(n13531), .IN3(n13532), .QN(n13530) );
  OR2X1 U34091 ( .IN1(n3822), .IN2(n13511), .Q(n13531) );
  OA221X1 U34092 ( .IN1(n3150), .IN2(n13533), .IN3(n18159), .IN4(n13534), 
        .IN5(n13504), .Q(n13532) );
  AO22X1 U34093 ( .IN1(test_so64), .IN2(n13495), .IN3(n2989), .IN4(n13496), 
        .Q(n17554) );
  NAND4X0 U34094 ( .IN1(n3151), .IN2(n13497), .IN3(n13498), .IN4(n13499), .QN(
        n13496) );
  OA22X1 U34095 ( .IN1(n13510), .IN2(n18159), .IN3(n13511), .IN4(n3824), .Q(
        n13498) );
  OA221X1 U34096 ( .IN1(n13500), .IN2(n3500), .IN3(n13501), .IN4(n3436), .IN5(
        n13502), .Q(n13499) );
  AO22X1 U34097 ( .IN1(s6_msel_gnt_p2[1]), .IN2(n13370), .IN3(n2981), .IN4(
        n13387), .Q(n17549) );
  NAND3X0 U34098 ( .IN1(n13388), .IN2(n13372), .IN3(n13389), .QN(n13387) );
  OA222X1 U34099 ( .IN1(n13385), .IN2(n3831), .IN3(n13390), .IN4(n3434), .IN5(
        n13391), .IN6(n3225), .Q(n13389) );
  OA21X1 U34100 ( .IN1(n13383), .IN2(n13395), .IN3(n13396), .Q(n13390) );
  AO22X1 U34101 ( .IN1(s6_msel_gnt_p2[0]), .IN2(n13370), .IN3(n2981), .IN4(
        n13401), .Q(n17550) );
  NAND3X0 U34102 ( .IN1(n13388), .IN2(n13402), .IN3(n13403), .QN(n13401) );
  OR2X1 U34103 ( .IN1(n3830), .IN2(n13385), .Q(n13402) );
  OA221X1 U34104 ( .IN1(n3147), .IN2(n13404), .IN3(n18165), .IN4(n13405), 
        .IN5(n13379), .Q(n13403) );
  AO22X1 U34105 ( .IN1(s6_msel_gnt_p2[2]), .IN2(n13370), .IN3(n2981), .IN4(
        n13371), .Q(n17548) );
  NAND4X0 U34106 ( .IN1(n3148), .IN2(n13372), .IN3(n13373), .IN4(n13374), .QN(
        n13371) );
  OA22X1 U34107 ( .IN1(n13384), .IN2(n18165), .IN3(n13385), .IN4(n3832), .Q(
        n13373) );
  OA221X1 U34108 ( .IN1(n13375), .IN2(n3498), .IN3(n13376), .IN4(n3434), .IN5(
        n13377), .Q(n13374) );
  AO22X1 U34109 ( .IN1(s14_msel_gnt_p1[1]), .IN2(n11329), .IN3(n2861), .IN4(
        n11347), .Q(n17345) );
  NAND3X0 U34110 ( .IN1(n11348), .IN2(n11331), .IN3(n11349), .QN(n11347) );
  OA222X1 U34111 ( .IN1(n11345), .IN2(n4183), .IN3(n11350), .IN4(n3404), .IN5(
        n11351), .IN6(n3195), .Q(n11349) );
  OA21X1 U34112 ( .IN1(n11342), .IN2(n11355), .IN3(n11356), .Q(n11350) );
  AO22X1 U34113 ( .IN1(s14_msel_gnt_p1[0]), .IN2(n11329), .IN3(n2861), .IN4(
        n11364), .Q(n17346) );
  NAND3X0 U34114 ( .IN1(n11348), .IN2(n11365), .IN3(n11366), .QN(n11364) );
  OR2X1 U34115 ( .IN1(n4182), .IN2(n11345), .Q(n11365) );
  OA221X1 U34116 ( .IN1(n3102), .IN2(n11367), .IN3(n18160), .IN4(n11368), 
        .IN5(n11338), .Q(n11366) );
  AO22X1 U34117 ( .IN1(s14_msel_gnt_p1[2]), .IN2(n11329), .IN3(n2861), .IN4(
        n11330), .Q(n17344) );
  NAND4X0 U34118 ( .IN1(n3103), .IN2(n11331), .IN3(n11332), .IN4(n11333), .QN(
        n11330) );
  OA22X1 U34119 ( .IN1(n11344), .IN2(n18160), .IN3(n11345), .IN4(n4184), .Q(
        n11332) );
  OA221X1 U34120 ( .IN1(n11334), .IN2(n3468), .IN3(n11335), .IN4(n3404), .IN5(
        n11336), .Q(n11333) );
  AO22X1 U34121 ( .IN1(test_so95), .IN2(n11204), .IN3(n2853), .IN4(n11221), 
        .Q(n17339) );
  NAND3X0 U34122 ( .IN1(n11222), .IN2(n11206), .IN3(n11223), .QN(n11221) );
  OA222X1 U34123 ( .IN1(n11219), .IN2(n4191), .IN3(n11224), .IN4(n3402), .IN5(
        n11225), .IN6(n3193), .Q(n11223) );
  OA21X1 U34124 ( .IN1(n11217), .IN2(n11229), .IN3(n11230), .Q(n11224) );
  AO22X1 U34125 ( .IN1(s14_msel_gnt_p2_0_), .IN2(n11204), .IN3(n2853), .IN4(
        n11235), .Q(n17340) );
  NAND3X0 U34126 ( .IN1(n11222), .IN2(n11236), .IN3(n11237), .QN(n11235) );
  OR2X1 U34127 ( .IN1(n4190), .IN2(n11219), .Q(n11236) );
  OA221X1 U34128 ( .IN1(n3099), .IN2(n11238), .IN3(n18166), .IN4(n11239), 
        .IN5(n11213), .Q(n11237) );
  AO22X1 U34129 ( .IN1(s14_msel_gnt_p2_2_), .IN2(n11204), .IN3(n2853), .IN4(
        n11205), .Q(n17338) );
  NAND4X0 U34130 ( .IN1(n3100), .IN2(n11206), .IN3(n11207), .IN4(n11208), .QN(
        n11205) );
  OA22X1 U34131 ( .IN1(n11218), .IN2(n18166), .IN3(n11219), .IN4(n4192), .Q(
        n11207) );
  OA221X1 U34132 ( .IN1(n11209), .IN2(n3466), .IN3(n11210), .IN4(n3402), .IN5(
        n11211), .Q(n11208) );
  AO22X1 U34133 ( .IN1(test_so60), .IN2(n13186), .IN3(n3005), .IN4(n13204), 
        .Q(n17525) );
  NAND3X0 U34134 ( .IN1(n13205), .IN2(n13188), .IN3(n13206), .QN(n13204) );
  OA222X1 U34135 ( .IN1(n13202), .IN2(n3778), .IN3(n13207), .IN4(n3440), .IN5(
        n13208), .IN6(n3231), .Q(n13206) );
  OA21X1 U34136 ( .IN1(n13199), .IN2(n13212), .IN3(n13213), .Q(n13207) );
  AO22X1 U34137 ( .IN1(s5_msel_gnt_p1_0_), .IN2(n13186), .IN3(n3005), .IN4(
        n13221), .Q(n17526) );
  NAND3X0 U34138 ( .IN1(n13205), .IN2(n13222), .IN3(n13223), .QN(n13221) );
  OR2X1 U34139 ( .IN1(n3777), .IN2(n13202), .Q(n13222) );
  OA221X1 U34140 ( .IN1(n3156), .IN2(n13224), .IN3(n18167), .IN4(n13225), 
        .IN5(n13195), .Q(n13223) );
  AO22X1 U34141 ( .IN1(s5_msel_gnt_p1_2_), .IN2(n13186), .IN3(n3005), .IN4(
        n13187), .Q(n17524) );
  NAND4X0 U34142 ( .IN1(n3157), .IN2(n13188), .IN3(n13189), .IN4(n13190), .QN(
        n13187) );
  OA22X1 U34143 ( .IN1(n13201), .IN2(n18167), .IN3(n13202), .IN4(n3779), .Q(
        n13189) );
  OA221X1 U34144 ( .IN1(n13191), .IN2(n3504), .IN3(n13192), .IN4(n3440), .IN5(
        n13193), .Q(n13190) );
  AO22X1 U34145 ( .IN1(s5_msel_gnt_p2[1]), .IN2(n13061), .IN3(n2997), .IN4(
        n13078), .Q(n17519) );
  NAND3X0 U34146 ( .IN1(n13079), .IN2(n13063), .IN3(n13080), .QN(n13078) );
  OA222X1 U34147 ( .IN1(n13076), .IN2(n3786), .IN3(n13081), .IN4(n3438), .IN5(
        n13082), .IN6(n3229), .Q(n13080) );
  OA21X1 U34148 ( .IN1(n13074), .IN2(n13086), .IN3(n13087), .Q(n13081) );
  AO22X1 U34149 ( .IN1(s5_msel_gnt_p2[0]), .IN2(n13061), .IN3(n2997), .IN4(
        n13092), .Q(n17520) );
  NAND3X0 U34150 ( .IN1(n13079), .IN2(n13093), .IN3(n13094), .QN(n13092) );
  OR2X1 U34151 ( .IN1(n3785), .IN2(n13076), .Q(n13093) );
  OA221X1 U34152 ( .IN1(n3153), .IN2(n13095), .IN3(n18168), .IN4(n13096), 
        .IN5(n13070), .Q(n13094) );
  AO22X1 U34153 ( .IN1(s5_msel_gnt_p2[2]), .IN2(n13061), .IN3(n2997), .IN4(
        n13062), .Q(n17518) );
  NAND4X0 U34154 ( .IN1(n3154), .IN2(n13063), .IN3(n13064), .IN4(n13065), .QN(
        n13062) );
  OA22X1 U34155 ( .IN1(n13075), .IN2(n18168), .IN3(n13076), .IN4(n3787), .Q(
        n13064) );
  OA221X1 U34156 ( .IN1(n13066), .IN2(n3502), .IN3(n13067), .IN4(n3438), .IN5(
        n13068), .Q(n13065) );
  AO22X1 U34157 ( .IN1(s4_msel_gnt_p1_1_), .IN2(n12877), .IN3(n3021), .IN4(
        n12895), .Q(n17495) );
  NAND3X0 U34158 ( .IN1(n12896), .IN2(n12879), .IN3(n12897), .QN(n12895) );
  OA222X1 U34159 ( .IN1(n12893), .IN2(n3733), .IN3(n12898), .IN4(n3444), .IN5(
        n12899), .IN6(n3235), .Q(n12897) );
  OA21X1 U34160 ( .IN1(n12890), .IN2(n12903), .IN3(n12904), .Q(n12898) );
  AO22X1 U34161 ( .IN1(test_so56), .IN2(n12877), .IN3(n3021), .IN4(n12912), 
        .Q(n17496) );
  NAND3X0 U34162 ( .IN1(n12896), .IN2(n12913), .IN3(n12914), .QN(n12912) );
  OR2X1 U34163 ( .IN1(n3732), .IN2(n12893), .Q(n12913) );
  OA221X1 U34164 ( .IN1(n3162), .IN2(n12915), .IN3(n18169), .IN4(n12916), 
        .IN5(n12886), .Q(n12914) );
  AO22X1 U34165 ( .IN1(s4_msel_gnt_p1_2_), .IN2(n12877), .IN3(n3021), .IN4(
        n12878), .Q(n17494) );
  NAND4X0 U34166 ( .IN1(n3163), .IN2(n12879), .IN3(n12880), .IN4(n12881), .QN(
        n12878) );
  OA22X1 U34167 ( .IN1(n12892), .IN2(n18169), .IN3(n12893), .IN4(n3734), .Q(
        n12880) );
  OA221X1 U34168 ( .IN1(n12882), .IN2(n3508), .IN3(n12883), .IN4(n3444), .IN5(
        n12884), .Q(n12881) );
  AO22X1 U34169 ( .IN1(s4_msel_gnt_p2[1]), .IN2(n12752), .IN3(n3013), .IN4(
        n12769), .Q(n17489) );
  NAND3X0 U34170 ( .IN1(n12770), .IN2(n12754), .IN3(n12771), .QN(n12769) );
  OA222X1 U34171 ( .IN1(n12767), .IN2(n3741), .IN3(n12772), .IN4(n3442), .IN5(
        n12773), .IN6(n3233), .Q(n12771) );
  OA21X1 U34172 ( .IN1(n12765), .IN2(n12777), .IN3(n12778), .Q(n12772) );
  AO22X1 U34173 ( .IN1(s4_msel_gnt_p2[0]), .IN2(n12752), .IN3(n3013), .IN4(
        n12783), .Q(n17490) );
  NAND3X0 U34174 ( .IN1(n12770), .IN2(n12784), .IN3(n12785), .QN(n12783) );
  OR2X1 U34175 ( .IN1(n3740), .IN2(n12767), .Q(n12784) );
  OA221X1 U34176 ( .IN1(n3159), .IN2(n12786), .IN3(n18170), .IN4(n12787), 
        .IN5(n12761), .Q(n12785) );
  AO22X1 U34177 ( .IN1(s4_msel_gnt_p2[2]), .IN2(n12752), .IN3(n3013), .IN4(
        n12753), .Q(n17488) );
  NAND4X0 U34178 ( .IN1(n3160), .IN2(n12754), .IN3(n12755), .IN4(n12756), .QN(
        n12753) );
  OA22X1 U34179 ( .IN1(n12766), .IN2(n18170), .IN3(n12767), .IN4(n3742), .Q(
        n12755) );
  OA221X1 U34180 ( .IN1(n12757), .IN2(n3506), .IN3(n12758), .IN4(n3442), .IN5(
        n12759), .Q(n12756) );
  AO22X1 U34181 ( .IN1(s13_msel_gnt_p1[1]), .IN2(n11020), .IN3(n2877), .IN4(
        n11038), .Q(n17315) );
  NAND3X0 U34182 ( .IN1(n11039), .IN2(n11022), .IN3(n11040), .QN(n11038) );
  OA222X1 U34183 ( .IN1(n11036), .IN2(n4138), .IN3(n11041), .IN4(n3408), .IN5(
        n11042), .IN6(n3199), .Q(n11040) );
  OA21X1 U34184 ( .IN1(n11033), .IN2(n11046), .IN3(n11047), .Q(n11041) );
  AO22X1 U34185 ( .IN1(s13_msel_gnt_p1[0]), .IN2(n11020), .IN3(n2877), .IN4(
        n11055), .Q(n17316) );
  NAND3X0 U34186 ( .IN1(n11039), .IN2(n11056), .IN3(n11057), .QN(n11055) );
  OR2X1 U34187 ( .IN1(n4137), .IN2(n11036), .Q(n11056) );
  OA221X1 U34188 ( .IN1(n3108), .IN2(n11058), .IN3(n18171), .IN4(n11059), 
        .IN5(n11029), .Q(n11057) );
  AO22X1 U34189 ( .IN1(s13_msel_gnt_p1[2]), .IN2(n11020), .IN3(n2877), .IN4(
        n11021), .Q(n17314) );
  NAND4X0 U34190 ( .IN1(n3109), .IN2(n11022), .IN3(n11023), .IN4(n11024), .QN(
        n11021) );
  OA22X1 U34191 ( .IN1(n11035), .IN2(n18171), .IN3(n11036), .IN4(n4139), .Q(
        n11023) );
  OA221X1 U34192 ( .IN1(n11025), .IN2(n3472), .IN3(n11026), .IN4(n3408), .IN5(
        n11027), .Q(n11024) );
  AO22X1 U34193 ( .IN1(s13_msel_gnt_p2_1_), .IN2(n10895), .IN3(n2869), .IN4(
        n10912), .Q(n17309) );
  NAND3X0 U34194 ( .IN1(n10913), .IN2(n10897), .IN3(n10914), .QN(n10912) );
  OA222X1 U34195 ( .IN1(n10910), .IN2(n4146), .IN3(n10915), .IN4(n3406), .IN5(
        n10916), .IN6(n3197), .Q(n10914) );
  OA21X1 U34196 ( .IN1(n10908), .IN2(n10920), .IN3(n10921), .Q(n10915) );
  AO22X1 U34197 ( .IN1(test_so91), .IN2(n10895), .IN3(n2869), .IN4(n10926), 
        .Q(n17310) );
  NAND3X0 U34198 ( .IN1(n10913), .IN2(n10927), .IN3(n10928), .QN(n10926) );
  OR2X1 U34199 ( .IN1(n4145), .IN2(n10910), .Q(n10927) );
  OA221X1 U34200 ( .IN1(n3105), .IN2(n10929), .IN3(n18172), .IN4(n10930), 
        .IN5(n10904), .Q(n10928) );
  AO22X1 U34201 ( .IN1(s13_msel_gnt_p2_2_), .IN2(n10895), .IN3(n2869), .IN4(
        n10896), .Q(n17308) );
  NAND4X0 U34202 ( .IN1(n3106), .IN2(n10897), .IN3(n10898), .IN4(n10899), .QN(
        n10896) );
  OA22X1 U34203 ( .IN1(n10909), .IN2(n18172), .IN3(n10910), .IN4(n4147), .Q(
        n10898) );
  OA221X1 U34204 ( .IN1(n10900), .IN2(n3470), .IN3(n10901), .IN4(n3406), .IN5(
        n10902), .Q(n10899) );
  AO22X1 U34205 ( .IN1(s12_msel_gnt_p1_1_), .IN2(n10710), .IN3(n2893), .IN4(
        n10728), .Q(n17285) );
  NAND3X0 U34206 ( .IN1(n10729), .IN2(n10712), .IN3(n10730), .QN(n10728) );
  OA222X1 U34207 ( .IN1(n10726), .IN2(n4093), .IN3(n10731), .IN4(n3412), .IN5(
        n10732), .IN6(n3203), .Q(n10730) );
  OA21X1 U34208 ( .IN1(n10723), .IN2(n10736), .IN3(n10737), .Q(n10731) );
  AO22X1 U34209 ( .IN1(s12_msel_gnt_p1_0_), .IN2(n10710), .IN3(n2893), .IN4(
        n10745), .Q(n17286) );
  NAND3X0 U34210 ( .IN1(n10729), .IN2(n10746), .IN3(n10747), .QN(n10745) );
  OR2X1 U34211 ( .IN1(n4092), .IN2(n10726), .Q(n10746) );
  OA221X1 U34212 ( .IN1(n3114), .IN2(n10748), .IN3(n18173), .IN4(n10749), 
        .IN5(n10719), .Q(n10747) );
  AO22X1 U34213 ( .IN1(test_so87), .IN2(n10710), .IN3(n2893), .IN4(n10711), 
        .Q(n17284) );
  NAND4X0 U34214 ( .IN1(n3115), .IN2(n10712), .IN3(n10713), .IN4(n10714), .QN(
        n10711) );
  OA22X1 U34215 ( .IN1(n10725), .IN2(n18173), .IN3(n10726), .IN4(n4094), .Q(
        n10713) );
  OA221X1 U34216 ( .IN1(n10715), .IN2(n3476), .IN3(n10716), .IN4(n3412), .IN5(
        n10717), .Q(n10714) );
  AO22X1 U34217 ( .IN1(s12_msel_gnt_p2[1]), .IN2(n10585), .IN3(n2885), .IN4(
        n10602), .Q(n17279) );
  NAND3X0 U34218 ( .IN1(n10603), .IN2(n10587), .IN3(n10604), .QN(n10602) );
  OA222X1 U34219 ( .IN1(n10600), .IN2(n4101), .IN3(n10605), .IN4(n3410), .IN5(
        n10606), .IN6(n3201), .Q(n10604) );
  OA21X1 U34220 ( .IN1(n10598), .IN2(n10610), .IN3(n10611), .Q(n10605) );
  AO22X1 U34221 ( .IN1(s12_msel_gnt_p2[0]), .IN2(n10585), .IN3(n2885), .IN4(
        n10616), .Q(n17280) );
  NAND3X0 U34222 ( .IN1(n10603), .IN2(n10617), .IN3(n10618), .QN(n10616) );
  OR2X1 U34223 ( .IN1(n4100), .IN2(n10600), .Q(n10617) );
  OA221X1 U34224 ( .IN1(n3111), .IN2(n10619), .IN3(n18174), .IN4(n10620), 
        .IN5(n10594), .Q(n10618) );
  AO22X1 U34225 ( .IN1(s12_msel_gnt_p2[2]), .IN2(n10585), .IN3(n2885), .IN4(
        n10586), .Q(n17278) );
  NAND4X0 U34226 ( .IN1(n3112), .IN2(n10587), .IN3(n10588), .IN4(n10589), .QN(
        n10586) );
  OA22X1 U34227 ( .IN1(n10599), .IN2(n18174), .IN3(n10600), .IN4(n4102), .Q(
        n10588) );
  OA221X1 U34228 ( .IN1(n10590), .IN2(n3474), .IN3(n10591), .IN4(n3410), .IN5(
        n10592), .Q(n10589) );
  AO22X1 U34229 ( .IN1(s3_msel_gnt_p1[1]), .IN2(n12568), .IN3(n3037), .IN4(
        n12586), .Q(n17465) );
  NAND3X0 U34230 ( .IN1(n12587), .IN2(n12570), .IN3(n12588), .QN(n12586) );
  OA222X1 U34231 ( .IN1(n12584), .IN2(n3688), .IN3(n12589), .IN4(n3448), .IN5(
        n12590), .IN6(n3239), .Q(n12588) );
  OA21X1 U34232 ( .IN1(n12581), .IN2(n12594), .IN3(n12595), .Q(n12589) );
  AO22X1 U34233 ( .IN1(s3_msel_gnt_p1[0]), .IN2(n12568), .IN3(n3037), .IN4(
        n12603), .Q(n17466) );
  NAND3X0 U34234 ( .IN1(n12587), .IN2(n12604), .IN3(n12605), .QN(n12603) );
  OR2X1 U34235 ( .IN1(n3687), .IN2(n12584), .Q(n12604) );
  OA221X1 U34236 ( .IN1(n3168), .IN2(n12606), .IN3(n18175), .IN4(n12607), 
        .IN5(n12577), .Q(n12605) );
  AO22X1 U34237 ( .IN1(s3_msel_gnt_p1[2]), .IN2(n12568), .IN3(n3037), .IN4(
        n12569), .Q(n17464) );
  NAND4X0 U34238 ( .IN1(n3169), .IN2(n12570), .IN3(n12571), .IN4(n12572), .QN(
        n12569) );
  OA22X1 U34239 ( .IN1(n12583), .IN2(n18175), .IN3(n12584), .IN4(n3689), .Q(
        n12571) );
  OA221X1 U34240 ( .IN1(n12573), .IN2(n3512), .IN3(n12574), .IN4(n3448), .IN5(
        n12575), .Q(n12572) );
  AO22X1 U34241 ( .IN1(s3_msel_gnt_p2_1_), .IN2(n12443), .IN3(n3029), .IN4(
        n12460), .Q(n17459) );
  NAND3X0 U34242 ( .IN1(n12461), .IN2(n12445), .IN3(n12462), .QN(n12460) );
  OA222X1 U34243 ( .IN1(n12458), .IN2(n3696), .IN3(n12463), .IN4(n3446), .IN5(
        n12464), .IN6(n3237), .Q(n12462) );
  OA21X1 U34244 ( .IN1(n12456), .IN2(n12468), .IN3(n12469), .Q(n12463) );
  AO22X1 U34245 ( .IN1(s3_msel_gnt_p2_0_), .IN2(n12443), .IN3(n3029), .IN4(
        n12474), .Q(n17460) );
  NAND3X0 U34246 ( .IN1(n12461), .IN2(n12475), .IN3(n12476), .QN(n12474) );
  OR2X1 U34247 ( .IN1(n3695), .IN2(n12458), .Q(n12475) );
  OA221X1 U34248 ( .IN1(n3165), .IN2(n12477), .IN3(n18176), .IN4(n12478), 
        .IN5(n12452), .Q(n12476) );
  AO22X1 U34249 ( .IN1(test_so53), .IN2(n12443), .IN3(n3029), .IN4(n12444), 
        .Q(n17458) );
  NAND4X0 U34250 ( .IN1(n3166), .IN2(n12445), .IN3(n12446), .IN4(n12447), .QN(
        n12444) );
  OA22X1 U34251 ( .IN1(n12457), .IN2(n18176), .IN3(n12458), .IN4(n3697), .Q(
        n12446) );
  OA221X1 U34252 ( .IN1(n12448), .IN2(n3510), .IN3(n12449), .IN4(n3446), .IN5(
        n12450), .Q(n12447) );
  AO22X1 U34253 ( .IN1(s2_msel_gnt_p1[1]), .IN2(n12259), .IN3(n3053), .IN4(
        n12277), .Q(n17435) );
  NAND3X0 U34254 ( .IN1(n12278), .IN2(n12261), .IN3(n12279), .QN(n12277) );
  OA222X1 U34255 ( .IN1(n12275), .IN2(n3643), .IN3(n12280), .IN4(n3452), .IN5(
        n12281), .IN6(n3243), .Q(n12279) );
  OA21X1 U34256 ( .IN1(n12272), .IN2(n12285), .IN3(n12286), .Q(n12280) );
  AO22X1 U34257 ( .IN1(s2_msel_gnt_p1[0]), .IN2(n12259), .IN3(n3053), .IN4(
        n12294), .Q(n17436) );
  NAND3X0 U34258 ( .IN1(n12278), .IN2(n12295), .IN3(n12296), .QN(n12294) );
  OR2X1 U34259 ( .IN1(n3642), .IN2(n12275), .Q(n12295) );
  OA221X1 U34260 ( .IN1(n3174), .IN2(n12297), .IN3(n18161), .IN4(n12298), 
        .IN5(n12268), .Q(n12296) );
  AO22X1 U34261 ( .IN1(s2_msel_gnt_p1[2]), .IN2(n12259), .IN3(n3053), .IN4(
        n12260), .Q(n17434) );
  NAND4X0 U34262 ( .IN1(n3175), .IN2(n12261), .IN3(n12262), .IN4(n12263), .QN(
        n12260) );
  OA22X1 U34263 ( .IN1(n12274), .IN2(n18161), .IN3(n12275), .IN4(n3644), .Q(
        n12262) );
  OA221X1 U34264 ( .IN1(n12264), .IN2(n3516), .IN3(n12265), .IN4(n3452), .IN5(
        n12266), .Q(n12263) );
  AO22X1 U34265 ( .IN1(test_so49), .IN2(n12134), .IN3(n3045), .IN4(n12151), 
        .Q(n17429) );
  NAND3X0 U34266 ( .IN1(n12152), .IN2(n12136), .IN3(n12153), .QN(n12151) );
  OA222X1 U34267 ( .IN1(n12149), .IN2(n3651), .IN3(n12154), .IN4(n3450), .IN5(
        n12155), .IN6(n3241), .Q(n12153) );
  OA21X1 U34268 ( .IN1(n12147), .IN2(n12159), .IN3(n12160), .Q(n12154) );
  AO22X1 U34269 ( .IN1(s2_msel_gnt_p2_0_), .IN2(n12134), .IN3(n3045), .IN4(
        n12165), .Q(n17430) );
  NAND3X0 U34270 ( .IN1(n12152), .IN2(n12166), .IN3(n12167), .QN(n12165) );
  OR2X1 U34271 ( .IN1(n3650), .IN2(n12149), .Q(n12166) );
  OA221X1 U34272 ( .IN1(n3171), .IN2(n12168), .IN3(n18177), .IN4(n12169), 
        .IN5(n12143), .Q(n12167) );
  AO22X1 U34273 ( .IN1(s2_msel_gnt_p2_2_), .IN2(n12134), .IN3(n3045), .IN4(
        n12135), .Q(n17428) );
  NAND4X0 U34274 ( .IN1(n3172), .IN2(n12136), .IN3(n12137), .IN4(n12138), .QN(
        n12135) );
  OA22X1 U34275 ( .IN1(n12148), .IN2(n18177), .IN3(n12149), .IN4(n3652), .Q(
        n12137) );
  OA221X1 U34276 ( .IN1(n12139), .IN2(n3514), .IN3(n12140), .IN4(n3450), .IN5(
        n12141), .Q(n12138) );
  AO22X1 U34277 ( .IN1(test_so83), .IN2(n10401), .IN3(n2909), .IN4(n10419), 
        .Q(n17255) );
  NAND3X0 U34278 ( .IN1(n10420), .IN2(n10403), .IN3(n10421), .QN(n10419) );
  OA222X1 U34279 ( .IN1(n10417), .IN2(n4048), .IN3(n10422), .IN4(n3416), .IN5(
        n10423), .IN6(n3207), .Q(n10421) );
  OA21X1 U34280 ( .IN1(n10414), .IN2(n10427), .IN3(n10428), .Q(n10422) );
  AO22X1 U34281 ( .IN1(s11_msel_gnt_p1_0_), .IN2(n10401), .IN3(n2909), .IN4(
        n10436), .Q(n17256) );
  NAND3X0 U34282 ( .IN1(n10420), .IN2(n10437), .IN3(n10438), .QN(n10436) );
  OR2X1 U34283 ( .IN1(n4047), .IN2(n10417), .Q(n10437) );
  OA221X1 U34284 ( .IN1(n3120), .IN2(n10439), .IN3(n18178), .IN4(n10440), 
        .IN5(n10410), .Q(n10438) );
  AO22X1 U34285 ( .IN1(s11_msel_gnt_p1_2_), .IN2(n10401), .IN3(n2909), .IN4(
        n10402), .Q(n17254) );
  NAND4X0 U34286 ( .IN1(n3121), .IN2(n10403), .IN3(n10404), .IN4(n10405), .QN(
        n10402) );
  OA22X1 U34287 ( .IN1(n10416), .IN2(n18178), .IN3(n10417), .IN4(n4049), .Q(
        n10404) );
  OA221X1 U34288 ( .IN1(n10406), .IN2(n3480), .IN3(n10407), .IN4(n3416), .IN5(
        n10408), .Q(n10405) );
  AO22X1 U34289 ( .IN1(s11_msel_gnt_p2[1]), .IN2(n10276), .IN3(n2901), .IN4(
        n10293), .Q(n17249) );
  NAND3X0 U34290 ( .IN1(n10294), .IN2(n10278), .IN3(n10295), .QN(n10293) );
  OA222X1 U34291 ( .IN1(n10291), .IN2(n4056), .IN3(n10296), .IN4(n3414), .IN5(
        n10297), .IN6(n3205), .Q(n10295) );
  OA21X1 U34292 ( .IN1(n10289), .IN2(n10301), .IN3(n10302), .Q(n10296) );
  AO22X1 U34293 ( .IN1(s11_msel_gnt_p2[0]), .IN2(n10276), .IN3(n2901), .IN4(
        n10307), .Q(n17250) );
  NAND3X0 U34294 ( .IN1(n10294), .IN2(n10308), .IN3(n10309), .QN(n10307) );
  OR2X1 U34295 ( .IN1(n4055), .IN2(n10291), .Q(n10308) );
  OA221X1 U34296 ( .IN1(n3117), .IN2(n10310), .IN3(n18179), .IN4(n10311), 
        .IN5(n10285), .Q(n10309) );
  AO22X1 U34297 ( .IN1(s11_msel_gnt_p2[2]), .IN2(n10276), .IN3(n2901), .IN4(
        n10277), .Q(n17248) );
  NAND4X0 U34298 ( .IN1(n3118), .IN2(n10278), .IN3(n10279), .IN4(n10280), .QN(
        n10277) );
  OA22X1 U34299 ( .IN1(n10290), .IN2(n18179), .IN3(n10291), .IN4(n4057), .Q(
        n10279) );
  OA221X1 U34300 ( .IN1(n10281), .IN2(n3478), .IN3(n10282), .IN4(n3414), .IN5(
        n10283), .Q(n10280) );
  AO22X1 U34301 ( .IN1(s10_msel_gnt_p1_1_), .IN2(n10091), .IN3(n2925), .IN4(
        n10109), .Q(n17225) );
  NAND3X0 U34302 ( .IN1(n10110), .IN2(n10093), .IN3(n10111), .QN(n10109) );
  OA222X1 U34303 ( .IN1(n10107), .IN2(n4003), .IN3(n10112), .IN4(n3420), .IN5(
        n10113), .IN6(n3211), .Q(n10111) );
  OA21X1 U34304 ( .IN1(n10104), .IN2(n10117), .IN3(n10118), .Q(n10112) );
  AO22X1 U34305 ( .IN1(test_so79), .IN2(n10091), .IN3(n2925), .IN4(n10126), 
        .Q(n17226) );
  NAND3X0 U34306 ( .IN1(n10110), .IN2(n10127), .IN3(n10128), .QN(n10126) );
  OR2X1 U34307 ( .IN1(n4002), .IN2(n10107), .Q(n10127) );
  OA221X1 U34308 ( .IN1(n3126), .IN2(n10129), .IN3(n18180), .IN4(n10130), 
        .IN5(n10100), .Q(n10128) );
  AO22X1 U34309 ( .IN1(s10_msel_gnt_p1_2_), .IN2(n10091), .IN3(n2925), .IN4(
        n10092), .Q(n17224) );
  NAND4X0 U34310 ( .IN1(n3127), .IN2(n10093), .IN3(n10094), .IN4(n10095), .QN(
        n10092) );
  OA22X1 U34311 ( .IN1(n10106), .IN2(n18180), .IN3(n10107), .IN4(n4004), .Q(
        n10094) );
  OA221X1 U34312 ( .IN1(n10096), .IN2(n3484), .IN3(n10097), .IN4(n3420), .IN5(
        n10098), .Q(n10095) );
  AO22X1 U34313 ( .IN1(s10_msel_gnt_p2[1]), .IN2(n9966), .IN3(n2917), .IN4(
        n9983), .Q(n17219) );
  NAND3X0 U34314 ( .IN1(n9984), .IN2(n9968), .IN3(n9985), .QN(n9983) );
  OA222X1 U34315 ( .IN1(n9981), .IN2(n4011), .IN3(n9986), .IN4(n3418), .IN5(
        n9987), .IN6(n3209), .Q(n9985) );
  OA21X1 U34316 ( .IN1(n9979), .IN2(n9991), .IN3(n9992), .Q(n9986) );
  AO22X1 U34317 ( .IN1(s10_msel_gnt_p2[0]), .IN2(n9966), .IN3(n2917), .IN4(
        n9997), .Q(n17220) );
  NAND3X0 U34318 ( .IN1(n9984), .IN2(n9998), .IN3(n9999), .QN(n9997) );
  OR2X1 U34319 ( .IN1(n4010), .IN2(n9981), .Q(n9998) );
  OA221X1 U34320 ( .IN1(n3123), .IN2(n10000), .IN3(n18181), .IN4(n10001), 
        .IN5(n9975), .Q(n9999) );
  AO22X1 U34321 ( .IN1(s10_msel_gnt_p2[2]), .IN2(n9966), .IN3(n2917), .IN4(
        n9967), .Q(n17218) );
  NAND4X0 U34322 ( .IN1(n3124), .IN2(n9968), .IN3(n9969), .IN4(n9970), .QN(
        n9967) );
  OA22X1 U34323 ( .IN1(n9980), .IN2(n18181), .IN3(n9981), .IN4(n4012), .Q(
        n9969) );
  OA221X1 U34324 ( .IN1(n9971), .IN2(n3482), .IN3(n9972), .IN4(n3418), .IN5(
        n9973), .Q(n9970) );
  AO22X1 U34325 ( .IN1(s1_msel_gnt_p1[1]), .IN2(n11949), .IN3(n3069), .IN4(
        n11967), .Q(n17405) );
  NAND3X0 U34326 ( .IN1(n11968), .IN2(n11951), .IN3(n11969), .QN(n11967) );
  OA222X1 U34327 ( .IN1(n11965), .IN2(n3598), .IN3(n11970), .IN4(n3456), .IN5(
        n11971), .IN6(n3247), .Q(n11969) );
  OA21X1 U34328 ( .IN1(n11962), .IN2(n11975), .IN3(n11976), .Q(n11970) );
  AO22X1 U34329 ( .IN1(s1_msel_gnt_p1[0]), .IN2(n11949), .IN3(n3069), .IN4(
        n11984), .Q(n17406) );
  NAND3X0 U34330 ( .IN1(n11968), .IN2(n11985), .IN3(n11986), .QN(n11984) );
  OR2X1 U34331 ( .IN1(n3597), .IN2(n11965), .Q(n11985) );
  OA221X1 U34332 ( .IN1(n3180), .IN2(n11987), .IN3(n18182), .IN4(n11988), 
        .IN5(n11958), .Q(n11986) );
  AO22X1 U34333 ( .IN1(s1_msel_gnt_p1[2]), .IN2(n11949), .IN3(n3069), .IN4(
        n11950), .Q(n17404) );
  NAND4X0 U34334 ( .IN1(n3181), .IN2(n11951), .IN3(n11952), .IN4(n11953), .QN(
        n11950) );
  OA22X1 U34335 ( .IN1(n11964), .IN2(n18182), .IN3(n11965), .IN4(n3599), .Q(
        n11952) );
  OA221X1 U34336 ( .IN1(n11954), .IN2(n3520), .IN3(n11955), .IN4(n3456), .IN5(
        n11956), .Q(n11953) );
  AO22X1 U34337 ( .IN1(s1_msel_gnt_p2_1_), .IN2(n11824), .IN3(n3061), .IN4(
        n11841), .Q(n17399) );
  NAND3X0 U34338 ( .IN1(n11842), .IN2(n11826), .IN3(n11843), .QN(n11841) );
  OA222X1 U34339 ( .IN1(n11839), .IN2(n3606), .IN3(n11844), .IN4(n3454), .IN5(
        n11845), .IN6(n3245), .Q(n11843) );
  OA21X1 U34340 ( .IN1(n11837), .IN2(n11849), .IN3(n11850), .Q(n11844) );
  AO22X1 U34341 ( .IN1(test_so45), .IN2(n11824), .IN3(n3061), .IN4(n11855), 
        .Q(n17400) );
  NAND3X0 U34342 ( .IN1(n11842), .IN2(n11856), .IN3(n11857), .QN(n11855) );
  OR2X1 U34343 ( .IN1(n3605), .IN2(n11839), .Q(n11856) );
  OA221X1 U34344 ( .IN1(n3177), .IN2(n11858), .IN3(n18183), .IN4(n11859), 
        .IN5(n11833), .Q(n11857) );
  AO22X1 U34345 ( .IN1(s1_msel_gnt_p2_2_), .IN2(n11824), .IN3(n3061), .IN4(
        n11825), .Q(n17398) );
  NAND4X0 U34346 ( .IN1(n3178), .IN2(n11826), .IN3(n11827), .IN4(n11828), .QN(
        n11825) );
  OA22X1 U34347 ( .IN1(n11838), .IN2(n18183), .IN3(n11839), .IN4(n3607), .Q(
        n11827) );
  OA221X1 U34348 ( .IN1(n11829), .IN2(n3518), .IN3(n11830), .IN4(n3454), .IN5(
        n11831), .Q(n11828) );
  AO22X1 U34349 ( .IN1(s0_msel_gnt_p1_1_), .IN2(n11639), .IN3(n3085), .IN4(
        n11657), .Q(n17375) );
  NAND3X0 U34350 ( .IN1(n11658), .IN2(n11641), .IN3(n11659), .QN(n11657) );
  OA222X1 U34351 ( .IN1(n11655), .IN2(n3553), .IN3(n11660), .IN4(n3460), .IN5(
        n11661), .IN6(n3251), .Q(n11659) );
  OA21X1 U34352 ( .IN1(n11652), .IN2(n11665), .IN3(n11666), .Q(n11660) );
  AO22X1 U34353 ( .IN1(s0_msel_gnt_p1_0_), .IN2(n11639), .IN3(n3085), .IN4(
        n11674), .Q(n17376) );
  NAND3X0 U34354 ( .IN1(n11658), .IN2(n11675), .IN3(n11676), .QN(n11674) );
  OR2X1 U34355 ( .IN1(n3552), .IN2(n11655), .Q(n11675) );
  OA221X1 U34356 ( .IN1(n3186), .IN2(n11677), .IN3(n18184), .IN4(n11678), 
        .IN5(n11648), .Q(n11676) );
  AO22X1 U34357 ( .IN1(test_so41), .IN2(n11639), .IN3(n3085), .IN4(n11640), 
        .Q(n17374) );
  NAND4X0 U34358 ( .IN1(n3187), .IN2(n11641), .IN3(n11642), .IN4(n11643), .QN(
        n11640) );
  OA22X1 U34359 ( .IN1(n11654), .IN2(n18184), .IN3(n11655), .IN4(n3554), .Q(
        n11642) );
  OA221X1 U34360 ( .IN1(n11644), .IN2(n3524), .IN3(n11645), .IN4(n3460), .IN5(
        n11646), .Q(n11643) );
  AO22X1 U34361 ( .IN1(s0_msel_gnt_p2[1]), .IN2(n11514), .IN3(n3077), .IN4(
        n11531), .Q(n17369) );
  NAND3X0 U34362 ( .IN1(n11532), .IN2(n11516), .IN3(n11533), .QN(n11531) );
  OA222X1 U34363 ( .IN1(n11529), .IN2(n3561), .IN3(n11534), .IN4(n3458), .IN5(
        n11535), .IN6(n3249), .Q(n11533) );
  OA21X1 U34364 ( .IN1(n11527), .IN2(n11539), .IN3(n11540), .Q(n11534) );
  AO22X1 U34365 ( .IN1(s0_msel_gnt_p2[0]), .IN2(n11514), .IN3(n3077), .IN4(
        n11545), .Q(n17370) );
  NAND3X0 U34366 ( .IN1(n11532), .IN2(n11546), .IN3(n11547), .QN(n11545) );
  OR2X1 U34367 ( .IN1(n3560), .IN2(n11529), .Q(n11546) );
  OA221X1 U34368 ( .IN1(n3183), .IN2(n11548), .IN3(n18185), .IN4(n11549), 
        .IN5(n11523), .Q(n11547) );
  AO22X1 U34369 ( .IN1(s0_msel_gnt_p2[2]), .IN2(n11514), .IN3(n3077), .IN4(
        n11515), .Q(n17368) );
  NAND4X0 U34370 ( .IN1(n3184), .IN2(n11516), .IN3(n11517), .IN4(n11518), .QN(
        n11515) );
  OA22X1 U34371 ( .IN1(n11528), .IN2(n18185), .IN3(n11529), .IN4(n3562), .Q(
        n11517) );
  OA221X1 U34372 ( .IN1(n11519), .IN2(n3522), .IN3(n11520), .IN4(n3458), .IN5(
        n11521), .Q(n11518) );
  AO22X1 U34373 ( .IN1(s9_msel_gnt_p1[1]), .IN2(n9781), .IN3(n2941), .IN4(
        n9799), .Q(n17195) );
  NAND3X0 U34374 ( .IN1(n9800), .IN2(n9783), .IN3(n9801), .QN(n9799) );
  OA222X1 U34375 ( .IN1(n9797), .IN2(n3958), .IN3(n9802), .IN4(n3424), .IN5(
        n9803), .IN6(n3215), .Q(n9801) );
  OA21X1 U34376 ( .IN1(n9794), .IN2(n9807), .IN3(n9808), .Q(n9802) );
  AO22X1 U34377 ( .IN1(s9_msel_gnt_p1[0]), .IN2(n9781), .IN3(n2941), .IN4(
        n9816), .Q(n17196) );
  NAND3X0 U34378 ( .IN1(n9800), .IN2(n9817), .IN3(n9818), .QN(n9816) );
  OR2X1 U34379 ( .IN1(n3957), .IN2(n9797), .Q(n9817) );
  OA221X1 U34380 ( .IN1(n3132), .IN2(n9819), .IN3(n18162), .IN4(n9820), .IN5(
        n9790), .Q(n9818) );
  AO22X1 U34381 ( .IN1(s9_msel_gnt_p1[2]), .IN2(n9781), .IN3(n2941), .IN4(
        n9782), .Q(n17194) );
  NAND4X0 U34382 ( .IN1(n3133), .IN2(n9783), .IN3(n9784), .IN4(n9785), .QN(
        n9782) );
  OA22X1 U34383 ( .IN1(n9796), .IN2(n18162), .IN3(n9797), .IN4(n3959), .Q(
        n9784) );
  OA221X1 U34384 ( .IN1(n9786), .IN2(n3488), .IN3(n9787), .IN4(n3424), .IN5(
        n9788), .Q(n9785) );
  AO22X1 U34385 ( .IN1(s9_msel_gnt_p2_1_), .IN2(n9656), .IN3(n2933), .IN4(
        n9673), .Q(n17189) );
  NAND3X0 U34386 ( .IN1(n9674), .IN2(n9658), .IN3(n9675), .QN(n9673) );
  OA222X1 U34387 ( .IN1(n9671), .IN2(n3966), .IN3(n9676), .IN4(n3422), .IN5(
        n9677), .IN6(n3213), .Q(n9675) );
  OA21X1 U34388 ( .IN1(n9669), .IN2(n9681), .IN3(n9682), .Q(n9676) );
  AO22X1 U34389 ( .IN1(s9_msel_gnt_p2_0_), .IN2(n9656), .IN3(n2933), .IN4(
        n9687), .Q(n17190) );
  NAND3X0 U34390 ( .IN1(n9674), .IN2(n9688), .IN3(n9689), .QN(n9687) );
  OR2X1 U34391 ( .IN1(n3965), .IN2(n9671), .Q(n9688) );
  OA221X1 U34392 ( .IN1(n3129), .IN2(n9690), .IN3(n18186), .IN4(n9691), .IN5(
        n9665), .Q(n9689) );
  AO22X1 U34393 ( .IN1(test_so76), .IN2(n9656), .IN3(n2933), .IN4(n9657), .Q(
        n17188) );
  NAND4X0 U34394 ( .IN1(n3130), .IN2(n9658), .IN3(n9659), .IN4(n9660), .QN(
        n9657) );
  OA22X1 U34395 ( .IN1(n9670), .IN2(n18186), .IN3(n9671), .IN4(n3967), .Q(
        n9659) );
  OA221X1 U34396 ( .IN1(n9661), .IN2(n3486), .IN3(n9662), .IN4(n3422), .IN5(
        n9663), .Q(n9660) );
  AO22X1 U34397 ( .IN1(s8_msel_gnt_p1[1]), .IN2(n9470), .IN3(n2957), .IN4(
        n9488), .Q(n17165) );
  NAND3X0 U34398 ( .IN1(n9489), .IN2(n9472), .IN3(n9490), .QN(n9488) );
  OA222X1 U34399 ( .IN1(n9486), .IN2(n3913), .IN3(n9491), .IN4(n3428), .IN5(
        n9492), .IN6(n3219), .Q(n9490) );
  OA21X1 U34400 ( .IN1(n9483), .IN2(n9496), .IN3(n9497), .Q(n9491) );
  AO22X1 U34401 ( .IN1(s8_msel_gnt_p1[0]), .IN2(n9470), .IN3(n2957), .IN4(
        n9505), .Q(n17166) );
  NAND3X0 U34402 ( .IN1(n9489), .IN2(n9506), .IN3(n9507), .QN(n9505) );
  OR2X1 U34403 ( .IN1(n3912), .IN2(n9486), .Q(n9506) );
  OA221X1 U34404 ( .IN1(n3138), .IN2(n9508), .IN3(n18187), .IN4(n9509), .IN5(
        n9479), .Q(n9507) );
  AO22X1 U34405 ( .IN1(s8_msel_gnt_p1[2]), .IN2(n9470), .IN3(n2957), .IN4(
        n9471), .Q(n17164) );
  NAND4X0 U34406 ( .IN1(n3139), .IN2(n9472), .IN3(n9473), .IN4(n9474), .QN(
        n9471) );
  OA22X1 U34407 ( .IN1(n9485), .IN2(n18187), .IN3(n9486), .IN4(n3914), .Q(
        n9473) );
  OA221X1 U34408 ( .IN1(n9475), .IN2(n3492), .IN3(n9476), .IN4(n3428), .IN5(
        n9477), .Q(n9474) );
  AO22X1 U34409 ( .IN1(test_so72), .IN2(n9345), .IN3(n2949), .IN4(n9362), .Q(
        n17159) );
  NAND3X0 U34410 ( .IN1(n9363), .IN2(n9347), .IN3(n9364), .QN(n9362) );
  OA222X1 U34411 ( .IN1(n9360), .IN2(n3921), .IN3(n9365), .IN4(n3426), .IN5(
        n9366), .IN6(n3217), .Q(n9364) );
  OA21X1 U34412 ( .IN1(n9358), .IN2(n9370), .IN3(n9371), .Q(n9365) );
  AO22X1 U34413 ( .IN1(s8_msel_gnt_p2_0_), .IN2(n9345), .IN3(n2949), .IN4(
        n9376), .Q(n17160) );
  NAND3X0 U34414 ( .IN1(n9363), .IN2(n9377), .IN3(n9378), .QN(n9376) );
  OR2X1 U34415 ( .IN1(n3920), .IN2(n9360), .Q(n9377) );
  OA221X1 U34416 ( .IN1(n3135), .IN2(n9379), .IN3(n18188), .IN4(n9380), .IN5(
        n9354), .Q(n9378) );
  AO22X1 U34417 ( .IN1(s8_msel_gnt_p2_2_), .IN2(n9345), .IN3(n2949), .IN4(
        n9346), .Q(n17158) );
  NAND4X0 U34418 ( .IN1(n3136), .IN2(n9347), .IN3(n9348), .IN4(n9349), .QN(
        n9346) );
  OA22X1 U34419 ( .IN1(n9359), .IN2(n18188), .IN3(n9360), .IN4(n3922), .Q(
        n9348) );
  OA221X1 U34420 ( .IN1(n9350), .IN2(n3490), .IN3(n9351), .IN4(n3426), .IN5(
        n9352), .Q(n9349) );
  AO22X1 U34421 ( .IN1(s15_msel_gnt_p0_1_), .IN2(n14001), .IN3(n2837), .IN4(
        n14023), .Q(n17610) );
  NAND3X0 U34422 ( .IN1(n14024), .IN2(n14010), .IN3(n14025), .QN(n14023) );
  OA222X1 U34423 ( .IN1(n14007), .IN2(n4220), .IN3(n14026), .IN4(n3398), .IN5(
        n14027), .IN6(n3189), .Q(n14025) );
  OA21X1 U34424 ( .IN1(n14028), .IN2(n14029), .IN3(n14030), .Q(n14027) );
  AO22X1 U34425 ( .IN1(s15_msel_gnt_p0_0_), .IN2(n14001), .IN3(n2837), .IN4(
        n14040), .Q(n17611) );
  NAND3X0 U34426 ( .IN1(n14024), .IN2(n14041), .IN3(n14042), .QN(n14040) );
  OR2X1 U34427 ( .IN1(n4219), .IN2(n14007), .Q(n14041) );
  AO22X1 U34428 ( .IN1(test_so98), .IN2(n14001), .IN3(n2837), .IN4(n14002), 
        .Q(n17609) );
  NAND4X0 U34429 ( .IN1(n14003), .IN2(n14004), .IN3(n14005), .IN4(n14006), 
        .QN(n14002) );
  NAND3X0 U34430 ( .IN1(n14019), .IN2(n3254), .IN3(n14020), .QN(n14003) );
  AOI22X1 U34431 ( .IN1(test_so36), .IN2(n18820), .IN3(s15_data_i[0]), .IN4(
        n18819), .QN(n14808) );
  AOI22X1 U34432 ( .IN1(rf_rf_dout_1_), .IN2(n18820), .IN3(s15_data_i[1]), 
        .IN4(n18819), .QN(n14709) );
  AOI22X1 U34433 ( .IN1(rf_rf_dout_2_), .IN2(n18820), .IN3(s15_data_i[2]), 
        .IN4(n18819), .QN(n14610) );
  AOI22X1 U34434 ( .IN1(rf_rf_dout_3_), .IN2(n17780), .IN3(s15_data_i[3]), 
        .IN4(n18819), .QN(n14583) );
  AOI22X1 U34435 ( .IN1(rf_rf_dout_4_), .IN2(n18820), .IN3(s15_data_i[4]), 
        .IN4(n18819), .QN(n14574) );
  AOI22X1 U34436 ( .IN1(rf_rf_dout_5_), .IN2(n17780), .IN3(s15_data_i[5]), 
        .IN4(n18818), .QN(n14565) );
  AOI22X1 U34437 ( .IN1(test_so37), .IN2(n18820), .IN3(s15_data_i[6]), .IN4(
        n18819), .QN(n14556) );
  AOI22X1 U34438 ( .IN1(rf_rf_dout_7_), .IN2(n17780), .IN3(s15_data_i[7]), 
        .IN4(n18818), .QN(n14547) );
  AOI22X1 U34439 ( .IN1(rf_rf_dout_8_), .IN2(n17780), .IN3(s15_data_i[8]), 
        .IN4(n18819), .QN(n14538) );
  AOI22X1 U34440 ( .IN1(rf_rf_dout_9_), .IN2(n17780), .IN3(s15_data_i[9]), 
        .IN4(n18819), .QN(n14514) );
  AOI22X1 U34441 ( .IN1(rf_rf_dout_10_), .IN2(n17780), .IN3(s15_data_i[10]), 
        .IN4(n18816), .QN(n14799) );
  AOI22X1 U34442 ( .IN1(rf_rf_dout_11_), .IN2(n17780), .IN3(s15_data_i[11]), 
        .IN4(n18819), .QN(n14790) );
  AOI22X1 U34443 ( .IN1(test_so38), .IN2(n17780), .IN3(s15_data_i[12]), .IN4(
        n18819), .QN(n14781) );
  AOI22X1 U34444 ( .IN1(rf_rf_dout_13_), .IN2(n18820), .IN3(s15_data_i[13]), 
        .IN4(n18819), .QN(n14772) );
  AOI22X1 U34445 ( .IN1(rf_rf_dout_14_), .IN2(n18820), .IN3(s15_data_i[14]), 
        .IN4(n18819), .QN(n14763) );
  AOI22X1 U34446 ( .IN1(rf_rf_dout_15_), .IN2(n18820), .IN3(s15_data_i[15]), 
        .IN4(n18819), .QN(n14754) );
  AOI22X1 U34447 ( .IN1(rf_rf_ack), .IN2(n17780), .IN3(s15_ack_i), .IN4(n18817), .QN(n14851) );
  NOR2X0 U34448 ( .IN1(n17095), .IN2(n17096), .QN(n17764) );
  NAND4X0 U34449 ( .IN1(n17097), .IN2(n17098), .IN3(n17099), .IN4(n17100), 
        .QN(n17096) );
  NAND4X0 U34450 ( .IN1(n17101), .IN2(n17102), .IN3(n17103), .IN4(n17104), 
        .QN(n17095) );
  NAND3X0 U34451 ( .IN1(m1s15_cyc), .IN2(n19645), .IN3(s15_m1_cyc_r), .QN(
        n17098) );
  NAND2X0 U34452 ( .IN1(s15_data_i[16]), .IN2(n18818), .QN(n14745) );
  NAND2X0 U34453 ( .IN1(s15_data_i[17]), .IN2(n18818), .QN(n14736) );
  NAND2X0 U34454 ( .IN1(s15_data_i[19]), .IN2(n18818), .QN(n14718) );
  NAND2X0 U34455 ( .IN1(s15_data_i[20]), .IN2(n18818), .QN(n14700) );
  NAND2X0 U34456 ( .IN1(s15_data_i[21]), .IN2(n18818), .QN(n14691) );
  NAND2X0 U34457 ( .IN1(s15_data_i[23]), .IN2(n18818), .QN(n14673) );
  NAND2X0 U34458 ( .IN1(s15_data_i[24]), .IN2(n18818), .QN(n14664) );
  NAND2X0 U34459 ( .IN1(s15_data_i[25]), .IN2(n18818), .QN(n14655) );
  NAND2X0 U34460 ( .IN1(s15_data_i[18]), .IN2(n18817), .QN(n14727) );
  NAND2X0 U34461 ( .IN1(s15_data_i[22]), .IN2(n18817), .QN(n14682) );
  NAND2X0 U34462 ( .IN1(s15_data_i[26]), .IN2(n18817), .QN(n14646) );
  NAND2X0 U34463 ( .IN1(s15_data_i[27]), .IN2(n18817), .QN(n14637) );
  NAND2X0 U34464 ( .IN1(s15_data_i[28]), .IN2(n18817), .QN(n14628) );
  NAND2X0 U34465 ( .IN1(s15_data_i[29]), .IN2(n18817), .QN(n14619) );
  NAND2X0 U34466 ( .IN1(s15_data_i[30]), .IN2(n18817), .QN(n14601) );
  NAND2X0 U34467 ( .IN1(s15_data_i[31]), .IN2(n18817), .QN(n14592) );
  NAND2X0 U34468 ( .IN1(s15_rty_i), .IN2(n18816), .QN(n14497) );
  NAND2X0 U34469 ( .IN1(s15_err_i), .IN2(n18817), .QN(n14506) );
  NAND3X0 U34470 ( .IN1(conf7_9_), .IN2(n18333), .IN3(conf7_8_), .QN(n13913)
         );
  NAND3X0 U34471 ( .IN1(conf6_9_), .IN2(n18332), .IN3(conf6_8_), .QN(n13604)
         );
  NAND3X0 U34472 ( .IN1(conf14_9_), .IN2(n18331), .IN3(conf14_8_), .QN(n11438)
         );
  NAND3X0 U34473 ( .IN1(conf5_9_), .IN2(n18330), .IN3(conf5_8_), .QN(n13295)
         );
  NAND3X0 U34474 ( .IN1(conf4_9_), .IN2(n18329), .IN3(conf4_8_), .QN(n12986)
         );
  NAND3X0 U34475 ( .IN1(conf13_9_), .IN2(n18328), .IN3(conf13_8_), .QN(n11129)
         );
  NAND3X0 U34476 ( .IN1(conf12_9_), .IN2(n18327), .IN3(conf12_8_), .QN(n10819)
         );
  NAND3X0 U34477 ( .IN1(conf3_9_), .IN2(n18326), .IN3(conf3_8_), .QN(n12677)
         );
  NAND3X0 U34478 ( .IN1(conf2_9_), .IN2(n18325), .IN3(conf2_8_), .QN(n12368)
         );
  NAND3X0 U34479 ( .IN1(conf11_9_), .IN2(n18324), .IN3(conf11_8_), .QN(n10510)
         );
  NAND3X0 U34480 ( .IN1(conf10_9_), .IN2(n18323), .IN3(conf10_8_), .QN(n10200)
         );
  NAND3X0 U34481 ( .IN1(conf1_9_), .IN2(n18322), .IN3(conf1_8_), .QN(n12058)
         );
  NAND3X0 U34482 ( .IN1(conf0_9_), .IN2(n18321), .IN3(conf0_8_), .QN(n11748)
         );
  NAND3X0 U34483 ( .IN1(conf9_9_), .IN2(n18320), .IN3(conf9_8_), .QN(n9890) );
  NAND3X0 U34484 ( .IN1(conf8_9_), .IN2(n18319), .IN3(conf8_8_), .QN(n9579) );
  OA221X1 U34485 ( .IN1(n13874), .IN2(n3885), .IN3(n13875), .IN4(n13876), 
        .IN5(n13877), .Q(n13873) );
  ISOLANDX1 U34486 ( .D(n13878), .ISO(n13879), .Q(n13877) );
  OA221X1 U34487 ( .IN1(n13565), .IN2(n3840), .IN3(n13566), .IN4(n13567), 
        .IN5(n13568), .Q(n13564) );
  ISOLANDX1 U34488 ( .D(n13569), .ISO(n13570), .Q(n13568) );
  OA221X1 U34489 ( .IN1(n11399), .IN2(n4200), .IN3(n11400), .IN4(n11401), 
        .IN5(n11402), .Q(n11398) );
  ISOLANDX1 U34490 ( .D(n11403), .ISO(n11404), .Q(n11402) );
  OA221X1 U34491 ( .IN1(n13256), .IN2(n3795), .IN3(n13257), .IN4(n13258), 
        .IN5(n13259), .Q(n13255) );
  ISOLANDX1 U34492 ( .D(n13260), .ISO(n13261), .Q(n13259) );
  OA221X1 U34493 ( .IN1(n12947), .IN2(n3750), .IN3(n12948), .IN4(n12949), 
        .IN5(n12950), .Q(n12946) );
  ISOLANDX1 U34494 ( .D(n12951), .ISO(n12952), .Q(n12950) );
  OA221X1 U34495 ( .IN1(n11090), .IN2(n4155), .IN3(n11091), .IN4(n11092), 
        .IN5(n11093), .Q(n11089) );
  ISOLANDX1 U34496 ( .D(n11094), .ISO(n11095), .Q(n11093) );
  OA221X1 U34497 ( .IN1(n10780), .IN2(n4110), .IN3(n10781), .IN4(n10782), 
        .IN5(n10783), .Q(n10779) );
  ISOLANDX1 U34498 ( .D(n10784), .ISO(n10785), .Q(n10783) );
  OA221X1 U34499 ( .IN1(n12638), .IN2(n3705), .IN3(n12639), .IN4(n12640), 
        .IN5(n12641), .Q(n12637) );
  ISOLANDX1 U34500 ( .D(n12642), .ISO(n12643), .Q(n12641) );
  OA221X1 U34501 ( .IN1(n12329), .IN2(n3660), .IN3(n12330), .IN4(n12331), 
        .IN5(n12332), .Q(n12328) );
  ISOLANDX1 U34502 ( .D(n12333), .ISO(n12334), .Q(n12332) );
  OA221X1 U34503 ( .IN1(n10471), .IN2(n4065), .IN3(n10472), .IN4(n10473), 
        .IN5(n10474), .Q(n10470) );
  ISOLANDX1 U34504 ( .D(n10475), .ISO(n10476), .Q(n10474) );
  OA221X1 U34505 ( .IN1(n10161), .IN2(n4020), .IN3(n10162), .IN4(n10163), 
        .IN5(n10164), .Q(n10160) );
  ISOLANDX1 U34506 ( .D(n10165), .ISO(n10166), .Q(n10164) );
  OA221X1 U34507 ( .IN1(n12019), .IN2(n3615), .IN3(n12020), .IN4(n12021), 
        .IN5(n12022), .Q(n12018) );
  ISOLANDX1 U34508 ( .D(n12023), .ISO(n12024), .Q(n12022) );
  OA221X1 U34509 ( .IN1(n11709), .IN2(n3570), .IN3(n11710), .IN4(n11711), 
        .IN5(n11712), .Q(n11708) );
  ISOLANDX1 U34510 ( .D(n11713), .ISO(n11714), .Q(n11712) );
  OA221X1 U34511 ( .IN1(n9851), .IN2(n3975), .IN3(n9852), .IN4(n9853), .IN5(
        n9854), .Q(n9850) );
  ISOLANDX1 U34512 ( .D(n9855), .ISO(n9856), .Q(n9854) );
  OA221X1 U34513 ( .IN1(n9540), .IN2(n3930), .IN3(n9541), .IN4(n9542), .IN5(
        n9543), .Q(n9539) );
  ISOLANDX1 U34514 ( .D(n9544), .ISO(n9545), .Q(n9543) );
  OA221X1 U34515 ( .IN1(n14148), .IN2(n4245), .IN3(n14149), .IN4(n14150), 
        .IN5(n14151), .Q(n14147) );
  ISOLANDX1 U34516 ( .D(n14152), .ISO(n14153), .Q(n14151) );
  AO22X1 U34517 ( .IN1(s7_msel_gnt_p3[1]), .IN2(n13868), .IN3(n2977), .IN4(
        n13889), .Q(n17588) );
  NAND3X0 U34518 ( .IN1(n13890), .IN2(n13878), .IN3(n13891), .QN(n13889) );
  OA222X1 U34519 ( .IN1(n13874), .IN2(n3884), .IN3(n13892), .IN4(n13883), 
        .IN5(n13893), .IN6(n13894), .Q(n13891) );
  OA21X1 U34520 ( .IN1(n13886), .IN2(n13898), .IN3(n13899), .Q(n13892) );
  AO22X1 U34521 ( .IN1(s7_msel_gnt_p3[2]), .IN2(n13868), .IN3(n2977), .IN4(
        n13869), .Q(n17587) );
  NAND4X0 U34522 ( .IN1(n13870), .IN2(n13871), .IN3(n13872), .IN4(n13873), 
        .QN(n13869) );
  NAND3X0 U34523 ( .IN1(n13887), .IN2(n13888), .IN3(n3390), .QN(n13870) );
  OA22X1 U34524 ( .IN1(n13880), .IN2(n13881), .IN3(n13882), .IN4(n13883), .Q(
        n13872) );
  AO22X1 U34525 ( .IN1(s7_msel_gnt_p3[0]), .IN2(n13868), .IN3(n2977), .IN4(
        n13904), .Q(n17589) );
  NAND3X0 U34526 ( .IN1(n13890), .IN2(n13905), .IN3(n13906), .QN(n13904) );
  OR2X1 U34527 ( .IN1(n3883), .IN2(n13874), .Q(n13905) );
  OA221X1 U34528 ( .IN1(n13907), .IN2(n13908), .IN3(n13909), .IN4(n13910), 
        .IN5(n13871), .Q(n13906) );
  AO22X1 U34529 ( .IN1(s6_msel_gnt_p3_1_), .IN2(n13559), .IN3(n2993), .IN4(
        n13580), .Q(n17558) );
  NAND3X0 U34530 ( .IN1(n13581), .IN2(n13569), .IN3(n13582), .QN(n13580) );
  OA222X1 U34531 ( .IN1(n13565), .IN2(n3839), .IN3(n13583), .IN4(n13574), 
        .IN5(n13584), .IN6(n13585), .Q(n13582) );
  OA21X1 U34532 ( .IN1(n13577), .IN2(n13589), .IN3(n13590), .Q(n13583) );
  AO22X1 U34533 ( .IN1(test_so65), .IN2(n13559), .IN3(n2993), .IN4(n13560), 
        .Q(n17557) );
  NAND4X0 U34534 ( .IN1(n13561), .IN2(n13562), .IN3(n13563), .IN4(n13564), 
        .QN(n13560) );
  NAND3X0 U34535 ( .IN1(n13578), .IN2(n13579), .IN3(n3391), .QN(n13561) );
  OA22X1 U34536 ( .IN1(n13571), .IN2(n13572), .IN3(n13573), .IN4(n13574), .Q(
        n13563) );
  AO22X1 U34537 ( .IN1(s6_msel_gnt_p3_0_), .IN2(n13559), .IN3(n2993), .IN4(
        n13595), .Q(n17559) );
  NAND3X0 U34538 ( .IN1(n13581), .IN2(n13596), .IN3(n13597), .QN(n13595) );
  OR2X1 U34539 ( .IN1(n3838), .IN2(n13565), .Q(n13596) );
  OA221X1 U34540 ( .IN1(n13598), .IN2(n13599), .IN3(n13600), .IN4(n13601), 
        .IN5(n13562), .Q(n13597) );
  AO22X1 U34541 ( .IN1(s14_msel_gnt_p3[1]), .IN2(n11393), .IN3(n2865), .IN4(
        n11414), .Q(n17348) );
  NAND3X0 U34542 ( .IN1(n11415), .IN2(n11403), .IN3(n11416), .QN(n11414) );
  OA222X1 U34543 ( .IN1(n11399), .IN2(n4199), .IN3(n11417), .IN4(n11408), 
        .IN5(n11418), .IN6(n11419), .Q(n11416) );
  OA21X1 U34544 ( .IN1(n11411), .IN2(n11423), .IN3(n11424), .Q(n11417) );
  AO22X1 U34545 ( .IN1(s14_msel_gnt_p3[2]), .IN2(n11393), .IN3(n2865), .IN4(
        n11394), .Q(n17347) );
  NAND4X0 U34546 ( .IN1(n11395), .IN2(n11396), .IN3(n11397), .IN4(n11398), 
        .QN(n11394) );
  NAND3X0 U34547 ( .IN1(n11412), .IN2(n11413), .IN3(n3383), .QN(n11395) );
  OA22X1 U34548 ( .IN1(n11405), .IN2(n11406), .IN3(n11407), .IN4(n11408), .Q(
        n11397) );
  AO22X1 U34549 ( .IN1(s14_msel_gnt_p3[0]), .IN2(n11393), .IN3(n2865), .IN4(
        n11429), .Q(n17349) );
  NAND3X0 U34550 ( .IN1(n11415), .IN2(n11430), .IN3(n11431), .QN(n11429) );
  OR2X1 U34551 ( .IN1(n4198), .IN2(n11399), .Q(n11430) );
  OA221X1 U34552 ( .IN1(n11432), .IN2(n11433), .IN3(n11434), .IN4(n11435), 
        .IN5(n11396), .Q(n11431) );
  AO22X1 U34553 ( .IN1(test_so61), .IN2(n13250), .IN3(n3009), .IN4(n13271), 
        .Q(n17528) );
  NAND3X0 U34554 ( .IN1(n13272), .IN2(n13260), .IN3(n13273), .QN(n13271) );
  OA222X1 U34555 ( .IN1(n13256), .IN2(n3794), .IN3(n13274), .IN4(n13265), 
        .IN5(n13275), .IN6(n13276), .Q(n13273) );
  OA21X1 U34556 ( .IN1(n13268), .IN2(n13280), .IN3(n13281), .Q(n13274) );
  AO22X1 U34557 ( .IN1(s5_msel_gnt_p3_2_), .IN2(n13250), .IN3(n3009), .IN4(
        n13251), .Q(n17527) );
  NAND4X0 U34558 ( .IN1(n13252), .IN2(n13253), .IN3(n13254), .IN4(n13255), 
        .QN(n13251) );
  NAND3X0 U34559 ( .IN1(n13269), .IN2(n13270), .IN3(n3392), .QN(n13252) );
  OA22X1 U34560 ( .IN1(n13262), .IN2(n13263), .IN3(n13264), .IN4(n13265), .Q(
        n13254) );
  AO22X1 U34561 ( .IN1(s5_msel_gnt_p3_0_), .IN2(n13250), .IN3(n3009), .IN4(
        n13286), .Q(n17529) );
  NAND3X0 U34562 ( .IN1(n13272), .IN2(n13287), .IN3(n13288), .QN(n13286) );
  OR2X1 U34563 ( .IN1(n3793), .IN2(n13256), .Q(n13287) );
  OA221X1 U34564 ( .IN1(n13289), .IN2(n13290), .IN3(n13291), .IN4(n13292), 
        .IN5(n13253), .Q(n13288) );
  AO22X1 U34565 ( .IN1(s4_msel_gnt_p3_1_), .IN2(n12941), .IN3(n3025), .IN4(
        n12962), .Q(n17498) );
  NAND3X0 U34566 ( .IN1(n12963), .IN2(n12951), .IN3(n12964), .QN(n12962) );
  OA222X1 U34567 ( .IN1(n12947), .IN2(n3749), .IN3(n12965), .IN4(n12956), 
        .IN5(n12966), .IN6(n12967), .Q(n12964) );
  OA21X1 U34568 ( .IN1(n12959), .IN2(n12971), .IN3(n12972), .Q(n12965) );
  AO22X1 U34569 ( .IN1(s4_msel_gnt_p3_2_), .IN2(n12941), .IN3(n3025), .IN4(
        n12942), .Q(n17497) );
  NAND4X0 U34570 ( .IN1(n12943), .IN2(n12944), .IN3(n12945), .IN4(n12946), 
        .QN(n12942) );
  NAND3X0 U34571 ( .IN1(n12960), .IN2(n12961), .IN3(n3393), .QN(n12943) );
  OA22X1 U34572 ( .IN1(n12953), .IN2(n12954), .IN3(n12955), .IN4(n12956), .Q(
        n12945) );
  AO22X1 U34573 ( .IN1(test_so57), .IN2(n12941), .IN3(n3025), .IN4(n12977), 
        .Q(n17499) );
  NAND3X0 U34574 ( .IN1(n12963), .IN2(n12978), .IN3(n12979), .QN(n12977) );
  OR2X1 U34575 ( .IN1(n3748), .IN2(n12947), .Q(n12978) );
  OA221X1 U34576 ( .IN1(n12980), .IN2(n12981), .IN3(n12982), .IN4(n12983), 
        .IN5(n12944), .Q(n12979) );
  AO22X1 U34577 ( .IN1(s13_msel_gnt_p3[1]), .IN2(n11084), .IN3(n2881), .IN4(
        n11105), .Q(n17318) );
  NAND3X0 U34578 ( .IN1(n11106), .IN2(n11094), .IN3(n11107), .QN(n11105) );
  OA222X1 U34579 ( .IN1(n11090), .IN2(n4154), .IN3(n11108), .IN4(n11099), 
        .IN5(n11109), .IN6(n11110), .Q(n11107) );
  OA21X1 U34580 ( .IN1(n11102), .IN2(n11114), .IN3(n11115), .Q(n11108) );
  AO22X1 U34581 ( .IN1(s13_msel_gnt_p3[2]), .IN2(n11084), .IN3(n2881), .IN4(
        n11085), .Q(n17317) );
  NAND4X0 U34582 ( .IN1(n11086), .IN2(n11087), .IN3(n11088), .IN4(n11089), 
        .QN(n11085) );
  NAND3X0 U34583 ( .IN1(n11103), .IN2(n11104), .IN3(n3384), .QN(n11086) );
  OA22X1 U34584 ( .IN1(n11096), .IN2(n11097), .IN3(n11098), .IN4(n11099), .Q(
        n11088) );
  AO22X1 U34585 ( .IN1(s13_msel_gnt_p3[0]), .IN2(n11084), .IN3(n2881), .IN4(
        n11120), .Q(n17319) );
  NAND3X0 U34586 ( .IN1(n11106), .IN2(n11121), .IN3(n11122), .QN(n11120) );
  OR2X1 U34587 ( .IN1(n4153), .IN2(n11090), .Q(n11121) );
  OA221X1 U34588 ( .IN1(n11123), .IN2(n11124), .IN3(n11125), .IN4(n11126), 
        .IN5(n11087), .Q(n11122) );
  AO22X1 U34589 ( .IN1(s12_msel_gnt_p3_1_), .IN2(n10774), .IN3(n2897), .IN4(
        n10795), .Q(n17288) );
  NAND3X0 U34590 ( .IN1(n10796), .IN2(n10784), .IN3(n10797), .QN(n10795) );
  OA222X1 U34591 ( .IN1(n10780), .IN2(n4109), .IN3(n10798), .IN4(n10789), 
        .IN5(n10799), .IN6(n10800), .Q(n10797) );
  OA21X1 U34592 ( .IN1(n10792), .IN2(n10804), .IN3(n10805), .Q(n10798) );
  AO22X1 U34593 ( .IN1(test_so88), .IN2(n10774), .IN3(n2897), .IN4(n10775), 
        .Q(n17287) );
  NAND4X0 U34594 ( .IN1(n10776), .IN2(n10777), .IN3(n10778), .IN4(n10779), 
        .QN(n10775) );
  NAND3X0 U34595 ( .IN1(n10793), .IN2(n10794), .IN3(n3385), .QN(n10776) );
  OA22X1 U34596 ( .IN1(n10786), .IN2(n10787), .IN3(n10788), .IN4(n10789), .Q(
        n10778) );
  AO22X1 U34597 ( .IN1(s12_msel_gnt_p3_0_), .IN2(n10774), .IN3(n2897), .IN4(
        n10810), .Q(n17289) );
  NAND3X0 U34598 ( .IN1(n10796), .IN2(n10811), .IN3(n10812), .QN(n10810) );
  OR2X1 U34599 ( .IN1(n4108), .IN2(n10780), .Q(n10811) );
  OA221X1 U34600 ( .IN1(n10813), .IN2(n10814), .IN3(n10815), .IN4(n10816), 
        .IN5(n10777), .Q(n10812) );
  AO22X1 U34601 ( .IN1(s3_msel_gnt_p3[1]), .IN2(n12632), .IN3(n3041), .IN4(
        n12653), .Q(n17468) );
  NAND3X0 U34602 ( .IN1(n12654), .IN2(n12642), .IN3(n12655), .QN(n12653) );
  OA222X1 U34603 ( .IN1(n12638), .IN2(n3704), .IN3(n12656), .IN4(n12647), 
        .IN5(n12657), .IN6(n12658), .Q(n12655) );
  OA21X1 U34604 ( .IN1(n12650), .IN2(n12662), .IN3(n12663), .Q(n12656) );
  AO22X1 U34605 ( .IN1(s3_msel_gnt_p3[2]), .IN2(n12632), .IN3(n3041), .IN4(
        n12633), .Q(n17467) );
  NAND4X0 U34606 ( .IN1(n12634), .IN2(n12635), .IN3(n12636), .IN4(n12637), 
        .QN(n12633) );
  NAND3X0 U34607 ( .IN1(n12651), .IN2(n12652), .IN3(n3394), .QN(n12634) );
  OA22X1 U34608 ( .IN1(n12644), .IN2(n12645), .IN3(n12646), .IN4(n12647), .Q(
        n12636) );
  AO22X1 U34609 ( .IN1(s3_msel_gnt_p3[0]), .IN2(n12632), .IN3(n3041), .IN4(
        n12668), .Q(n17469) );
  NAND3X0 U34610 ( .IN1(n12654), .IN2(n12669), .IN3(n12670), .QN(n12668) );
  OR2X1 U34611 ( .IN1(n3703), .IN2(n12638), .Q(n12669) );
  OA221X1 U34612 ( .IN1(n12671), .IN2(n12672), .IN3(n12673), .IN4(n12674), 
        .IN5(n12635), .Q(n12670) );
  AO22X1 U34613 ( .IN1(s2_msel_gnt_p3[1]), .IN2(n12323), .IN3(n3057), .IN4(
        n12344), .Q(n17438) );
  NAND3X0 U34614 ( .IN1(n12345), .IN2(n12333), .IN3(n12346), .QN(n12344) );
  OA222X1 U34615 ( .IN1(n12329), .IN2(n3659), .IN3(n12347), .IN4(n12338), 
        .IN5(n12348), .IN6(n12349), .Q(n12346) );
  OA21X1 U34616 ( .IN1(n12341), .IN2(n12353), .IN3(n12354), .Q(n12347) );
  AO22X1 U34617 ( .IN1(s2_msel_gnt_p3[2]), .IN2(n12323), .IN3(n3057), .IN4(
        n12324), .Q(n17437) );
  NAND4X0 U34618 ( .IN1(n12325), .IN2(n12326), .IN3(n12327), .IN4(n12328), 
        .QN(n12324) );
  NAND3X0 U34619 ( .IN1(n12342), .IN2(n12343), .IN3(n3395), .QN(n12325) );
  OA22X1 U34620 ( .IN1(n12335), .IN2(n12336), .IN3(n12337), .IN4(n12338), .Q(
        n12327) );
  AO22X1 U34621 ( .IN1(s2_msel_gnt_p3[0]), .IN2(n12323), .IN3(n3057), .IN4(
        n12359), .Q(n17439) );
  NAND3X0 U34622 ( .IN1(n12345), .IN2(n12360), .IN3(n12361), .QN(n12359) );
  OR2X1 U34623 ( .IN1(n3658), .IN2(n12329), .Q(n12360) );
  OA221X1 U34624 ( .IN1(n12362), .IN2(n12363), .IN3(n12364), .IN4(n12365), 
        .IN5(n12326), .Q(n12361) );
  AO22X1 U34625 ( .IN1(test_so84), .IN2(n10465), .IN3(n2913), .IN4(n10486), 
        .Q(n17258) );
  NAND3X0 U34626 ( .IN1(n10487), .IN2(n10475), .IN3(n10488), .QN(n10486) );
  OA222X1 U34627 ( .IN1(n10471), .IN2(n4064), .IN3(n10489), .IN4(n10480), 
        .IN5(n10490), .IN6(n10491), .Q(n10488) );
  OA21X1 U34628 ( .IN1(n10483), .IN2(n10495), .IN3(n10496), .Q(n10489) );
  AO22X1 U34629 ( .IN1(s11_msel_gnt_p3_2_), .IN2(n10465), .IN3(n2913), .IN4(
        n10466), .Q(n17257) );
  NAND4X0 U34630 ( .IN1(n10467), .IN2(n10468), .IN3(n10469), .IN4(n10470), 
        .QN(n10466) );
  NAND3X0 U34631 ( .IN1(n10484), .IN2(n10485), .IN3(n3386), .QN(n10467) );
  OA22X1 U34632 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .IN4(n10480), .Q(
        n10469) );
  AO22X1 U34633 ( .IN1(s11_msel_gnt_p3_0_), .IN2(n10465), .IN3(n2913), .IN4(
        n10501), .Q(n17259) );
  NAND3X0 U34634 ( .IN1(n10487), .IN2(n10502), .IN3(n10503), .QN(n10501) );
  OR2X1 U34635 ( .IN1(n4063), .IN2(n10471), .Q(n10502) );
  OA221X1 U34636 ( .IN1(n10504), .IN2(n10505), .IN3(n10506), .IN4(n10507), 
        .IN5(n10468), .Q(n10503) );
  AO22X1 U34637 ( .IN1(s10_msel_gnt_p3_1_), .IN2(n10155), .IN3(n2929), .IN4(
        n10176), .Q(n17228) );
  NAND3X0 U34638 ( .IN1(n10177), .IN2(n10165), .IN3(n10178), .QN(n10176) );
  OA222X1 U34639 ( .IN1(n10161), .IN2(n4019), .IN3(n10179), .IN4(n10170), 
        .IN5(n10180), .IN6(n10181), .Q(n10178) );
  OA21X1 U34640 ( .IN1(n10173), .IN2(n10185), .IN3(n10186), .Q(n10179) );
  AO22X1 U34641 ( .IN1(s10_msel_gnt_p3_2_), .IN2(n10155), .IN3(n2929), .IN4(
        n10156), .Q(n17227) );
  NAND4X0 U34642 ( .IN1(n10157), .IN2(n10158), .IN3(n10159), .IN4(n10160), 
        .QN(n10156) );
  NAND3X0 U34643 ( .IN1(n10174), .IN2(n10175), .IN3(n3387), .QN(n10157) );
  OA22X1 U34644 ( .IN1(n10167), .IN2(n10168), .IN3(n10169), .IN4(n10170), .Q(
        n10159) );
  AO22X1 U34645 ( .IN1(test_so80), .IN2(n10155), .IN3(n2929), .IN4(n10191), 
        .Q(n17229) );
  NAND3X0 U34646 ( .IN1(n10177), .IN2(n10192), .IN3(n10193), .QN(n10191) );
  OR2X1 U34647 ( .IN1(n4018), .IN2(n10161), .Q(n10192) );
  OA221X1 U34648 ( .IN1(n10194), .IN2(n10195), .IN3(n10196), .IN4(n10197), 
        .IN5(n10158), .Q(n10193) );
  AO22X1 U34649 ( .IN1(s1_msel_gnt_p3[1]), .IN2(n12013), .IN3(n3073), .IN4(
        n12034), .Q(n17408) );
  NAND3X0 U34650 ( .IN1(n12035), .IN2(n12023), .IN3(n12036), .QN(n12034) );
  OA222X1 U34651 ( .IN1(n12019), .IN2(n3614), .IN3(n12037), .IN4(n12028), 
        .IN5(n12038), .IN6(n12039), .Q(n12036) );
  OA21X1 U34652 ( .IN1(n12031), .IN2(n12043), .IN3(n12044), .Q(n12037) );
  AO22X1 U34653 ( .IN1(s1_msel_gnt_p3[2]), .IN2(n12013), .IN3(n3073), .IN4(
        n12014), .Q(n17407) );
  NAND4X0 U34654 ( .IN1(n12015), .IN2(n12016), .IN3(n12017), .IN4(n12018), 
        .QN(n12014) );
  NAND3X0 U34655 ( .IN1(n12032), .IN2(n12033), .IN3(n3396), .QN(n12015) );
  OA22X1 U34656 ( .IN1(n12025), .IN2(n12026), .IN3(n12027), .IN4(n12028), .Q(
        n12017) );
  AO22X1 U34657 ( .IN1(s1_msel_gnt_p3[0]), .IN2(n12013), .IN3(n3073), .IN4(
        n12049), .Q(n17409) );
  NAND3X0 U34658 ( .IN1(n12035), .IN2(n12050), .IN3(n12051), .QN(n12049) );
  OR2X1 U34659 ( .IN1(n3613), .IN2(n12019), .Q(n12050) );
  OA221X1 U34660 ( .IN1(n12052), .IN2(n12053), .IN3(n12054), .IN4(n12055), 
        .IN5(n12016), .Q(n12051) );
  AO22X1 U34661 ( .IN1(s0_msel_gnt_p3_1_), .IN2(n11703), .IN3(n3089), .IN4(
        n11724), .Q(n17378) );
  NAND3X0 U34662 ( .IN1(n11725), .IN2(n11713), .IN3(n11726), .QN(n11724) );
  OA222X1 U34663 ( .IN1(n11709), .IN2(n3569), .IN3(n11727), .IN4(n11718), 
        .IN5(n11728), .IN6(n11729), .Q(n11726) );
  OA21X1 U34664 ( .IN1(n11721), .IN2(n11733), .IN3(n11734), .Q(n11727) );
  AO22X1 U34665 ( .IN1(test_so42), .IN2(n11703), .IN3(n3089), .IN4(n11704), 
        .Q(n17377) );
  NAND4X0 U34666 ( .IN1(n11705), .IN2(n11706), .IN3(n11707), .IN4(n11708), 
        .QN(n11704) );
  NAND3X0 U34667 ( .IN1(n11722), .IN2(n11723), .IN3(n3397), .QN(n11705) );
  OA22X1 U34668 ( .IN1(n11715), .IN2(n11716), .IN3(n11717), .IN4(n11718), .Q(
        n11707) );
  AO22X1 U34669 ( .IN1(s0_msel_gnt_p3_0_), .IN2(n11703), .IN3(n3089), .IN4(
        n11739), .Q(n17379) );
  NAND3X0 U34670 ( .IN1(n11725), .IN2(n11740), .IN3(n11741), .QN(n11739) );
  OR2X1 U34671 ( .IN1(n3568), .IN2(n11709), .Q(n11740) );
  OA221X1 U34672 ( .IN1(n11742), .IN2(n11743), .IN3(n11744), .IN4(n11745), 
        .IN5(n11706), .Q(n11741) );
  AO22X1 U34673 ( .IN1(s9_msel_gnt_p3[1]), .IN2(n9845), .IN3(n2945), .IN4(
        n9866), .Q(n17198) );
  NAND3X0 U34674 ( .IN1(n9867), .IN2(n9855), .IN3(n9868), .QN(n9866) );
  OA222X1 U34675 ( .IN1(n9851), .IN2(n3974), .IN3(n9869), .IN4(n9860), .IN5(
        n9870), .IN6(n9871), .Q(n9868) );
  OA21X1 U34676 ( .IN1(n9863), .IN2(n9875), .IN3(n9876), .Q(n9869) );
  AO22X1 U34677 ( .IN1(s9_msel_gnt_p3[2]), .IN2(n9845), .IN3(n2945), .IN4(
        n9846), .Q(n17197) );
  NAND4X0 U34678 ( .IN1(n9847), .IN2(n9848), .IN3(n9849), .IN4(n9850), .QN(
        n9846) );
  NAND3X0 U34679 ( .IN1(n9864), .IN2(n9865), .IN3(n3388), .QN(n9847) );
  OA22X1 U34680 ( .IN1(n9857), .IN2(n9858), .IN3(n9859), .IN4(n9860), .Q(n9849) );
  AO22X1 U34681 ( .IN1(s9_msel_gnt_p3[0]), .IN2(n9845), .IN3(n2945), .IN4(
        n9881), .Q(n17199) );
  NAND3X0 U34682 ( .IN1(n9867), .IN2(n9882), .IN3(n9883), .QN(n9881) );
  OR2X1 U34683 ( .IN1(n3973), .IN2(n9851), .Q(n9882) );
  OA221X1 U34684 ( .IN1(n9884), .IN2(n9885), .IN3(n9886), .IN4(n9887), .IN5(
        n9848), .Q(n9883) );
  AO22X1 U34685 ( .IN1(s8_msel_gnt_p3[1]), .IN2(n9534), .IN3(n2961), .IN4(
        n9555), .Q(n17168) );
  NAND3X0 U34686 ( .IN1(n9556), .IN2(n9544), .IN3(n9557), .QN(n9555) );
  OA222X1 U34687 ( .IN1(n9540), .IN2(n3929), .IN3(n9558), .IN4(n9549), .IN5(
        n9559), .IN6(n9560), .Q(n9557) );
  OA21X1 U34688 ( .IN1(n9552), .IN2(n9564), .IN3(n9565), .Q(n9558) );
  AO22X1 U34689 ( .IN1(s8_msel_gnt_p3[2]), .IN2(n9534), .IN3(n2961), .IN4(
        n9535), .Q(n17167) );
  NAND4X0 U34690 ( .IN1(n9536), .IN2(n9537), .IN3(n9538), .IN4(n9539), .QN(
        n9535) );
  NAND3X0 U34691 ( .IN1(n9553), .IN2(n9554), .IN3(n3389), .QN(n9536) );
  OA22X1 U34692 ( .IN1(n9546), .IN2(n9547), .IN3(n9548), .IN4(n9549), .Q(n9538) );
  AO22X1 U34693 ( .IN1(s8_msel_gnt_p3[0]), .IN2(n9534), .IN3(n2961), .IN4(
        n9570), .Q(n17169) );
  NAND3X0 U34694 ( .IN1(n9556), .IN2(n9571), .IN3(n9572), .QN(n9570) );
  OR2X1 U34695 ( .IN1(n3928), .IN2(n9540), .Q(n9571) );
  OA221X1 U34696 ( .IN1(n9573), .IN2(n9574), .IN3(n9575), .IN4(n9576), .IN5(
        n9537), .Q(n9572) );
  AO22X1 U34697 ( .IN1(s15_msel_gnt_p1[1]), .IN2(n13935), .IN3(n2843), .IN4(
        n13955), .Q(n17607) );
  NAND3X0 U34698 ( .IN1(n13956), .IN2(n13937), .IN3(n13957), .QN(n13955) );
  OA222X1 U34699 ( .IN1(n13953), .IN2(n4228), .IN3(n13958), .IN4(n3400), .IN5(
        n13959), .IN6(n3191), .Q(n13957) );
  OA21X1 U34700 ( .IN1(n13949), .IN2(n13963), .IN3(n13964), .Q(n13958) );
  AO22X1 U34701 ( .IN1(s15_msel_gnt_p1[0]), .IN2(n13935), .IN3(n2843), .IN4(
        n13972), .Q(n17608) );
  NAND3X0 U34702 ( .IN1(n13956), .IN2(n13973), .IN3(n13974), .QN(n13972) );
  OR2X1 U34703 ( .IN1(n4227), .IN2(n13953), .Q(n13973) );
  OA221X1 U34704 ( .IN1(n3095), .IN2(n13975), .IN3(n18157), .IN4(n13976), 
        .IN5(n13945), .Q(n13974) );
  AO22X1 U34705 ( .IN1(s15_msel_gnt_p1[2]), .IN2(n13935), .IN3(n2843), .IN4(
        n13936), .Q(n17606) );
  NAND4X0 U34706 ( .IN1(n3096), .IN2(n13937), .IN3(n13938), .IN4(n13939), .QN(
        n13936) );
  OA221X1 U34707 ( .IN1(n13940), .IN2(n3464), .IN3(n13941), .IN4(n3400), .IN5(
        n13942), .Q(n13939) );
  OA22X1 U34708 ( .IN1(n13951), .IN2(n18157), .IN3(n13953), .IN4(n4229), .Q(
        n13938) );
  AO22X1 U34709 ( .IN1(s15_msel_gnt_p3[1]), .IN2(n14142), .IN3(n2840), .IN4(
        n14163), .Q(n17616) );
  NAND3X0 U34710 ( .IN1(n14164), .IN2(n14152), .IN3(n14165), .QN(n14163) );
  OA222X1 U34711 ( .IN1(n14148), .IN2(n4244), .IN3(n14166), .IN4(n14157), 
        .IN5(n14167), .IN6(n14168), .Q(n14165) );
  OA21X1 U34712 ( .IN1(n14160), .IN2(n14172), .IN3(n14173), .Q(n14166) );
  AO22X1 U34713 ( .IN1(s15_msel_gnt_p3[2]), .IN2(n14142), .IN3(n2840), .IN4(
        n14143), .Q(n17615) );
  NAND4X0 U34714 ( .IN1(n14144), .IN2(n14145), .IN3(n14146), .IN4(n14147), 
        .QN(n14143) );
  NAND3X0 U34715 ( .IN1(n14161), .IN2(n14162), .IN3(n3381), .QN(n14144) );
  OA22X1 U34716 ( .IN1(n14154), .IN2(n14155), .IN3(n14156), .IN4(n14157), .Q(
        n14146) );
  AO22X1 U34717 ( .IN1(s15_msel_gnt_p3[0]), .IN2(n14142), .IN3(n2840), .IN4(
        n14178), .Q(n17617) );
  NAND3X0 U34718 ( .IN1(n14164), .IN2(n14179), .IN3(n14180), .QN(n14178) );
  OR2X1 U34719 ( .IN1(n4243), .IN2(n14148), .Q(n14179) );
  OA221X1 U34720 ( .IN1(n14181), .IN2(n14182), .IN3(n14183), .IN4(n14184), 
        .IN5(n14145), .Q(n14180) );
  AO22X1 U34721 ( .IN1(s15_msel_gnt_p2_1_), .IN2(n14076), .IN3(n2848), .IN4(
        n14095), .Q(n17613) );
  NAND3X0 U34722 ( .IN1(n14096), .IN2(n14078), .IN3(n14097), .QN(n14095) );
  OA222X1 U34723 ( .IN1(n14093), .IN2(n4236), .IN3(n14098), .IN4(n3401), .IN5(
        n14099), .IN6(n3192), .Q(n14097) );
  OA21X1 U34724 ( .IN1(n14089), .IN2(n14103), .IN3(n14104), .Q(n14098) );
  AO22X1 U34725 ( .IN1(s15_msel_gnt_p2_0_), .IN2(n14076), .IN3(n2848), .IN4(
        n14112), .Q(n17614) );
  NAND3X0 U34726 ( .IN1(n14096), .IN2(n14113), .IN3(n14114), .QN(n14112) );
  OR2X1 U34727 ( .IN1(n4235), .IN2(n14093), .Q(n14113) );
  OA221X1 U34728 ( .IN1(n3097), .IN2(n14115), .IN3(n18158), .IN4(n14116), 
        .IN5(n14085), .Q(n14114) );
  AO22X1 U34729 ( .IN1(test_so99), .IN2(n14076), .IN3(n2848), .IN4(n14077), 
        .Q(n17612) );
  NAND4X0 U34730 ( .IN1(n3098), .IN2(n14078), .IN3(n14079), .IN4(n14080), .QN(
        n14077) );
  OA221X1 U34731 ( .IN1(n14081), .IN2(n3465), .IN3(n14082), .IN4(n3401), .IN5(
        n14083), .Q(n14080) );
  OA22X1 U34732 ( .IN1(n14091), .IN2(n18158), .IN3(n14093), .IN4(n4237), .Q(
        n14079) );
  AO221X1 U34733 ( .IN1(n13632), .IN2(n13629), .IN3(n13627), .IN4(
        s7_msel_pri_out_1_), .IN5(n13628), .Q(n17577) );
  AO221X1 U34734 ( .IN1(n13323), .IN2(n13320), .IN3(n13318), .IN4(
        s6_msel_pri_out_1_), .IN5(n13319), .Q(n17547) );
  AO221X1 U34735 ( .IN1(n11157), .IN2(n11154), .IN3(n11152), .IN4(test_so96), 
        .IN5(n11153), .Q(n17337) );
  AO221X1 U34736 ( .IN1(n13014), .IN2(n13011), .IN3(n13009), .IN4(
        s5_msel_pri_out_1_), .IN5(n13010), .Q(n17517) );
  AO221X1 U34737 ( .IN1(n12705), .IN2(n12702), .IN3(n12700), .IN4(
        s4_msel_pri_out_1_), .IN5(n12701), .Q(n17487) );
  AO221X1 U34738 ( .IN1(n10848), .IN2(n10845), .IN3(n10843), .IN4(
        s13_msel_pri_out_1_), .IN5(n10844), .Q(n17307) );
  AO221X1 U34739 ( .IN1(n10538), .IN2(n10535), .IN3(n10533), .IN4(
        s12_msel_pri_out_1_), .IN5(n10534), .Q(n17277) );
  AO221X1 U34740 ( .IN1(n12396), .IN2(n12393), .IN3(n12391), .IN4(
        s3_msel_pri_out_1_), .IN5(n12392), .Q(n17457) );
  AO221X1 U34741 ( .IN1(n12087), .IN2(n12084), .IN3(n12082), .IN4(test_so50), 
        .IN5(n12083), .Q(n17427) );
  AO221X1 U34742 ( .IN1(n10229), .IN2(n10226), .IN3(n10224), .IN4(
        s11_msel_pri_out_1_), .IN5(n10225), .Q(n17247) );
  AO221X1 U34743 ( .IN1(n9919), .IN2(n9916), .IN3(n9914), .IN4(
        s10_msel_pri_out_1_), .IN5(n9915), .Q(n17217) );
  AO221X1 U34744 ( .IN1(n11777), .IN2(n11774), .IN3(n11772), .IN4(
        s1_msel_pri_out_1_), .IN5(n11773), .Q(n17397) );
  AO221X1 U34745 ( .IN1(n11467), .IN2(n11464), .IN3(n11462), .IN4(
        s0_msel_pri_out_1_), .IN5(n11463), .Q(n17367) );
  AO221X1 U34746 ( .IN1(n9609), .IN2(n9606), .IN3(n9604), .IN4(
        s9_msel_pri_out_1_), .IN5(n9605), .Q(n17187) );
  AO221X1 U34747 ( .IN1(n9298), .IN2(n9295), .IN3(n9293), .IN4(test_so73), 
        .IN5(n9294), .Q(n17157) );
  AO221X1 U34748 ( .IN1(n13626), .IN2(n2969), .IN3(n13627), .IN4(test_so69), 
        .IN5(n13628), .Q(n17576) );
  INVX0 U34749 ( .IN(n13629), .QN(n2969) );
  OA21X1 U34750 ( .IN1(n13630), .IN2(n13631), .IN3(n13632), .Q(n13626) );
  NAND4X0 U34751 ( .IN1(n2974), .IN2(n3144), .IN3(n3322), .IN4(n3223), .QN(
        n13631) );
  AO221X1 U34752 ( .IN1(n13317), .IN2(n2985), .IN3(n13318), .IN4(
        s6_msel_pri_out_0_), .IN5(n13319), .Q(n17546) );
  INVX0 U34753 ( .IN(n13320), .QN(n2985) );
  OA21X1 U34754 ( .IN1(n13321), .IN2(n13322), .IN3(n13323), .Q(n13317) );
  NAND4X0 U34755 ( .IN1(n2990), .IN2(n3150), .IN3(n3330), .IN4(n3227), .QN(
        n13322) );
  AO221X1 U34756 ( .IN1(n11151), .IN2(n2857), .IN3(n11152), .IN4(
        s14_msel_pri_out_0_), .IN5(n11153), .Q(n17336) );
  INVX0 U34757 ( .IN(n11154), .QN(n2857) );
  OA21X1 U34758 ( .IN1(n11155), .IN2(n11156), .IN3(n11157), .Q(n11151) );
  NAND4X0 U34759 ( .IN1(n2862), .IN2(n3102), .IN3(n3266), .IN4(n3195), .QN(
        n11156) );
  AO221X1 U34760 ( .IN1(n13008), .IN2(n3001), .IN3(n13009), .IN4(
        s5_msel_pri_out_0_), .IN5(n13010), .Q(n17516) );
  INVX0 U34761 ( .IN(n13011), .QN(n3001) );
  OA21X1 U34762 ( .IN1(n13012), .IN2(n13013), .IN3(n13014), .Q(n13008) );
  NAND4X0 U34763 ( .IN1(n3006), .IN2(n3156), .IN3(n3338), .IN4(n3231), .QN(
        n13013) );
  AO221X1 U34764 ( .IN1(n12699), .IN2(n3017), .IN3(n12700), .IN4(
        s4_msel_pri_out_0_), .IN5(n12701), .Q(n17486) );
  INVX0 U34765 ( .IN(n12702), .QN(n3017) );
  OA21X1 U34766 ( .IN1(n12703), .IN2(n12704), .IN3(n12705), .Q(n12699) );
  NAND4X0 U34767 ( .IN1(n3022), .IN2(n3162), .IN3(n3346), .IN4(n3235), .QN(
        n12704) );
  AO221X1 U34768 ( .IN1(n10842), .IN2(n2873), .IN3(n10843), .IN4(test_so92), 
        .IN5(n10844), .Q(n17306) );
  INVX0 U34769 ( .IN(n10845), .QN(n2873) );
  OA21X1 U34770 ( .IN1(n10846), .IN2(n10847), .IN3(n10848), .Q(n10842) );
  NAND4X0 U34771 ( .IN1(n2878), .IN2(n3108), .IN3(n3274), .IN4(n3199), .QN(
        n10847) );
  AO221X1 U34772 ( .IN1(n10532), .IN2(n2889), .IN3(n10533), .IN4(
        s12_msel_pri_out_0_), .IN5(n10534), .Q(n17276) );
  INVX0 U34773 ( .IN(n10535), .QN(n2889) );
  OA21X1 U34774 ( .IN1(n10536), .IN2(n10537), .IN3(n10538), .Q(n10532) );
  NAND4X0 U34775 ( .IN1(n2894), .IN2(n3114), .IN3(n3282), .IN4(n3203), .QN(
        n10537) );
  AO221X1 U34776 ( .IN1(n12390), .IN2(n3033), .IN3(n12391), .IN4(
        s3_msel_pri_out_0_), .IN5(n12392), .Q(n17456) );
  INVX0 U34777 ( .IN(n12393), .QN(n3033) );
  OA21X1 U34778 ( .IN1(n12394), .IN2(n12395), .IN3(n12396), .Q(n12390) );
  NAND4X0 U34779 ( .IN1(n3038), .IN2(n3168), .IN3(n3354), .IN4(n3239), .QN(
        n12395) );
  AO221X1 U34780 ( .IN1(n12081), .IN2(n3049), .IN3(n12082), .IN4(
        s2_msel_pri_out_0_), .IN5(n12083), .Q(n17426) );
  INVX0 U34781 ( .IN(n12084), .QN(n3049) );
  OA21X1 U34782 ( .IN1(n12085), .IN2(n12086), .IN3(n12087), .Q(n12081) );
  NAND4X0 U34783 ( .IN1(n3054), .IN2(n3174), .IN3(n3362), .IN4(n3243), .QN(
        n12086) );
  AO221X1 U34784 ( .IN1(n10223), .IN2(n2905), .IN3(n10224), .IN4(
        s11_msel_pri_out_0_), .IN5(n10225), .Q(n17246) );
  INVX0 U34785 ( .IN(n10226), .QN(n2905) );
  OA21X1 U34786 ( .IN1(n10227), .IN2(n10228), .IN3(n10229), .Q(n10223) );
  NAND4X0 U34787 ( .IN1(n2910), .IN2(n3120), .IN3(n3290), .IN4(n3207), .QN(
        n10228) );
  AO221X1 U34788 ( .IN1(n9913), .IN2(n2921), .IN3(n9914), .IN4(
        s10_msel_pri_out_0_), .IN5(n9915), .Q(n17216) );
  INVX0 U34789 ( .IN(n9916), .QN(n2921) );
  OA21X1 U34790 ( .IN1(n9917), .IN2(n9918), .IN3(n9919), .Q(n9913) );
  NAND4X0 U34791 ( .IN1(n2926), .IN2(n3126), .IN3(n3298), .IN4(n3211), .QN(
        n9918) );
  AO221X1 U34792 ( .IN1(n11771), .IN2(n3065), .IN3(n11772), .IN4(test_so46), 
        .IN5(n11773), .Q(n17396) );
  INVX0 U34793 ( .IN(n11774), .QN(n3065) );
  OA21X1 U34794 ( .IN1(n11775), .IN2(n11776), .IN3(n11777), .Q(n11771) );
  NAND4X0 U34795 ( .IN1(n3070), .IN2(n3180), .IN3(n3370), .IN4(n3247), .QN(
        n11776) );
  AO221X1 U34796 ( .IN1(n11461), .IN2(n3081), .IN3(n11462), .IN4(
        s0_msel_pri_out_0_), .IN5(n11463), .Q(n17366) );
  INVX0 U34797 ( .IN(n11464), .QN(n3081) );
  OA21X1 U34798 ( .IN1(n11465), .IN2(n11466), .IN3(n11467), .Q(n11461) );
  NAND4X0 U34799 ( .IN1(n3086), .IN2(n3186), .IN3(n3378), .IN4(n3251), .QN(
        n11466) );
  AO221X1 U34800 ( .IN1(n9603), .IN2(n2937), .IN3(n9604), .IN4(
        s9_msel_pri_out_0_), .IN5(n9605), .Q(n17186) );
  INVX0 U34801 ( .IN(n9606), .QN(n2937) );
  OA21X1 U34802 ( .IN1(n9607), .IN2(n9608), .IN3(n9609), .Q(n9603) );
  NAND4X0 U34803 ( .IN1(n2942), .IN2(n3132), .IN3(n3306), .IN4(n3215), .QN(
        n9608) );
  AO221X1 U34804 ( .IN1(n9292), .IN2(n2953), .IN3(n9293), .IN4(
        s8_msel_pri_out_0_), .IN5(n9294), .Q(n17156) );
  INVX0 U34805 ( .IN(n9295), .QN(n2953) );
  OA21X1 U34806 ( .IN1(n9296), .IN2(n9297), .IN3(n9298), .Q(n9292) );
  NAND4X0 U34807 ( .IN1(n2958), .IN2(n3138), .IN3(n3314), .IN4(n3219), .QN(
        n9297) );
  AND3X1 U34808 ( .IN1(s15_we_o), .IN2(n4502), .IN3(n18820), .Q(rf_N18) );
  OA21X1 U34809 ( .IN1(n13635), .IN2(n13636), .IN3(n13632), .Q(n13628) );
  NAND4X0 U34810 ( .IN1(n13637), .IN2(n13638), .IN3(n13639), .IN4(n13640), 
        .QN(n13636) );
  NAND4X0 U34811 ( .IN1(n13653), .IN2(n13654), .IN3(n13655), .IN4(n13656), 
        .QN(n13635) );
  NAND4X0 U34812 ( .IN1(m0s7_cyc), .IN2(n13650), .IN3(n13651), .IN4(n13652), 
        .QN(n13637) );
  OA21X1 U34813 ( .IN1(n13326), .IN2(n13327), .IN3(n13323), .Q(n13319) );
  NAND4X0 U34814 ( .IN1(n13328), .IN2(n13329), .IN3(n13330), .IN4(n13331), 
        .QN(n13327) );
  NAND4X0 U34815 ( .IN1(n13344), .IN2(n13345), .IN3(n13346), .IN4(n13347), 
        .QN(n13326) );
  NAND4X0 U34816 ( .IN1(test_so17), .IN2(n13341), .IN3(n13342), .IN4(n13343), 
        .QN(n13328) );
  OA21X1 U34817 ( .IN1(n11160), .IN2(n11161), .IN3(n11157), .Q(n11153) );
  NAND4X0 U34818 ( .IN1(n11162), .IN2(n11163), .IN3(n11164), .IN4(n11165), 
        .QN(n11161) );
  NAND4X0 U34819 ( .IN1(n11178), .IN2(n11179), .IN3(n11180), .IN4(n11181), 
        .QN(n11160) );
  NAND4X0 U34820 ( .IN1(m0s14_cyc), .IN2(n11175), .IN3(n11176), .IN4(n11177), 
        .QN(n11162) );
  OA21X1 U34821 ( .IN1(n13017), .IN2(n13018), .IN3(n13014), .Q(n13010) );
  NAND4X0 U34822 ( .IN1(n13019), .IN2(n13020), .IN3(n13021), .IN4(n13022), 
        .QN(n13018) );
  NAND4X0 U34823 ( .IN1(n13035), .IN2(n13036), .IN3(n13037), .IN4(n13038), 
        .QN(n13017) );
  NAND4X0 U34824 ( .IN1(m0s5_cyc), .IN2(n13032), .IN3(n13033), .IN4(n13034), 
        .QN(n13019) );
  OA21X1 U34825 ( .IN1(n12708), .IN2(n12709), .IN3(n12705), .Q(n12701) );
  NAND4X0 U34826 ( .IN1(n12710), .IN2(n12711), .IN3(n12712), .IN4(n12713), 
        .QN(n12709) );
  NAND4X0 U34827 ( .IN1(n12726), .IN2(n12727), .IN3(n12728), .IN4(n12729), 
        .QN(n12708) );
  NAND4X0 U34828 ( .IN1(m0s4_cyc), .IN2(n12723), .IN3(n12724), .IN4(n12725), 
        .QN(n12710) );
  OA21X1 U34829 ( .IN1(n10851), .IN2(n10852), .IN3(n10848), .Q(n10844) );
  NAND4X0 U34830 ( .IN1(n10853), .IN2(n10854), .IN3(n10855), .IN4(n10856), 
        .QN(n10852) );
  NAND4X0 U34831 ( .IN1(n10869), .IN2(n10870), .IN3(n10871), .IN4(n10872), 
        .QN(n10851) );
  NAND4X0 U34832 ( .IN1(test_so18), .IN2(n10866), .IN3(n10867), .IN4(n10868), 
        .QN(n10853) );
  OA21X1 U34833 ( .IN1(n10541), .IN2(n10542), .IN3(n10538), .Q(n10534) );
  NAND4X0 U34834 ( .IN1(n10543), .IN2(n10544), .IN3(n10545), .IN4(n10546), 
        .QN(n10542) );
  NAND4X0 U34835 ( .IN1(n10559), .IN2(n10560), .IN3(n10561), .IN4(n10562), 
        .QN(n10541) );
  NAND4X0 U34836 ( .IN1(m0s12_cyc), .IN2(n10556), .IN3(n10557), .IN4(n10558), 
        .QN(n10543) );
  OA21X1 U34837 ( .IN1(n12399), .IN2(n12400), .IN3(n12396), .Q(n12392) );
  NAND4X0 U34838 ( .IN1(n12401), .IN2(n12402), .IN3(n12403), .IN4(n12404), 
        .QN(n12400) );
  NAND4X0 U34839 ( .IN1(n12417), .IN2(n12418), .IN3(n12419), .IN4(n12420), 
        .QN(n12399) );
  NAND4X0 U34840 ( .IN1(m0s3_cyc), .IN2(n12414), .IN3(n12415), .IN4(n12416), 
        .QN(n12401) );
  OA21X1 U34841 ( .IN1(n12090), .IN2(n12091), .IN3(n12087), .Q(n12083) );
  NAND4X0 U34842 ( .IN1(n12092), .IN2(n12093), .IN3(n12094), .IN4(n12095), 
        .QN(n12091) );
  NAND4X0 U34843 ( .IN1(n12108), .IN2(n12109), .IN3(n12110), .IN4(n12111), 
        .QN(n12090) );
  NAND4X0 U34844 ( .IN1(m0s2_cyc), .IN2(n12105), .IN3(n12106), .IN4(n12107), 
        .QN(n12092) );
  OA21X1 U34845 ( .IN1(n10232), .IN2(n10233), .IN3(n10229), .Q(n10225) );
  NAND4X0 U34846 ( .IN1(n10234), .IN2(n10235), .IN3(n10236), .IN4(n10237), 
        .QN(n10233) );
  NAND4X0 U34847 ( .IN1(n10250), .IN2(n10251), .IN3(n10252), .IN4(n10253), 
        .QN(n10232) );
  NAND4X0 U34848 ( .IN1(m0s11_cyc), .IN2(n10247), .IN3(n10248), .IN4(n10249), 
        .QN(n10234) );
  OA21X1 U34849 ( .IN1(n9922), .IN2(n9923), .IN3(n9919), .Q(n9915) );
  NAND4X0 U34850 ( .IN1(n9924), .IN2(n9925), .IN3(n9926), .IN4(n9927), .QN(
        n9923) );
  NAND4X0 U34851 ( .IN1(n9940), .IN2(n9941), .IN3(n9942), .IN4(n9943), .QN(
        n9922) );
  NAND4X0 U34852 ( .IN1(m0s10_cyc), .IN2(n9937), .IN3(n9938), .IN4(n9939), 
        .QN(n9924) );
  OA21X1 U34853 ( .IN1(n11780), .IN2(n11781), .IN3(n11777), .Q(n11773) );
  NAND4X0 U34854 ( .IN1(n11782), .IN2(n11783), .IN3(n11784), .IN4(n11785), 
        .QN(n11781) );
  NAND4X0 U34855 ( .IN1(n11798), .IN2(n11799), .IN3(n11800), .IN4(n11801), 
        .QN(n11780) );
  NAND4X0 U34856 ( .IN1(m0s1_cyc), .IN2(n11795), .IN3(n11796), .IN4(n11797), 
        .QN(n11782) );
  OA21X1 U34857 ( .IN1(n11470), .IN2(n11471), .IN3(n11467), .Q(n11463) );
  NAND4X0 U34858 ( .IN1(n11472), .IN2(n11473), .IN3(n11474), .IN4(n11475), 
        .QN(n11471) );
  NAND4X0 U34859 ( .IN1(n11488), .IN2(n11489), .IN3(n11490), .IN4(n11491), 
        .QN(n11470) );
  NAND4X0 U34860 ( .IN1(m0s0_cyc), .IN2(n11485), .IN3(n11486), .IN4(n11487), 
        .QN(n11472) );
  OA21X1 U34861 ( .IN1(n9612), .IN2(n9613), .IN3(n9609), .Q(n9605) );
  NAND4X0 U34862 ( .IN1(n9614), .IN2(n9615), .IN3(n9616), .IN4(n9617), .QN(
        n9613) );
  NAND4X0 U34863 ( .IN1(n9630), .IN2(n9631), .IN3(n9632), .IN4(n9633), .QN(
        n9612) );
  NAND4X0 U34864 ( .IN1(m0s9_cyc), .IN2(n9627), .IN3(n9628), .IN4(n9629), .QN(
        n9614) );
  OA21X1 U34865 ( .IN1(n9301), .IN2(n9302), .IN3(n9298), .Q(n9294) );
  NAND4X0 U34866 ( .IN1(n9303), .IN2(n9304), .IN3(n9305), .IN4(n9306), .QN(
        n9302) );
  NAND4X0 U34867 ( .IN1(n9319), .IN2(n9320), .IN3(n9321), .IN4(n9322), .QN(
        n9301) );
  NAND4X0 U34868 ( .IN1(m0s8_cyc), .IN2(n9316), .IN3(n9317), .IN4(n9318), .QN(
        n9303) );
  NOR2X0 U34869 ( .IN1(n14410), .IN2(n14411), .QN(n17772) );
  NAND4X0 U34870 ( .IN1(n14412), .IN2(n14413), .IN3(n14414), .IN4(n14415), 
        .QN(n14411) );
  NAND4X0 U34871 ( .IN1(n14416), .IN2(n14417), .IN3(n14418), .IN4(n14419), 
        .QN(n14410) );
  NAND3X0 U34872 ( .IN1(m1s7_cyc), .IN2(n20567), .IN3(s7_m1_cyc_r), .QN(n14413) );
  NOR2X0 U34873 ( .IN1(n14420), .IN2(n14421), .QN(n17773) );
  NAND4X0 U34874 ( .IN1(n14422), .IN2(n14423), .IN3(n14424), .IN4(n14425), 
        .QN(n14421) );
  NAND4X0 U34875 ( .IN1(n14426), .IN2(n14427), .IN3(n14428), .IN4(n14429), 
        .QN(n14420) );
  NAND3X0 U34876 ( .IN1(m1s6_cyc), .IN2(n20435), .IN3(test_so62), .QN(n14423)
         );
  NOR2X0 U34877 ( .IN1(n14340), .IN2(n14341), .QN(n17765) );
  NAND4X0 U34878 ( .IN1(n14342), .IN2(n14343), .IN3(n14344), .IN4(n14345), 
        .QN(n14341) );
  NAND4X0 U34879 ( .IN1(n14346), .IN2(n14347), .IN3(n14348), .IN4(n14349), 
        .QN(n14340) );
  NAND3X0 U34880 ( .IN1(m1s14_cyc), .IN2(n19513), .IN3(s14_m1_cyc_r), .QN(
        n14343) );
  NAND4X0 U34881 ( .IN1(n14432), .IN2(n14433), .IN3(n14434), .IN4(n14435), 
        .QN(n14431) );
  NAND4X0 U34882 ( .IN1(n14436), .IN2(n14437), .IN3(n14438), .IN4(n14439), 
        .QN(n14430) );
  NAND3X0 U34883 ( .IN1(m1s5_cyc), .IN2(n20303), .IN3(s5_m1_cyc_r), .QN(n14433) );
  NAND4X0 U34884 ( .IN1(n14442), .IN2(n14443), .IN3(n14444), .IN4(n14445), 
        .QN(n14441) );
  NAND4X0 U34885 ( .IN1(n14446), .IN2(n14447), .IN3(n14448), .IN4(n14449), 
        .QN(n14440) );
  NAND3X0 U34886 ( .IN1(test_so19), .IN2(n20171), .IN3(s4_m1_cyc_r), .QN(
        n14443) );
  NAND4X0 U34887 ( .IN1(n14352), .IN2(n14353), .IN3(n14354), .IN4(n14355), 
        .QN(n14351) );
  NAND4X0 U34888 ( .IN1(n14356), .IN2(n14357), .IN3(n14358), .IN4(n14359), 
        .QN(n14350) );
  NAND3X0 U34889 ( .IN1(m1s13_cyc), .IN2(n19381), .IN3(s13_m1_cyc_r), .QN(
        n14353) );
  NAND4X0 U34890 ( .IN1(n14362), .IN2(n14363), .IN3(n14364), .IN4(n14365), 
        .QN(n14361) );
  NAND4X0 U34891 ( .IN1(n14366), .IN2(n14367), .IN3(n14368), .IN4(n14369), 
        .QN(n14360) );
  NAND3X0 U34892 ( .IN1(m1s12_cyc), .IN2(n19249), .IN3(test_so85), .QN(n14363)
         );
  NOR2X0 U34893 ( .IN1(n14450), .IN2(n14451), .QN(n17776) );
  NAND4X0 U34894 ( .IN1(n14452), .IN2(n14453), .IN3(n14454), .IN4(n14455), 
        .QN(n14451) );
  NAND4X0 U34895 ( .IN1(n14456), .IN2(n14457), .IN3(n14458), .IN4(n14459), 
        .QN(n14450) );
  NAND3X0 U34896 ( .IN1(m1s3_cyc), .IN2(n20040), .IN3(s3_m1_cyc_r), .QN(n14453) );
  NOR2X0 U34897 ( .IN1(n14460), .IN2(n14461), .QN(n17777) );
  NAND4X0 U34898 ( .IN1(n14462), .IN2(n14463), .IN3(n14464), .IN4(n14465), 
        .QN(n14461) );
  NAND4X0 U34899 ( .IN1(n14466), .IN2(n14467), .IN3(n14468), .IN4(n14469), 
        .QN(n14460) );
  NAND3X0 U34900 ( .IN1(m1s2_cyc), .IN2(n19909), .IN3(s2_m1_cyc_r), .QN(n14463) );
  NAND4X0 U34901 ( .IN1(n14372), .IN2(n14373), .IN3(n14374), .IN4(n14375), 
        .QN(n14371) );
  NAND4X0 U34902 ( .IN1(n14376), .IN2(n14377), .IN3(n14378), .IN4(n14379), 
        .QN(n14370) );
  NAND3X0 U34903 ( .IN1(test_so20), .IN2(n19117), .IN3(s11_m1_cyc_r), .QN(
        n14373) );
  NAND4X0 U34904 ( .IN1(n14382), .IN2(n14383), .IN3(n14384), .IN4(n14385), 
        .QN(n14381) );
  NAND4X0 U34905 ( .IN1(n14386), .IN2(n14387), .IN3(n14388), .IN4(n14389), 
        .QN(n14380) );
  NAND3X0 U34906 ( .IN1(m1s10_cyc), .IN2(n18985), .IN3(s10_m1_cyc_r), .QN(
        n14383) );
  NAND4X0 U34907 ( .IN1(n14472), .IN2(n14473), .IN3(n14474), .IN4(n14475), 
        .QN(n14471) );
  NAND4X0 U34908 ( .IN1(n14476), .IN2(n14477), .IN3(n14478), .IN4(n14479), 
        .QN(n14470) );
  NAND3X0 U34909 ( .IN1(m1s1_cyc), .IN2(n19777), .IN3(s1_m1_cyc_r), .QN(n14473) );
  NAND4X0 U34910 ( .IN1(n14482), .IN2(n14483), .IN3(n14484), .IN4(n14485), 
        .QN(n14481) );
  NAND4X0 U34911 ( .IN1(n14486), .IN2(n14487), .IN3(n14488), .IN4(n14489), 
        .QN(n14480) );
  NAND3X0 U34912 ( .IN1(m1s0_cyc), .IN2(n18853), .IN3(test_so39), .QN(n14483)
         );
  NOR2X0 U34913 ( .IN1(n14390), .IN2(n14391), .QN(n17770) );
  NAND4X0 U34914 ( .IN1(n14392), .IN2(n14393), .IN3(n14394), .IN4(n14395), 
        .QN(n14391) );
  NAND4X0 U34915 ( .IN1(n14396), .IN2(n14397), .IN3(n14398), .IN4(n14399), 
        .QN(n14390) );
  NAND3X0 U34916 ( .IN1(m0s9_cyc), .IN2(n20807), .IN3(s9_m0_cyc_r), .QN(n14392) );
  NAND4X0 U34917 ( .IN1(n14402), .IN2(n14403), .IN3(n14404), .IN4(n14405), 
        .QN(n14401) );
  NAND4X0 U34918 ( .IN1(n14406), .IN2(n14407), .IN3(n14408), .IN4(n14409), 
        .QN(n14400) );
  NAND3X0 U34919 ( .IN1(m1s8_cyc), .IN2(n20699), .IN3(s8_m1_cyc_r), .QN(n14403) );
  AO221X1 U34920 ( .IN1(n14275), .IN2(n14272), .IN3(n14270), .IN4(
        s15_msel_pri_out_1_), .IN5(n14271), .Q(n17634) );
  AO221X1 U34921 ( .IN1(n14269), .IN2(n2847), .IN3(n14270), .IN4(
        s15_msel_pri_out_0_), .IN5(n14271), .Q(n17633) );
  INVX0 U34922 ( .IN(n14272), .QN(n2847) );
  OA21X1 U34923 ( .IN1(n14273), .IN2(n14274), .IN3(n14275), .Q(n14269) );
  NAND4X0 U34924 ( .IN1(n3191), .IN2(n3095), .IN3(n13944), .IN4(n3258), .QN(
        n14274) );
  NAND3X0 U34925 ( .IN1(n18333), .IN2(n20621), .IN3(s7_m4_cyc_r), .QN(n14416)
         );
  NAND3X0 U34926 ( .IN1(n18332), .IN2(n20489), .IN3(s6_m4_cyc_r), .QN(n14426)
         );
  NAND3X0 U34927 ( .IN1(n18331), .IN2(n19567), .IN3(s14_m4_cyc_r), .QN(n14346)
         );
  NAND3X0 U34928 ( .IN1(n18330), .IN2(n20360), .IN3(s5_m4_cyc_r), .QN(n14436)
         );
  NAND3X0 U34929 ( .IN1(n18329), .IN2(n20228), .IN3(s4_m4_cyc_r), .QN(n14446)
         );
  NAND3X0 U34930 ( .IN1(n18328), .IN2(n19438), .IN3(s13_m4_cyc_r), .QN(n14356)
         );
  NAND3X0 U34931 ( .IN1(n18327), .IN2(n19306), .IN3(s12_m4_cyc_r), .QN(n14366)
         );
  NAND3X0 U34932 ( .IN1(n18326), .IN2(n20096), .IN3(test_so51), .QN(n14456) );
  NAND3X0 U34933 ( .IN1(n18325), .IN2(n19962), .IN3(s2_m4_cyc_r), .QN(n14466)
         );
  NAND3X0 U34934 ( .IN1(n18324), .IN2(n19174), .IN3(s11_m4_cyc_r), .QN(n14376)
         );
  NAND3X0 U34935 ( .IN1(n18323), .IN2(n19042), .IN3(s10_m4_cyc_r), .QN(n14386)
         );
  NAND3X0 U34936 ( .IN1(n18322), .IN2(n19834), .IN3(s1_m4_cyc_r), .QN(n14476)
         );
  NAND3X0 U34937 ( .IN1(n18321), .IN2(n18910), .IN3(s0_m4_cyc_r), .QN(n14486)
         );
  NAND3X0 U34938 ( .IN1(n18320), .IN2(n20843), .IN3(test_so74), .QN(n14396) );
  NAND3X0 U34939 ( .IN1(n18319), .IN2(n20756), .IN3(s8_m4_cyc_r), .QN(n14406)
         );
  NOR2X0 U34940 ( .IN1(rf_rf_ack), .IN2(n18816), .QN(rf_N19) );
  AO22X1 U34941 ( .IN1(n14328), .IN2(m5s15_cyc), .IN3(n14329), .IN4(n17782), 
        .Q(n17683) );
  AO22X1 U34942 ( .IN1(n14328), .IN2(test_so28), .IN3(n14329), .IN4(n17829), 
        .Q(n17669) );
  AO22X1 U34943 ( .IN1(n14328), .IN2(m5s3_cyc), .IN3(n14329), .IN4(n17797), 
        .Q(n17671) );
  AO22X1 U34944 ( .IN1(n14328), .IN2(m5s5_cyc), .IN3(n14329), .IN4(n17799), 
        .Q(n17673) );
  AO22X1 U34945 ( .IN1(n14328), .IN2(m5s9_cyc), .IN3(n14329), .IN4(n17874), 
        .Q(n17677) );
  AO22X1 U34946 ( .IN1(n14328), .IN2(m5s11_cyc), .IN3(n14329), .IN4(n17821), 
        .Q(n17679) );
  AO22X1 U34947 ( .IN1(n14328), .IN2(test_so30), .IN3(n14329), .IN4(n17812), 
        .Q(n17681) );
  AO22X1 U34948 ( .IN1(n14328), .IN2(m5s6_cyc), .IN3(n14329), .IN4(n17872), 
        .Q(n17674) );
  NAND4X0 U34949 ( .IN1(m5s6_cyc), .IN2(n13354), .IN3(n13355), .IN4(n13356), 
        .QN(n13345) );
  NAND4X0 U34950 ( .IN1(m5s5_cyc), .IN2(n13045), .IN3(n13046), .IN4(n13047), 
        .QN(n13036) );
  NAND4X0 U34951 ( .IN1(test_so30), .IN2(n10879), .IN3(n10880), .IN4(n10881), 
        .QN(n10870) );
  NAND4X0 U34952 ( .IN1(m5s3_cyc), .IN2(n12427), .IN3(n12428), .IN4(n12429), 
        .QN(n12418) );
  NAND4X0 U34953 ( .IN1(m5s11_cyc), .IN2(n10260), .IN3(n10261), .IN4(n10262), 
        .QN(n10251) );
  NAND4X0 U34954 ( .IN1(test_so28), .IN2(n11808), .IN3(n11809), .IN4(n11810), 
        .QN(n11799) );
  NAND4X0 U34955 ( .IN1(m5s9_cyc), .IN2(n9640), .IN3(n9641), .IN4(n9642), .QN(
        n9631) );
  NAND4X0 U34956 ( .IN1(m5s15_cyc), .IN2(n14300), .IN3(n14071), .IN4(n14282), 
        .QN(n14295) );
  OA21X1 U34957 ( .IN1(n14284), .IN2(n14285), .IN3(n14275), .Q(n14271) );
  NAND4X0 U34958 ( .IN1(n14286), .IN2(n14287), .IN3(n14288), .IN4(n14289), 
        .QN(n14285) );
  NAND4X0 U34959 ( .IN1(n14294), .IN2(n14295), .IN3(n14296), .IN4(n14297), 
        .QN(n14284) );
  NAND4X0 U34960 ( .IN1(m0s15_cyc), .IN2(n14293), .IN3(n14074), .IN4(n14281), 
        .QN(n14286) );
  NAND3X0 U34961 ( .IN1(m4s15_cyc), .IN2(n19702), .IN3(test_so97), .QN(n17101)
         );
  ISOLANDX1 U34962 ( .D(m4s15_cyc), .ISO(n14301), .Q(n14141) );
  AO221X1 U34963 ( .IN1(s15_msel_gnt_p3[2]), .IN2(n17120), .IN3(test_so99), 
        .IN4(n17121), .IN5(n17122), .Q(n17118) );
  AO22X1 U34964 ( .IN1(test_so98), .IN2(n17123), .IN3(s15_msel_gnt_p1[2]), 
        .IN4(n17124), .Q(n17122) );
  AO221X1 U34965 ( .IN1(s15_msel_gnt_p3[1]), .IN2(n17120), .IN3(
        s15_msel_gnt_p2_1_), .IN4(n17121), .IN5(n17126), .Q(n17117) );
  AO22X1 U34966 ( .IN1(s15_msel_gnt_p0_1_), .IN2(n17123), .IN3(
        s15_msel_gnt_p1[1]), .IN4(n17124), .Q(n17126) );
  AO221X1 U34967 ( .IN1(s15_msel_gnt_p3[0]), .IN2(n17120), .IN3(
        s15_msel_gnt_p2_0_), .IN4(n17121), .IN5(n17125), .Q(n17119) );
  AO22X1 U34968 ( .IN1(s15_msel_gnt_p0_0_), .IN2(n17123), .IN3(
        s15_msel_gnt_p1[0]), .IN4(n17124), .Q(n17125) );
  NAND3X0 U34969 ( .IN1(conf15_9_), .IN2(m4s15_cyc), .IN3(conf15_8_), .QN(
        n14187) );
  ISOLANDX1 U34970 ( .D(m2s7_cyc), .ISO(n13644), .Q(n13769) );
  ISOLANDX1 U34971 ( .D(m2s6_cyc), .ISO(n13335), .Q(n13460) );
  ISOLANDX1 U34972 ( .D(m2s14_cyc), .ISO(n11169), .Q(n11294) );
  ISOLANDX1 U34973 ( .D(m2s5_cyc), .ISO(n13026), .Q(n13151) );
  ISOLANDX1 U34974 ( .D(m2s4_cyc), .ISO(n12717), .Q(n12842) );
  ISOLANDX1 U34975 ( .D(m2s13_cyc), .ISO(n10860), .Q(n10985) );
  ISOLANDX1 U34976 ( .D(m2s12_cyc), .ISO(n10550), .Q(n10675) );
  ISOLANDX1 U34977 ( .D(m2s3_cyc), .ISO(n12408), .Q(n12533) );
  ISOLANDX1 U34978 ( .D(test_so21), .ISO(n12099), .Q(n12224) );
  ISOLANDX1 U34979 ( .D(m2s11_cyc), .ISO(n10241), .Q(n10366) );
  ISOLANDX1 U34980 ( .D(m2s10_cyc), .ISO(n9931), .Q(n10056) );
  ISOLANDX1 U34981 ( .D(m2s1_cyc), .ISO(n11789), .Q(n11914) );
  ISOLANDX1 U34982 ( .D(m2s0_cyc), .ISO(n11479), .Q(n11604) );
  ISOLANDX1 U34983 ( .D(test_so22), .ISO(n9621), .Q(n9746) );
  ISOLANDX1 U34984 ( .D(m2s8_cyc), .ISO(n9310), .Q(n9435) );
  ISOLANDX1 U34985 ( .D(m2s15_cyc), .ISO(n14072), .Q(n14033) );
  ISOLANDX1 U34986 ( .D(m1s7_cyc), .ISO(n13647), .Q(n13772) );
  ISOLANDX1 U34987 ( .D(m1s6_cyc), .ISO(n13338), .Q(n13463) );
  ISOLANDX1 U34988 ( .D(m1s14_cyc), .ISO(n11172), .Q(n11297) );
  ISOLANDX1 U34989 ( .D(m1s5_cyc), .ISO(n13029), .Q(n13154) );
  ISOLANDX1 U34990 ( .D(test_so19), .ISO(n12720), .Q(n12845) );
  ISOLANDX1 U34991 ( .D(m1s13_cyc), .ISO(n10863), .Q(n10988) );
  ISOLANDX1 U34992 ( .D(m1s12_cyc), .ISO(n10553), .Q(n10678) );
  ISOLANDX1 U34993 ( .D(m1s3_cyc), .ISO(n12411), .Q(n12536) );
  ISOLANDX1 U34994 ( .D(m1s2_cyc), .ISO(n12102), .Q(n12227) );
  ISOLANDX1 U34995 ( .D(test_so20), .ISO(n10244), .Q(n10369) );
  ISOLANDX1 U34996 ( .D(m1s10_cyc), .ISO(n9934), .Q(n10059) );
  ISOLANDX1 U34997 ( .D(m1s1_cyc), .ISO(n11792), .Q(n11917) );
  ISOLANDX1 U34998 ( .D(m1s0_cyc), .ISO(n11482), .Q(n11607) );
  ISOLANDX1 U34999 ( .D(m1s9_cyc), .ISO(n9624), .Q(n9749) );
  ISOLANDX1 U35000 ( .D(m1s8_cyc), .ISO(n9313), .Q(n9438) );
  ISOLANDX1 U35001 ( .D(m1s15_cyc), .ISO(n14075), .Q(n14036) );
  ISOLANDX1 U35002 ( .D(m0s7_cyc), .ISO(n13650), .Q(n13786) );
  ISOLANDX1 U35003 ( .D(test_so17), .ISO(n13341), .Q(n13477) );
  ISOLANDX1 U35004 ( .D(m0s14_cyc), .ISO(n11175), .Q(n11311) );
  ISOLANDX1 U35005 ( .D(m0s5_cyc), .ISO(n13032), .Q(n13168) );
  ISOLANDX1 U35006 ( .D(m0s4_cyc), .ISO(n12723), .Q(n12859) );
  ISOLANDX1 U35007 ( .D(test_so18), .ISO(n10866), .Q(n11002) );
  ISOLANDX1 U35008 ( .D(m0s12_cyc), .ISO(n10556), .Q(n10692) );
  ISOLANDX1 U35009 ( .D(m0s3_cyc), .ISO(n12414), .Q(n12550) );
  ISOLANDX1 U35010 ( .D(m0s2_cyc), .ISO(n12105), .Q(n12241) );
  ISOLANDX1 U35011 ( .D(m0s11_cyc), .ISO(n10247), .Q(n10383) );
  ISOLANDX1 U35012 ( .D(m0s10_cyc), .ISO(n9937), .Q(n10073) );
  ISOLANDX1 U35013 ( .D(m0s1_cyc), .ISO(n11795), .Q(n11931) );
  ISOLANDX1 U35014 ( .D(m0s0_cyc), .ISO(n11485), .Q(n11621) );
  ISOLANDX1 U35015 ( .D(m0s9_cyc), .ISO(n9627), .Q(n9763) );
  ISOLANDX1 U35016 ( .D(m0s8_cyc), .ISO(n9316), .Q(n9452) );
  ISOLANDX1 U35017 ( .D(m0s15_cyc), .ISO(n14074), .Q(n14050) );
  NOR2X0 U35018 ( .IN1(n4213), .IN2(s15_msel_pri_out_0_), .QN(n17121) );
  NOR2X0 U35019 ( .IN1(n4213), .IN2(n4212), .QN(n17120) );
  NOR2X0 U35020 ( .IN1(s15_msel_pri_out_0_), .IN2(s15_msel_pri_out_1_), .QN(
        n17123) );
  NOR2X0 U35021 ( .IN1(n4212), .IN2(s15_msel_pri_out_1_), .QN(n17124) );
  NAND3X0 U35022 ( .IN1(n3860), .IN2(n3861), .IN3(n3859), .QN(n13773) );
  NAND3X0 U35023 ( .IN1(n3815), .IN2(n3816), .IN3(n3814), .QN(n13464) );
  NAND3X0 U35024 ( .IN1(n4175), .IN2(n4176), .IN3(n4174), .QN(n11298) );
  NAND3X0 U35025 ( .IN1(n3770), .IN2(n3771), .IN3(n3769), .QN(n13155) );
  NAND3X0 U35026 ( .IN1(n3725), .IN2(n3726), .IN3(n3724), .QN(n12846) );
  NAND3X0 U35027 ( .IN1(n4130), .IN2(n4131), .IN3(n4129), .QN(n10989) );
  NAND3X0 U35028 ( .IN1(n4085), .IN2(n4086), .IN3(n4084), .QN(n10679) );
  NAND3X0 U35029 ( .IN1(n3680), .IN2(n3681), .IN3(n3679), .QN(n12537) );
  NAND3X0 U35030 ( .IN1(n3635), .IN2(n3636), .IN3(n3634), .QN(n12228) );
  NAND3X0 U35031 ( .IN1(n4040), .IN2(n4041), .IN3(n4039), .QN(n10370) );
  NAND3X0 U35032 ( .IN1(n3995), .IN2(n3996), .IN3(n3994), .QN(n10060) );
  NAND3X0 U35033 ( .IN1(n3590), .IN2(n3591), .IN3(n3589), .QN(n11918) );
  NAND3X0 U35034 ( .IN1(n3545), .IN2(n3546), .IN3(n3544), .QN(n11608) );
  NAND3X0 U35035 ( .IN1(n3950), .IN2(n3951), .IN3(n3949), .QN(n9750) );
  NAND3X0 U35036 ( .IN1(n3905), .IN2(n3906), .IN3(n3904), .QN(n9439) );
  NAND3X0 U35037 ( .IN1(n4220), .IN2(n4221), .IN3(n4219), .QN(n14037) );
  NAND3X0 U35038 ( .IN1(n3860), .IN2(n3861), .IN3(test_so67), .QN(n13774) );
  NAND3X0 U35039 ( .IN1(n3815), .IN2(n3816), .IN3(s6_msel_gnt_p0[0]), .QN(
        n13465) );
  NAND3X0 U35040 ( .IN1(n4175), .IN2(n4176), .IN3(s14_msel_gnt_p0_0_), .QN(
        n11299) );
  NAND3X0 U35041 ( .IN1(n3770), .IN2(n3771), .IN3(s5_msel_gnt_p0[0]), .QN(
        n13156) );
  NAND3X0 U35042 ( .IN1(n3725), .IN2(n3726), .IN3(s4_msel_gnt_p0[0]), .QN(
        n12847) );
  NAND3X0 U35043 ( .IN1(n4130), .IN2(n4131), .IN3(test_so90), .QN(n10990) );
  NAND3X0 U35044 ( .IN1(n4085), .IN2(n4086), .IN3(s12_msel_gnt_p0[0]), .QN(
        n10680) );
  NAND3X0 U35045 ( .IN1(n3680), .IN2(n3681), .IN3(s3_msel_gnt_p0_0_), .QN(
        n12538) );
  NAND3X0 U35046 ( .IN1(n3635), .IN2(n3636), .IN3(s2_msel_gnt_p0_0_), .QN(
        n12229) );
  NAND3X0 U35047 ( .IN1(n4040), .IN2(n4041), .IN3(s11_msel_gnt_p0[0]), .QN(
        n10371) );
  NAND3X0 U35048 ( .IN1(n3995), .IN2(n3996), .IN3(s10_msel_gnt_p0[0]), .QN(
        n10061) );
  NAND3X0 U35049 ( .IN1(n3590), .IN2(n3591), .IN3(test_so44), .QN(n11919) );
  NAND3X0 U35050 ( .IN1(n3545), .IN2(n3546), .IN3(s0_msel_gnt_p0[0]), .QN(
        n11609) );
  NAND3X0 U35051 ( .IN1(n3950), .IN2(n3951), .IN3(s9_msel_gnt_p0_0_), .QN(
        n9751) );
  NAND3X0 U35052 ( .IN1(n3905), .IN2(n3906), .IN3(s8_msel_gnt_p0_0_), .QN(
        n9440) );
  NAND3X0 U35053 ( .IN1(n4220), .IN2(n4221), .IN3(s15_msel_gnt_p0_0_), .QN(
        n14038) );
  NAND3X0 U35054 ( .IN1(s7_msel_gnt_p0_1_), .IN2(s7_msel_gnt_p0_2_), .IN3(
        test_so67), .QN(n13799) );
  NAND3X0 U35055 ( .IN1(s6_msel_gnt_p0[1]), .IN2(s6_msel_gnt_p0[2]), .IN3(
        s6_msel_gnt_p0[0]), .QN(n13490) );
  NAND3X0 U35056 ( .IN1(test_so94), .IN2(s14_msel_gnt_p0_2_), .IN3(
        s14_msel_gnt_p0_0_), .QN(n11324) );
  NAND3X0 U35057 ( .IN1(s5_msel_gnt_p0[1]), .IN2(s5_msel_gnt_p0[2]), .IN3(
        s5_msel_gnt_p0[0]), .QN(n13181) );
  NAND3X0 U35058 ( .IN1(s4_msel_gnt_p0[1]), .IN2(s4_msel_gnt_p0[2]), .IN3(
        s4_msel_gnt_p0[0]), .QN(n12872) );
  NAND3X0 U35059 ( .IN1(s13_msel_gnt_p0_1_), .IN2(s13_msel_gnt_p0_2_), .IN3(
        test_so90), .QN(n11015) );
  NAND3X0 U35060 ( .IN1(s12_msel_gnt_p0[1]), .IN2(s12_msel_gnt_p0[2]), .IN3(
        s12_msel_gnt_p0[0]), .QN(n10705) );
  NAND3X0 U35061 ( .IN1(s3_msel_gnt_p0_1_), .IN2(test_so52), .IN3(
        s3_msel_gnt_p0_0_), .QN(n12563) );
  NAND3X0 U35062 ( .IN1(test_so48), .IN2(s2_msel_gnt_p0_2_), .IN3(
        s2_msel_gnt_p0_0_), .QN(n12254) );
  NAND3X0 U35063 ( .IN1(s11_msel_gnt_p0[1]), .IN2(s11_msel_gnt_p0[2]), .IN3(
        s11_msel_gnt_p0[0]), .QN(n10396) );
  NAND3X0 U35064 ( .IN1(s10_msel_gnt_p0[1]), .IN2(s10_msel_gnt_p0[2]), .IN3(
        s10_msel_gnt_p0[0]), .QN(n10086) );
  NAND3X0 U35065 ( .IN1(s1_msel_gnt_p0_1_), .IN2(s1_msel_gnt_p0_2_), .IN3(
        test_so44), .QN(n11944) );
  NAND3X0 U35066 ( .IN1(s0_msel_gnt_p0[1]), .IN2(s0_msel_gnt_p0[2]), .IN3(
        s0_msel_gnt_p0[0]), .QN(n11634) );
  NAND3X0 U35067 ( .IN1(s9_msel_gnt_p0_1_), .IN2(test_so75), .IN3(
        s9_msel_gnt_p0_0_), .QN(n9776) );
  NAND3X0 U35068 ( .IN1(test_so71), .IN2(s8_msel_gnt_p0_2_), .IN3(
        s8_msel_gnt_p0_0_), .QN(n9465) );
  NAND3X0 U35069 ( .IN1(s15_msel_gnt_p0_1_), .IN2(test_so98), .IN3(
        s15_msel_gnt_p0_0_), .QN(n14063) );
  NAND3X0 U35070 ( .IN1(test_so33), .IN2(n19735), .IN3(s15_m6_cyc_r), .QN(
        n17103) );
  NAND3X0 U35071 ( .IN1(m2s15_cyc), .IN2(n19669), .IN3(s15_m2_cyc_r), .QN(
        n17099) );
  NAND3X0 U35072 ( .IN1(m0s15_cyc), .IN2(n19636), .IN3(s15_m0_cyc_r), .QN(
        n17097) );
  NAND2X0 U35073 ( .IN1(conf7_9_), .IN2(n18152), .QN(n13668) );
  NAND2X0 U35074 ( .IN1(conf5_9_), .IN2(n17935), .QN(n13050) );
  NAND2X0 U35075 ( .IN1(conf4_9_), .IN2(n18066), .QN(n12741) );
  NAND2X0 U35076 ( .IN1(conf13_9_), .IN2(n17936), .QN(n10884) );
  NAND2X0 U35077 ( .IN1(conf12_9_), .IN2(n18083), .QN(n10574) );
  NAND2X0 U35078 ( .IN1(conf3_9_), .IN2(n18151), .QN(n12432) );
  NAND2X0 U35079 ( .IN1(conf11_9_), .IN2(n17937), .QN(n10265) );
  NAND2X0 U35080 ( .IN1(conf10_9_), .IN2(n18084), .QN(n9955) );
  NAND2X0 U35081 ( .IN1(conf1_9_), .IN2(n17938), .QN(n11813) );
  NAND2X0 U35082 ( .IN1(conf0_9_), .IN2(n18085), .QN(n11503) );
  NAND2X0 U35083 ( .IN1(conf8_9_), .IN2(n18065), .QN(n9334) );
  NAND2X0 U35084 ( .IN1(conf15_10_), .IN2(n17949), .QN(n14282) );
  NAND2X0 U35085 ( .IN1(conf6_11_), .IN2(n17941), .QN(n13356) );
  NAND2X0 U35086 ( .IN1(conf5_11_), .IN2(n18071), .QN(n13047) );
  NAND2X0 U35087 ( .IN1(conf13_11_), .IN2(n18072), .QN(n10881) );
  NAND2X0 U35088 ( .IN1(conf3_11_), .IN2(n18067), .QN(n12429) );
  NAND2X0 U35089 ( .IN1(conf11_11_), .IN2(n18073), .QN(n10262) );
  NAND2X0 U35090 ( .IN1(conf1_11_), .IN2(n18074), .QN(n11810) );
  NAND2X0 U35091 ( .IN1(conf9_11_), .IN2(n18068), .QN(n9642) );
  NAND2X0 U35092 ( .IN1(conf7_11_), .IN2(n18069), .QN(n13665) );
  NAND2X0 U35093 ( .IN1(conf14_11_), .IN2(n17942), .QN(n11190) );
  NAND2X0 U35094 ( .IN1(conf4_11_), .IN2(n17953), .QN(n12738) );
  NAND2X0 U35095 ( .IN1(conf12_11_), .IN2(n17954), .QN(n10571) );
  NAND2X0 U35096 ( .IN1(conf2_11_), .IN2(n17943), .QN(n12120) );
  NAND2X0 U35097 ( .IN1(conf10_11_), .IN2(n17955), .QN(n9952) );
  NAND2X0 U35098 ( .IN1(conf0_11_), .IN2(n17956), .QN(n11500) );
  NAND2X0 U35099 ( .IN1(conf8_11_), .IN2(n17944), .QN(n9331) );
  NAND2X0 U35100 ( .IN1(conf7_10_), .IN2(n17950), .QN(n13664) );
  NAND2X0 U35101 ( .IN1(conf6_10_), .IN2(n18075), .QN(n13355) );
  NAND2X0 U35102 ( .IN1(conf14_10_), .IN2(n18076), .QN(n11189) );
  NAND2X0 U35103 ( .IN1(conf5_10_), .IN2(n17960), .QN(n13046) );
  NAND2X0 U35104 ( .IN1(conf4_10_), .IN2(n18079), .QN(n12737) );
  NAND2X0 U35105 ( .IN1(conf13_10_), .IN2(n17961), .QN(n10880) );
  NAND2X0 U35106 ( .IN1(conf12_10_), .IN2(n18080), .QN(n10570) );
  NAND2X0 U35107 ( .IN1(conf3_10_), .IN2(n17951), .QN(n12428) );
  NAND2X0 U35108 ( .IN1(conf2_10_), .IN2(n18077), .QN(n12119) );
  NAND2X0 U35109 ( .IN1(conf11_10_), .IN2(n17962), .QN(n10261) );
  NAND2X0 U35110 ( .IN1(conf10_10_), .IN2(n18081), .QN(n9951) );
  NAND2X0 U35111 ( .IN1(conf1_10_), .IN2(n17963), .QN(n11809) );
  NAND2X0 U35112 ( .IN1(conf0_10_), .IN2(n18082), .QN(n11499) );
  NAND2X0 U35113 ( .IN1(conf9_10_), .IN2(n17952), .QN(n9641) );
  NAND2X0 U35114 ( .IN1(conf8_10_), .IN2(n18078), .QN(n9330) );
  NAND2X0 U35115 ( .IN1(conf15_11_), .IN2(n18070), .QN(n14300) );
  AO22X1 U35116 ( .IN1(n14330), .IN2(m4s15_cyc), .IN3(n14331), .IN4(n17788), 
        .Q(n17699) );
  INVX0 U35117 ( .IN(m7_addr_i[28]), .QN(n2277) );
  INVX0 U35118 ( .IN(m5_addr_i[28]), .QN(n2105) );
  INVX0 U35119 ( .IN(m3_addr_i[28]), .QN(n1933) );
  INVX0 U35120 ( .IN(m1_addr_i[28]), .QN(n1761) );
  INVX0 U35121 ( .IN(m7_addr_i[29]), .QN(n2276) );
  INVX0 U35122 ( .IN(m5_addr_i[29]), .QN(n2104) );
  INVX0 U35123 ( .IN(m3_addr_i[29]), .QN(n1932) );
  INVX0 U35124 ( .IN(m1_addr_i[29]), .QN(n1760) );
  INVX0 U35125 ( .IN(m7_addr_i[30]), .QN(n2275) );
  INVX0 U35126 ( .IN(m5_addr_i[30]), .QN(n2103) );
  INVX0 U35127 ( .IN(m3_addr_i[30]), .QN(n1931) );
  INVX0 U35128 ( .IN(m1_addr_i[30]), .QN(n1759) );
  INVX0 U35129 ( .IN(m6_addr_i[28]), .QN(n2191) );
  INVX0 U35130 ( .IN(m4_addr_i[28]), .QN(n2019) );
  INVX0 U35131 ( .IN(m2_addr_i[28]), .QN(n1847) );
  INVX0 U35132 ( .IN(m0_addr_i[28]), .QN(n1657) );
  INVX0 U35133 ( .IN(m7_addr_i[31]), .QN(n2274) );
  INVX0 U35134 ( .IN(m5_addr_i[31]), .QN(n2102) );
  INVX0 U35135 ( .IN(m3_addr_i[31]), .QN(n1930) );
  INVX0 U35136 ( .IN(m1_addr_i[31]), .QN(n1758) );
  INVX0 U35137 ( .IN(m6_addr_i[29]), .QN(n2190) );
  INVX0 U35138 ( .IN(m4_addr_i[29]), .QN(n2018) );
  INVX0 U35139 ( .IN(m2_addr_i[29]), .QN(n1846) );
  INVX0 U35140 ( .IN(m0_addr_i[29]), .QN(n1656) );
  INVX0 U35141 ( .IN(m6_addr_i[30]), .QN(n2189) );
  INVX0 U35142 ( .IN(m4_addr_i[30]), .QN(n2017) );
  INVX0 U35143 ( .IN(m2_addr_i[30]), .QN(n1845) );
  INVX0 U35144 ( .IN(m0_addr_i[30]), .QN(n1655) );
  INVX0 U35145 ( .IN(m6_addr_i[31]), .QN(n2188) );
  INVX0 U35146 ( .IN(m4_addr_i[31]), .QN(n2016) );
  INVX0 U35147 ( .IN(m2_addr_i[31]), .QN(n1844) );
  INVX0 U35148 ( .IN(m0_addr_i[31]), .QN(n1650) );
  NAND3X0 U35149 ( .IN1(n3859), .IN2(n3861), .IN3(s7_msel_gnt_p0_1_), .QN(
        n13771) );
  NAND3X0 U35150 ( .IN1(n3814), .IN2(n3816), .IN3(s6_msel_gnt_p0[1]), .QN(
        n13462) );
  NAND3X0 U35151 ( .IN1(n4174), .IN2(n4176), .IN3(test_so94), .QN(n11296) );
  NAND3X0 U35152 ( .IN1(n3769), .IN2(n3771), .IN3(s5_msel_gnt_p0[1]), .QN(
        n13153) );
  NAND3X0 U35153 ( .IN1(n3724), .IN2(n3726), .IN3(s4_msel_gnt_p0[1]), .QN(
        n12844) );
  NAND3X0 U35154 ( .IN1(n4129), .IN2(n4131), .IN3(s13_msel_gnt_p0_1_), .QN(
        n10987) );
  NAND3X0 U35155 ( .IN1(n4084), .IN2(n4086), .IN3(s12_msel_gnt_p0[1]), .QN(
        n10677) );
  NAND3X0 U35156 ( .IN1(n3679), .IN2(n3681), .IN3(s3_msel_gnt_p0_1_), .QN(
        n12535) );
  NAND3X0 U35157 ( .IN1(n3634), .IN2(n3636), .IN3(test_so48), .QN(n12226) );
  NAND3X0 U35158 ( .IN1(n4039), .IN2(n4041), .IN3(s11_msel_gnt_p0[1]), .QN(
        n10368) );
  NAND3X0 U35159 ( .IN1(n3994), .IN2(n3996), .IN3(s10_msel_gnt_p0[1]), .QN(
        n10058) );
  NAND3X0 U35160 ( .IN1(n3589), .IN2(n3591), .IN3(s1_msel_gnt_p0_1_), .QN(
        n11916) );
  NAND3X0 U35161 ( .IN1(n3544), .IN2(n3546), .IN3(s0_msel_gnt_p0[1]), .QN(
        n11606) );
  NAND3X0 U35162 ( .IN1(n3949), .IN2(n3951), .IN3(s9_msel_gnt_p0_1_), .QN(
        n9748) );
  NAND3X0 U35163 ( .IN1(n3904), .IN2(n3906), .IN3(test_so71), .QN(n9437) );
  NAND3X0 U35164 ( .IN1(n4219), .IN2(n4221), .IN3(s15_msel_gnt_p0_1_), .QN(
        n14035) );
  NAND3X0 U35165 ( .IN1(s7_msel_gnt_p0_1_), .IN2(n3861), .IN3(test_so67), .QN(
        n13752) );
  NAND3X0 U35166 ( .IN1(s6_msel_gnt_p0[1]), .IN2(n3816), .IN3(
        s6_msel_gnt_p0[0]), .QN(n13443) );
  NAND3X0 U35167 ( .IN1(test_so94), .IN2(n4176), .IN3(s14_msel_gnt_p0_0_), 
        .QN(n11277) );
  NAND3X0 U35168 ( .IN1(s5_msel_gnt_p0[1]), .IN2(n3771), .IN3(
        s5_msel_gnt_p0[0]), .QN(n13134) );
  NAND3X0 U35169 ( .IN1(s4_msel_gnt_p0[1]), .IN2(n3726), .IN3(
        s4_msel_gnt_p0[0]), .QN(n12825) );
  NAND3X0 U35170 ( .IN1(s13_msel_gnt_p0_1_), .IN2(n4131), .IN3(test_so90), 
        .QN(n10968) );
  NAND3X0 U35171 ( .IN1(s12_msel_gnt_p0[1]), .IN2(n4086), .IN3(
        s12_msel_gnt_p0[0]), .QN(n10658) );
  NAND3X0 U35172 ( .IN1(s3_msel_gnt_p0_1_), .IN2(n3681), .IN3(
        s3_msel_gnt_p0_0_), .QN(n12516) );
  NAND3X0 U35173 ( .IN1(test_so48), .IN2(n3636), .IN3(s2_msel_gnt_p0_0_), .QN(
        n12207) );
  NAND3X0 U35174 ( .IN1(s11_msel_gnt_p0[1]), .IN2(n4041), .IN3(
        s11_msel_gnt_p0[0]), .QN(n10349) );
  NAND3X0 U35175 ( .IN1(s10_msel_gnt_p0[1]), .IN2(n3996), .IN3(
        s10_msel_gnt_p0[0]), .QN(n10039) );
  NAND3X0 U35176 ( .IN1(s1_msel_gnt_p0_1_), .IN2(n3591), .IN3(test_so44), .QN(
        n11897) );
  NAND3X0 U35177 ( .IN1(s0_msel_gnt_p0[1]), .IN2(n3546), .IN3(
        s0_msel_gnt_p0[0]), .QN(n11587) );
  NAND3X0 U35178 ( .IN1(s9_msel_gnt_p0_1_), .IN2(n3951), .IN3(
        s9_msel_gnt_p0_0_), .QN(n9729) );
  NAND3X0 U35179 ( .IN1(test_so71), .IN2(n3906), .IN3(s8_msel_gnt_p0_0_), .QN(
        n9418) );
  NAND3X0 U35180 ( .IN1(s15_msel_gnt_p0_1_), .IN2(n4221), .IN3(
        s15_msel_gnt_p0_0_), .QN(n14016) );
  ISOLANDX1 U35181 ( .D(test_so24), .ISO(n13641), .Q(n13754) );
  ISOLANDX1 U35182 ( .D(m3s6_cyc), .ISO(n13332), .Q(n13445) );
  ISOLANDX1 U35183 ( .D(test_so25), .ISO(n11166), .Q(n11279) );
  ISOLANDX1 U35184 ( .D(m3s5_cyc), .ISO(n13023), .Q(n13136) );
  ISOLANDX1 U35185 ( .D(m3s4_cyc), .ISO(n12714), .Q(n12827) );
  ISOLANDX1 U35186 ( .D(m3s13_cyc), .ISO(n10857), .Q(n10970) );
  ISOLANDX1 U35187 ( .D(m3s12_cyc), .ISO(n10547), .Q(n10660) );
  ISOLANDX1 U35188 ( .D(m3s3_cyc), .ISO(n12405), .Q(n12518) );
  ISOLANDX1 U35189 ( .D(m3s2_cyc), .ISO(n12096), .Q(n12209) );
  ISOLANDX1 U35190 ( .D(m3s11_cyc), .ISO(n10238), .Q(n10351) );
  ISOLANDX1 U35191 ( .D(m3s10_cyc), .ISO(n9928), .Q(n10041) );
  ISOLANDX1 U35192 ( .D(m3s1_cyc), .ISO(n11786), .Q(n11899) );
  ISOLANDX1 U35193 ( .D(test_so23), .ISO(n11476), .Q(n11589) );
  ISOLANDX1 U35194 ( .D(m3s9_cyc), .ISO(n9618), .Q(n9731) );
  ISOLANDX1 U35195 ( .D(m3s8_cyc), .ISO(n9307), .Q(n9420) );
  ISOLANDX1 U35196 ( .D(m3s15_cyc), .ISO(n14073), .Q(n14018) );
  INVX0 U35197 ( .IN(m7_stb_i), .QN(n2311) );
  INVX0 U35198 ( .IN(m5_stb_i), .QN(n2139) );
  INVX0 U35199 ( .IN(m3_stb_i), .QN(n1967) );
  INVX0 U35200 ( .IN(m1_stb_i), .QN(n1795) );
  INVX0 U35201 ( .IN(m6_stb_i), .QN(n2225) );
  INVX0 U35202 ( .IN(m4_stb_i), .QN(n2053) );
  INVX0 U35203 ( .IN(m2_stb_i), .QN(n1881) );
  INVX0 U35204 ( .IN(m0_stb_i), .QN(n1709) );
  INVX0 U35205 ( .IN(m7_addr_i[24]), .QN(n2281) );
  INVX0 U35206 ( .IN(m5_addr_i[24]), .QN(n2109) );
  INVX0 U35207 ( .IN(m3_addr_i[24]), .QN(n1937) );
  INVX0 U35208 ( .IN(m1_addr_i[24]), .QN(n1765) );
  INVX0 U35209 ( .IN(m7_addr_i[25]), .QN(n2280) );
  INVX0 U35210 ( .IN(m5_addr_i[25]), .QN(n2108) );
  INVX0 U35211 ( .IN(m3_addr_i[25]), .QN(n1936) );
  INVX0 U35212 ( .IN(m1_addr_i[25]), .QN(n1764) );
  INVX0 U35213 ( .IN(m7_addr_i[26]), .QN(n2279) );
  INVX0 U35214 ( .IN(m5_addr_i[26]), .QN(n2107) );
  INVX0 U35215 ( .IN(m3_addr_i[26]), .QN(n1935) );
  INVX0 U35216 ( .IN(m1_addr_i[26]), .QN(n1763) );
  INVX0 U35217 ( .IN(m7_addr_i[27]), .QN(n2278) );
  INVX0 U35218 ( .IN(m5_addr_i[27]), .QN(n2106) );
  INVX0 U35219 ( .IN(m3_addr_i[27]), .QN(n1934) );
  INVX0 U35220 ( .IN(m1_addr_i[27]), .QN(n1762) );
  INVX0 U35221 ( .IN(m6_addr_i[24]), .QN(n2195) );
  INVX0 U35222 ( .IN(m4_addr_i[24]), .QN(n2023) );
  INVX0 U35223 ( .IN(m2_addr_i[24]), .QN(n1851) );
  INVX0 U35224 ( .IN(m0_addr_i[24]), .QN(n1661) );
  INVX0 U35225 ( .IN(m6_addr_i[25]), .QN(n2194) );
  INVX0 U35226 ( .IN(m4_addr_i[25]), .QN(n2022) );
  INVX0 U35227 ( .IN(m2_addr_i[25]), .QN(n1850) );
  INVX0 U35228 ( .IN(m0_addr_i[25]), .QN(n1660) );
  INVX0 U35229 ( .IN(m6_addr_i[26]), .QN(n2193) );
  INVX0 U35230 ( .IN(m4_addr_i[26]), .QN(n2021) );
  INVX0 U35231 ( .IN(m2_addr_i[26]), .QN(n1849) );
  INVX0 U35232 ( .IN(m0_addr_i[26]), .QN(n1659) );
  INVX0 U35233 ( .IN(m6_addr_i[27]), .QN(n2192) );
  INVX0 U35234 ( .IN(m4_addr_i[27]), .QN(n2020) );
  INVX0 U35235 ( .IN(m2_addr_i[27]), .QN(n1848) );
  INVX0 U35236 ( .IN(m0_addr_i[27]), .QN(n1658) );
  AO22X1 U35237 ( .IN1(n18409), .IN2(n18341), .IN3(test_so14), .IN4(n1693), 
        .Q(n921) );
  AO22X1 U35238 ( .IN1(n18408), .IN2(n18343), .IN3(conf13_1_), .IN4(n1693), 
        .Q(n922) );
  AO22X1 U35239 ( .IN1(n18409), .IN2(n18345), .IN3(conf13_2_), .IN4(n1693), 
        .Q(n923) );
  AO22X1 U35240 ( .IN1(n18408), .IN2(n18347), .IN3(conf13_3_), .IN4(n1693), 
        .Q(n924) );
  AO22X1 U35241 ( .IN1(n18409), .IN2(n18349), .IN3(conf13_4_), .IN4(n1693), 
        .Q(n925) );
  AO22X1 U35242 ( .IN1(n18408), .IN2(n18351), .IN3(conf13_5_), .IN4(n1693), 
        .Q(n926) );
  AO22X1 U35243 ( .IN1(n18409), .IN2(n18353), .IN3(conf13_6_), .IN4(n1693), 
        .Q(n927) );
  AO22X1 U35244 ( .IN1(n18408), .IN2(n18355), .IN3(conf13_7_), .IN4(n1693), 
        .Q(n928) );
  AO22X1 U35245 ( .IN1(n18409), .IN2(n18357), .IN3(conf13_8_), .IN4(n1693), 
        .Q(n929) );
  AO22X1 U35246 ( .IN1(n18408), .IN2(n18359), .IN3(conf13_9_), .IN4(n1693), 
        .Q(n930) );
  AO22X1 U35247 ( .IN1(n18409), .IN2(n18361), .IN3(conf13_10_), .IN4(n1693), 
        .Q(n931) );
  AO22X1 U35248 ( .IN1(n18408), .IN2(n18363), .IN3(conf13_11_), .IN4(n1693), 
        .Q(n932) );
  AO22X1 U35249 ( .IN1(n18409), .IN2(n18365), .IN3(conf13_12_), .IN4(n1693), 
        .Q(n933) );
  AO22X1 U35250 ( .IN1(n18408), .IN2(n18367), .IN3(conf13_13_), .IN4(n1693), 
        .Q(n934) );
  AO22X1 U35251 ( .IN1(n18409), .IN2(n18369), .IN3(conf13_14_), .IN4(n1693), 
        .Q(n935) );
  AO22X1 U35252 ( .IN1(n18408), .IN2(n18339), .IN3(conf13_15_), .IN4(n1693), 
        .Q(n936) );
  AO22X1 U35253 ( .IN1(n18413), .IN2(n18341), .IN3(test_so13), .IN4(n1681), 
        .Q(n971) );
  AO22X1 U35254 ( .IN1(n18412), .IN2(n18343), .IN3(conf12_1_), .IN4(n1681), 
        .Q(n972) );
  AO22X1 U35255 ( .IN1(n18413), .IN2(n18345), .IN3(conf12_2_), .IN4(n1681), 
        .Q(n973) );
  AO22X1 U35256 ( .IN1(n18412), .IN2(n18347), .IN3(conf12_3_), .IN4(n1681), 
        .Q(n974) );
  AO22X1 U35257 ( .IN1(n18413), .IN2(n18349), .IN3(conf12_4_), .IN4(n1681), 
        .Q(n975) );
  AO22X1 U35258 ( .IN1(n18412), .IN2(n18351), .IN3(conf12_5_), .IN4(n1681), 
        .Q(n976) );
  AO22X1 U35259 ( .IN1(n18413), .IN2(n18353), .IN3(conf12_6_), .IN4(n1681), 
        .Q(n977) );
  AO22X1 U35260 ( .IN1(n18412), .IN2(n18355), .IN3(conf12_7_), .IN4(n1681), 
        .Q(n978) );
  AO22X1 U35261 ( .IN1(n18413), .IN2(n18357), .IN3(conf12_8_), .IN4(n1681), 
        .Q(n979) );
  AO22X1 U35262 ( .IN1(n18412), .IN2(n18359), .IN3(conf12_9_), .IN4(n1681), 
        .Q(n980) );
  AO22X1 U35263 ( .IN1(n18413), .IN2(n18361), .IN3(conf12_10_), .IN4(n1681), 
        .Q(n981) );
  AO22X1 U35264 ( .IN1(n18412), .IN2(n18363), .IN3(conf12_11_), .IN4(n1681), 
        .Q(n982) );
  AO22X1 U35265 ( .IN1(n18413), .IN2(n18365), .IN3(conf12_12_), .IN4(n1681), 
        .Q(n983) );
  AO22X1 U35266 ( .IN1(n18412), .IN2(n18367), .IN3(conf12_13_), .IN4(n1681), 
        .Q(n984) );
  AO22X1 U35267 ( .IN1(n18413), .IN2(n18369), .IN3(conf12_14_), .IN4(n1681), 
        .Q(n985) );
  AO22X1 U35268 ( .IN1(n18412), .IN2(n18339), .IN3(conf12_15_), .IN4(n1681), 
        .Q(n986) );
  AO22X1 U35269 ( .IN1(n18417), .IN2(n18341), .IN3(test_so12), .IN4(n1694), 
        .Q(n1021) );
  AO22X1 U35270 ( .IN1(n18416), .IN2(n18343), .IN3(conf11_1_), .IN4(n1694), 
        .Q(n1022) );
  AO22X1 U35271 ( .IN1(n18417), .IN2(n18345), .IN3(conf11_2_), .IN4(n1694), 
        .Q(n1023) );
  AO22X1 U35272 ( .IN1(n18416), .IN2(n18347), .IN3(conf11_3_), .IN4(n1694), 
        .Q(n1024) );
  AO22X1 U35273 ( .IN1(n18417), .IN2(n18349), .IN3(conf11_4_), .IN4(n1694), 
        .Q(n1025) );
  AO22X1 U35274 ( .IN1(n18416), .IN2(n18351), .IN3(conf11_5_), .IN4(n1694), 
        .Q(n1026) );
  AO22X1 U35275 ( .IN1(n18417), .IN2(n18353), .IN3(conf11_6_), .IN4(n1694), 
        .Q(n1027) );
  AO22X1 U35276 ( .IN1(n18416), .IN2(n18355), .IN3(conf11_7_), .IN4(n1694), 
        .Q(n1028) );
  AO22X1 U35277 ( .IN1(n18417), .IN2(n18357), .IN3(conf11_8_), .IN4(n1694), 
        .Q(n1029) );
  AO22X1 U35278 ( .IN1(n18416), .IN2(n18359), .IN3(conf11_9_), .IN4(n1694), 
        .Q(n1030) );
  AO22X1 U35279 ( .IN1(n18417), .IN2(n18361), .IN3(conf11_10_), .IN4(n1694), 
        .Q(n1031) );
  AO22X1 U35280 ( .IN1(n18416), .IN2(n18363), .IN3(conf11_11_), .IN4(n1694), 
        .Q(n1032) );
  AO22X1 U35281 ( .IN1(n18417), .IN2(n18365), .IN3(conf11_12_), .IN4(n1694), 
        .Q(n1033) );
  AO22X1 U35282 ( .IN1(n18416), .IN2(n18367), .IN3(conf11_13_), .IN4(n1694), 
        .Q(n1034) );
  AO22X1 U35283 ( .IN1(n18417), .IN2(n18369), .IN3(conf11_14_), .IN4(n1694), 
        .Q(n1035) );
  AO22X1 U35284 ( .IN1(n18416), .IN2(n18339), .IN3(conf11_15_), .IN4(n1694), 
        .Q(n1036) );
  AO22X1 U35285 ( .IN1(n18421), .IN2(n18341), .IN3(test_so11), .IN4(n1682), 
        .Q(n1071) );
  AO22X1 U35286 ( .IN1(n18420), .IN2(n18343), .IN3(conf10_1_), .IN4(n1682), 
        .Q(n1072) );
  AO22X1 U35287 ( .IN1(n18421), .IN2(n18345), .IN3(conf10_2_), .IN4(n1682), 
        .Q(n1073) );
  AO22X1 U35288 ( .IN1(n18420), .IN2(n18347), .IN3(conf10_3_), .IN4(n1682), 
        .Q(n1074) );
  AO22X1 U35289 ( .IN1(n18421), .IN2(n18349), .IN3(conf10_4_), .IN4(n1682), 
        .Q(n1075) );
  AO22X1 U35290 ( .IN1(n18420), .IN2(n18351), .IN3(conf10_5_), .IN4(n1682), 
        .Q(n1076) );
  AO22X1 U35291 ( .IN1(n18421), .IN2(n18353), .IN3(conf10_6_), .IN4(n1682), 
        .Q(n1077) );
  AO22X1 U35292 ( .IN1(n18420), .IN2(n18355), .IN3(conf10_7_), .IN4(n1682), 
        .Q(n1078) );
  AO22X1 U35293 ( .IN1(n18421), .IN2(n18357), .IN3(conf10_8_), .IN4(n1682), 
        .Q(n1079) );
  AO22X1 U35294 ( .IN1(n18420), .IN2(n18359), .IN3(conf10_9_), .IN4(n1682), 
        .Q(n1080) );
  AO22X1 U35295 ( .IN1(n18421), .IN2(n18361), .IN3(conf10_10_), .IN4(n1682), 
        .Q(n1081) );
  AO22X1 U35296 ( .IN1(n18420), .IN2(n18363), .IN3(conf10_11_), .IN4(n1682), 
        .Q(n1082) );
  AO22X1 U35297 ( .IN1(n18421), .IN2(n18365), .IN3(conf10_12_), .IN4(n1682), 
        .Q(n1083) );
  AO22X1 U35298 ( .IN1(n18420), .IN2(n18367), .IN3(conf10_13_), .IN4(n1682), 
        .Q(n1084) );
  AO22X1 U35299 ( .IN1(n18421), .IN2(n18369), .IN3(conf10_14_), .IN4(n1682), 
        .Q(n1085) );
  AO22X1 U35300 ( .IN1(n18420), .IN2(n18339), .IN3(conf10_15_), .IN4(n1682), 
        .Q(n1086) );
  AO22X1 U35301 ( .IN1(n18425), .IN2(n18341), .IN3(test_so10), .IN4(n1695), 
        .Q(n1121) );
  AO22X1 U35302 ( .IN1(n18424), .IN2(n18343), .IN3(conf9_1_), .IN4(n1695), .Q(
        n1122) );
  AO22X1 U35303 ( .IN1(n18425), .IN2(n18345), .IN3(conf9_2_), .IN4(n1695), .Q(
        n1123) );
  AO22X1 U35304 ( .IN1(n18424), .IN2(n18347), .IN3(conf9_3_), .IN4(n1695), .Q(
        n1124) );
  AO22X1 U35305 ( .IN1(n18425), .IN2(n18349), .IN3(conf9_4_), .IN4(n1695), .Q(
        n1125) );
  AO22X1 U35306 ( .IN1(n18424), .IN2(n18351), .IN3(conf9_5_), .IN4(n1695), .Q(
        n1126) );
  AO22X1 U35307 ( .IN1(n18425), .IN2(n18353), .IN3(conf9_6_), .IN4(n1695), .Q(
        n1127) );
  AO22X1 U35308 ( .IN1(n18424), .IN2(n18355), .IN3(conf9_7_), .IN4(n1695), .Q(
        n1128) );
  AO22X1 U35309 ( .IN1(n18425), .IN2(n18357), .IN3(conf9_8_), .IN4(n1695), .Q(
        n1129) );
  AO22X1 U35310 ( .IN1(n18424), .IN2(n18359), .IN3(conf9_9_), .IN4(n1695), .Q(
        n1130) );
  AO22X1 U35311 ( .IN1(n18425), .IN2(n18361), .IN3(conf9_10_), .IN4(n1695), 
        .Q(n1131) );
  AO22X1 U35312 ( .IN1(n18424), .IN2(n18363), .IN3(conf9_11_), .IN4(n1695), 
        .Q(n1132) );
  AO22X1 U35313 ( .IN1(n18425), .IN2(n18365), .IN3(conf9_12_), .IN4(n1695), 
        .Q(n1133) );
  AO22X1 U35314 ( .IN1(n18424), .IN2(n18367), .IN3(conf9_13_), .IN4(n1695), 
        .Q(n1134) );
  AO22X1 U35315 ( .IN1(n18425), .IN2(n18369), .IN3(conf9_14_), .IN4(n1695), 
        .Q(n1135) );
  AO22X1 U35316 ( .IN1(n18424), .IN2(n18339), .IN3(conf9_15_), .IN4(n1695), 
        .Q(n1136) );
  AO22X1 U35317 ( .IN1(n18429), .IN2(n18341), .IN3(test_so9), .IN4(n1683), .Q(
        n1171) );
  AO22X1 U35318 ( .IN1(n18428), .IN2(n18343), .IN3(conf8_1_), .IN4(n1683), .Q(
        n1172) );
  AO22X1 U35319 ( .IN1(n18429), .IN2(n18345), .IN3(conf8_2_), .IN4(n1683), .Q(
        n1173) );
  AO22X1 U35320 ( .IN1(n18428), .IN2(n18347), .IN3(conf8_3_), .IN4(n1683), .Q(
        n1174) );
  AO22X1 U35321 ( .IN1(n18429), .IN2(n18349), .IN3(conf8_4_), .IN4(n1683), .Q(
        n1175) );
  AO22X1 U35322 ( .IN1(n18428), .IN2(n18351), .IN3(conf8_5_), .IN4(n1683), .Q(
        n1176) );
  AO22X1 U35323 ( .IN1(n18429), .IN2(n18353), .IN3(conf8_6_), .IN4(n1683), .Q(
        n1177) );
  AO22X1 U35324 ( .IN1(n18428), .IN2(n18355), .IN3(conf8_7_), .IN4(n1683), .Q(
        n1178) );
  AO22X1 U35325 ( .IN1(n18429), .IN2(n18357), .IN3(conf8_8_), .IN4(n1683), .Q(
        n1179) );
  AO22X1 U35326 ( .IN1(n18428), .IN2(n18359), .IN3(conf8_9_), .IN4(n1683), .Q(
        n1180) );
  AO22X1 U35327 ( .IN1(n18429), .IN2(n18361), .IN3(conf8_10_), .IN4(n1683), 
        .Q(n1181) );
  AO22X1 U35328 ( .IN1(n18428), .IN2(n18363), .IN3(conf8_11_), .IN4(n1683), 
        .Q(n1182) );
  AO22X1 U35329 ( .IN1(n18429), .IN2(n18365), .IN3(conf8_12_), .IN4(n1683), 
        .Q(n1183) );
  AO22X1 U35330 ( .IN1(n18428), .IN2(n18367), .IN3(conf8_13_), .IN4(n1683), 
        .Q(n1184) );
  AO22X1 U35331 ( .IN1(n18429), .IN2(n18369), .IN3(conf8_14_), .IN4(n1683), 
        .Q(n1185) );
  AO22X1 U35332 ( .IN1(n18428), .IN2(n18339), .IN3(conf8_15_), .IN4(n1683), 
        .Q(n1186) );
  AO22X1 U35333 ( .IN1(n18373), .IN2(n18341), .IN3(test_so8), .IN4(n1688), .Q(
        n1221) );
  AO22X1 U35334 ( .IN1(n18372), .IN2(n18343), .IN3(conf7_1_), .IN4(n1688), .Q(
        n1222) );
  AO22X1 U35335 ( .IN1(n18373), .IN2(n18345), .IN3(conf7_2_), .IN4(n1688), .Q(
        n1223) );
  AO22X1 U35336 ( .IN1(n18372), .IN2(n18347), .IN3(conf7_3_), .IN4(n1688), .Q(
        n1224) );
  AO22X1 U35337 ( .IN1(n18373), .IN2(n18349), .IN3(conf7_4_), .IN4(n1688), .Q(
        n1225) );
  AO22X1 U35338 ( .IN1(n18372), .IN2(n18351), .IN3(conf7_5_), .IN4(n1688), .Q(
        n1226) );
  AO22X1 U35339 ( .IN1(n18373), .IN2(n18353), .IN3(conf7_6_), .IN4(n1688), .Q(
        n1227) );
  AO22X1 U35340 ( .IN1(n18372), .IN2(n18355), .IN3(conf7_7_), .IN4(n1688), .Q(
        n1228) );
  AO22X1 U35341 ( .IN1(n18373), .IN2(n18357), .IN3(conf7_8_), .IN4(n1688), .Q(
        n1229) );
  AO22X1 U35342 ( .IN1(n18372), .IN2(n18359), .IN3(conf7_9_), .IN4(n1688), .Q(
        n1230) );
  AO22X1 U35343 ( .IN1(n18373), .IN2(n18361), .IN3(conf7_10_), .IN4(n1688), 
        .Q(n1231) );
  AO22X1 U35344 ( .IN1(n18372), .IN2(n18363), .IN3(conf7_11_), .IN4(n1688), 
        .Q(n1232) );
  AO22X1 U35345 ( .IN1(n18373), .IN2(n18365), .IN3(conf7_12_), .IN4(n1688), 
        .Q(n1233) );
  AO22X1 U35346 ( .IN1(n18372), .IN2(n18367), .IN3(conf7_13_), .IN4(n1688), 
        .Q(n1234) );
  AO22X1 U35347 ( .IN1(n18373), .IN2(n18369), .IN3(conf7_14_), .IN4(n1688), 
        .Q(n1235) );
  AO22X1 U35348 ( .IN1(n18372), .IN2(n18339), .IN3(conf7_15_), .IN4(n1688), 
        .Q(n1236) );
  AO22X1 U35349 ( .IN1(n18377), .IN2(n18341), .IN3(test_so7), .IN4(n1684), .Q(
        n1271) );
  AO22X1 U35350 ( .IN1(n18376), .IN2(n18343), .IN3(conf6_1_), .IN4(n1684), .Q(
        n1272) );
  AO22X1 U35351 ( .IN1(n18377), .IN2(n18345), .IN3(conf6_2_), .IN4(n1684), .Q(
        n1273) );
  AO22X1 U35352 ( .IN1(n18376), .IN2(n18347), .IN3(conf6_3_), .IN4(n1684), .Q(
        n1274) );
  AO22X1 U35353 ( .IN1(n18377), .IN2(n18349), .IN3(conf6_4_), .IN4(n1684), .Q(
        n1275) );
  AO22X1 U35354 ( .IN1(n18376), .IN2(n18351), .IN3(conf6_5_), .IN4(n1684), .Q(
        n1276) );
  AO22X1 U35355 ( .IN1(n18377), .IN2(n18353), .IN3(conf6_6_), .IN4(n1684), .Q(
        n1277) );
  AO22X1 U35356 ( .IN1(n18376), .IN2(n18355), .IN3(conf6_7_), .IN4(n1684), .Q(
        n1278) );
  AO22X1 U35357 ( .IN1(n18377), .IN2(n18357), .IN3(conf6_8_), .IN4(n1684), .Q(
        n1279) );
  AO22X1 U35358 ( .IN1(n18376), .IN2(n18359), .IN3(conf6_9_), .IN4(n1684), .Q(
        n1280) );
  AO22X1 U35359 ( .IN1(n18377), .IN2(n18361), .IN3(conf6_10_), .IN4(n1684), 
        .Q(n1281) );
  AO22X1 U35360 ( .IN1(n18376), .IN2(n18363), .IN3(conf6_11_), .IN4(n1684), 
        .Q(n1282) );
  AO22X1 U35361 ( .IN1(n18377), .IN2(n18365), .IN3(conf6_12_), .IN4(n1684), 
        .Q(n1283) );
  AO22X1 U35362 ( .IN1(n18376), .IN2(n18367), .IN3(conf6_13_), .IN4(n1684), 
        .Q(n1284) );
  AO22X1 U35363 ( .IN1(n18377), .IN2(n18369), .IN3(conf6_14_), .IN4(n1684), 
        .Q(n1285) );
  AO22X1 U35364 ( .IN1(n18376), .IN2(n18339), .IN3(conf6_15_), .IN4(n1684), 
        .Q(n1286) );
  AO22X1 U35365 ( .IN1(n18381), .IN2(n18341), .IN3(test_so6), .IN4(n1689), .Q(
        n1321) );
  AO22X1 U35366 ( .IN1(n18380), .IN2(n18343), .IN3(conf5_1_), .IN4(n1689), .Q(
        n1322) );
  AO22X1 U35367 ( .IN1(n18381), .IN2(n18345), .IN3(conf5_2_), .IN4(n1689), .Q(
        n1323) );
  AO22X1 U35368 ( .IN1(n18380), .IN2(n18347), .IN3(conf5_3_), .IN4(n1689), .Q(
        n1324) );
  AO22X1 U35369 ( .IN1(n18381), .IN2(n18349), .IN3(conf5_4_), .IN4(n1689), .Q(
        n1325) );
  AO22X1 U35370 ( .IN1(n18380), .IN2(n18351), .IN3(conf5_5_), .IN4(n1689), .Q(
        n1326) );
  AO22X1 U35371 ( .IN1(n18381), .IN2(n18353), .IN3(conf5_6_), .IN4(n1689), .Q(
        n1327) );
  AO22X1 U35372 ( .IN1(n18380), .IN2(n18355), .IN3(conf5_7_), .IN4(n1689), .Q(
        n1328) );
  AO22X1 U35373 ( .IN1(n18381), .IN2(n18357), .IN3(conf5_8_), .IN4(n1689), .Q(
        n1329) );
  AO22X1 U35374 ( .IN1(n18380), .IN2(n18359), .IN3(conf5_9_), .IN4(n1689), .Q(
        n1330) );
  AO22X1 U35375 ( .IN1(n18381), .IN2(n18361), .IN3(conf5_10_), .IN4(n1689), 
        .Q(n1331) );
  AO22X1 U35376 ( .IN1(n18380), .IN2(n18363), .IN3(conf5_11_), .IN4(n1689), 
        .Q(n1332) );
  AO22X1 U35377 ( .IN1(n18381), .IN2(n18365), .IN3(conf5_12_), .IN4(n1689), 
        .Q(n1333) );
  AO22X1 U35378 ( .IN1(n18380), .IN2(n18367), .IN3(conf5_13_), .IN4(n1689), 
        .Q(n1334) );
  AO22X1 U35379 ( .IN1(n18381), .IN2(n18369), .IN3(conf5_14_), .IN4(n1689), 
        .Q(n1335) );
  AO22X1 U35380 ( .IN1(n18380), .IN2(n18339), .IN3(conf5_15_), .IN4(n1689), 
        .Q(n1336) );
  AO22X1 U35381 ( .IN1(n18385), .IN2(n18341), .IN3(test_so5), .IN4(n1685), .Q(
        n1371) );
  AO22X1 U35382 ( .IN1(n18384), .IN2(n18343), .IN3(conf4_1_), .IN4(n1685), .Q(
        n1372) );
  AO22X1 U35383 ( .IN1(n18385), .IN2(n18345), .IN3(conf4_2_), .IN4(n1685), .Q(
        n1373) );
  AO22X1 U35384 ( .IN1(n18384), .IN2(n18347), .IN3(conf4_3_), .IN4(n1685), .Q(
        n1374) );
  AO22X1 U35385 ( .IN1(n18385), .IN2(n18349), .IN3(conf4_4_), .IN4(n1685), .Q(
        n1375) );
  AO22X1 U35386 ( .IN1(n18384), .IN2(n18351), .IN3(conf4_5_), .IN4(n1685), .Q(
        n1376) );
  AO22X1 U35387 ( .IN1(n18385), .IN2(n18353), .IN3(conf4_6_), .IN4(n1685), .Q(
        n1377) );
  AO22X1 U35388 ( .IN1(n18384), .IN2(n18355), .IN3(conf4_7_), .IN4(n1685), .Q(
        n1378) );
  AO22X1 U35389 ( .IN1(n18385), .IN2(n18357), .IN3(conf4_8_), .IN4(n1685), .Q(
        n1379) );
  AO22X1 U35390 ( .IN1(n18384), .IN2(n18359), .IN3(conf4_9_), .IN4(n1685), .Q(
        n1380) );
  AO22X1 U35391 ( .IN1(n18385), .IN2(n18361), .IN3(conf4_10_), .IN4(n1685), 
        .Q(n1381) );
  AO22X1 U35392 ( .IN1(n18384), .IN2(n18363), .IN3(conf4_11_), .IN4(n1685), 
        .Q(n1382) );
  AO22X1 U35393 ( .IN1(n18385), .IN2(n18365), .IN3(conf4_12_), .IN4(n1685), 
        .Q(n1383) );
  AO22X1 U35394 ( .IN1(n18384), .IN2(n18367), .IN3(conf4_13_), .IN4(n1685), 
        .Q(n1384) );
  AO22X1 U35395 ( .IN1(n18385), .IN2(n18369), .IN3(conf4_14_), .IN4(n1685), 
        .Q(n1385) );
  AO22X1 U35396 ( .IN1(n18384), .IN2(n18339), .IN3(conf4_15_), .IN4(n1685), 
        .Q(n1386) );
  AO22X1 U35397 ( .IN1(n18389), .IN2(n18341), .IN3(test_so4), .IN4(n1690), .Q(
        n1421) );
  AO22X1 U35398 ( .IN1(n18388), .IN2(n18343), .IN3(conf3_1_), .IN4(n1690), .Q(
        n1422) );
  AO22X1 U35399 ( .IN1(n18389), .IN2(n18345), .IN3(conf3_2_), .IN4(n1690), .Q(
        n1423) );
  AO22X1 U35400 ( .IN1(n18388), .IN2(n18347), .IN3(conf3_3_), .IN4(n1690), .Q(
        n1424) );
  AO22X1 U35401 ( .IN1(n18389), .IN2(n18349), .IN3(conf3_4_), .IN4(n1690), .Q(
        n1425) );
  AO22X1 U35402 ( .IN1(n18388), .IN2(n18351), .IN3(conf3_5_), .IN4(n1690), .Q(
        n1426) );
  AO22X1 U35403 ( .IN1(n18389), .IN2(n18353), .IN3(conf3_6_), .IN4(n1690), .Q(
        n1427) );
  AO22X1 U35404 ( .IN1(n18388), .IN2(n18355), .IN3(conf3_7_), .IN4(n1690), .Q(
        n1428) );
  AO22X1 U35405 ( .IN1(n18389), .IN2(n18357), .IN3(conf3_8_), .IN4(n1690), .Q(
        n1429) );
  AO22X1 U35406 ( .IN1(n18388), .IN2(n18359), .IN3(conf3_9_), .IN4(n1690), .Q(
        n1430) );
  AO22X1 U35407 ( .IN1(n18389), .IN2(n18361), .IN3(conf3_10_), .IN4(n1690), 
        .Q(n1431) );
  AO22X1 U35408 ( .IN1(n18388), .IN2(n18363), .IN3(conf3_11_), .IN4(n1690), 
        .Q(n1432) );
  AO22X1 U35409 ( .IN1(n18389), .IN2(n18365), .IN3(conf3_12_), .IN4(n1690), 
        .Q(n1433) );
  AO22X1 U35410 ( .IN1(n18388), .IN2(n18367), .IN3(conf3_13_), .IN4(n1690), 
        .Q(n1434) );
  AO22X1 U35411 ( .IN1(n18389), .IN2(n18369), .IN3(conf3_14_), .IN4(n1690), 
        .Q(n1435) );
  AO22X1 U35412 ( .IN1(n18388), .IN2(n18339), .IN3(conf3_15_), .IN4(n1690), 
        .Q(n1436) );
  AO22X1 U35413 ( .IN1(n18393), .IN2(n18341), .IN3(test_so3), .IN4(n1686), .Q(
        n1471) );
  AO22X1 U35414 ( .IN1(n18392), .IN2(n18343), .IN3(conf2_1_), .IN4(n1686), .Q(
        n1472) );
  AO22X1 U35415 ( .IN1(n18393), .IN2(n18345), .IN3(conf2_2_), .IN4(n1686), .Q(
        n1473) );
  AO22X1 U35416 ( .IN1(n18392), .IN2(n18347), .IN3(conf2_3_), .IN4(n1686), .Q(
        n1474) );
  AO22X1 U35417 ( .IN1(n18393), .IN2(n18349), .IN3(conf2_4_), .IN4(n1686), .Q(
        n1475) );
  AO22X1 U35418 ( .IN1(n18392), .IN2(n18351), .IN3(conf2_5_), .IN4(n1686), .Q(
        n1476) );
  AO22X1 U35419 ( .IN1(n18393), .IN2(n18353), .IN3(conf2_6_), .IN4(n1686), .Q(
        n1477) );
  AO22X1 U35420 ( .IN1(n18392), .IN2(n18355), .IN3(conf2_7_), .IN4(n1686), .Q(
        n1478) );
  AO22X1 U35421 ( .IN1(n18393), .IN2(n18357), .IN3(conf2_8_), .IN4(n1686), .Q(
        n1479) );
  AO22X1 U35422 ( .IN1(n18392), .IN2(n18359), .IN3(conf2_9_), .IN4(n1686), .Q(
        n1480) );
  AO22X1 U35423 ( .IN1(n18393), .IN2(n18361), .IN3(conf2_10_), .IN4(n1686), 
        .Q(n1481) );
  AO22X1 U35424 ( .IN1(n18392), .IN2(n18363), .IN3(conf2_11_), .IN4(n1686), 
        .Q(n1482) );
  AO22X1 U35425 ( .IN1(n18393), .IN2(n18365), .IN3(conf2_12_), .IN4(n1686), 
        .Q(n1483) );
  AO22X1 U35426 ( .IN1(n18392), .IN2(n18367), .IN3(conf2_13_), .IN4(n1686), 
        .Q(n1484) );
  AO22X1 U35427 ( .IN1(n18393), .IN2(n18369), .IN3(conf2_14_), .IN4(n1686), 
        .Q(n1485) );
  AO22X1 U35428 ( .IN1(n18392), .IN2(n18339), .IN3(conf2_15_), .IN4(n1686), 
        .Q(n1486) );
  AO22X1 U35429 ( .IN1(n18397), .IN2(n18341), .IN3(test_so2), .IN4(n1691), .Q(
        n1521) );
  AO22X1 U35430 ( .IN1(n18396), .IN2(n18343), .IN3(conf1_1_), .IN4(n1691), .Q(
        n1522) );
  AO22X1 U35431 ( .IN1(n18397), .IN2(n18345), .IN3(conf1_2_), .IN4(n1691), .Q(
        n1523) );
  AO22X1 U35432 ( .IN1(n18396), .IN2(n18347), .IN3(conf1_3_), .IN4(n1691), .Q(
        n1524) );
  AO22X1 U35433 ( .IN1(n18397), .IN2(n18349), .IN3(conf1_4_), .IN4(n1691), .Q(
        n1525) );
  AO22X1 U35434 ( .IN1(n18396), .IN2(n18351), .IN3(conf1_5_), .IN4(n1691), .Q(
        n1526) );
  AO22X1 U35435 ( .IN1(n18397), .IN2(n18353), .IN3(conf1_6_), .IN4(n1691), .Q(
        n1527) );
  AO22X1 U35436 ( .IN1(n18396), .IN2(n18355), .IN3(conf1_7_), .IN4(n1691), .Q(
        n1528) );
  AO22X1 U35437 ( .IN1(n18397), .IN2(n18357), .IN3(conf1_8_), .IN4(n1691), .Q(
        n1529) );
  AO22X1 U35438 ( .IN1(n18396), .IN2(n18359), .IN3(conf1_9_), .IN4(n1691), .Q(
        n1530) );
  AO22X1 U35439 ( .IN1(n18397), .IN2(n18361), .IN3(conf1_10_), .IN4(n1691), 
        .Q(n1531) );
  AO22X1 U35440 ( .IN1(n18396), .IN2(n18363), .IN3(conf1_11_), .IN4(n1691), 
        .Q(n1532) );
  AO22X1 U35441 ( .IN1(n18397), .IN2(n18365), .IN3(conf1_12_), .IN4(n1691), 
        .Q(n1533) );
  AO22X1 U35442 ( .IN1(n18396), .IN2(n18367), .IN3(conf1_13_), .IN4(n1691), 
        .Q(n1534) );
  AO22X1 U35443 ( .IN1(n18397), .IN2(n18369), .IN3(conf1_14_), .IN4(n1691), 
        .Q(n1535) );
  AO22X1 U35444 ( .IN1(n18396), .IN2(n18339), .IN3(conf1_15_), .IN4(n1691), 
        .Q(n1536) );
  AO22X1 U35445 ( .IN1(n18401), .IN2(n18341), .IN3(test_so1), .IN4(n1687), .Q(
        n1571) );
  AO22X1 U35446 ( .IN1(n18400), .IN2(n18343), .IN3(conf0_1_), .IN4(n1687), .Q(
        n1572) );
  AO22X1 U35447 ( .IN1(n18401), .IN2(n18345), .IN3(conf0_2_), .IN4(n1687), .Q(
        n1573) );
  AO22X1 U35448 ( .IN1(n18400), .IN2(n18347), .IN3(conf0_3_), .IN4(n1687), .Q(
        n1574) );
  AO22X1 U35449 ( .IN1(n18401), .IN2(n18349), .IN3(conf0_4_), .IN4(n1687), .Q(
        n1575) );
  AO22X1 U35450 ( .IN1(n18400), .IN2(n18351), .IN3(conf0_5_), .IN4(n1687), .Q(
        n1576) );
  AO22X1 U35451 ( .IN1(n18401), .IN2(n18353), .IN3(conf0_6_), .IN4(n1687), .Q(
        n1577) );
  AO22X1 U35452 ( .IN1(n18400), .IN2(n18355), .IN3(conf0_7_), .IN4(n1687), .Q(
        n1578) );
  AO22X1 U35453 ( .IN1(n18401), .IN2(n18357), .IN3(conf0_8_), .IN4(n1687), .Q(
        n1579) );
  AO22X1 U35454 ( .IN1(n18400), .IN2(n18359), .IN3(conf0_9_), .IN4(n1687), .Q(
        n1580) );
  AO22X1 U35455 ( .IN1(n18401), .IN2(n18361), .IN3(conf0_10_), .IN4(n1687), 
        .Q(n1581) );
  AO22X1 U35456 ( .IN1(n18400), .IN2(n18363), .IN3(conf0_11_), .IN4(n1687), 
        .Q(n1582) );
  AO22X1 U35457 ( .IN1(n18401), .IN2(n18365), .IN3(conf0_12_), .IN4(n1687), 
        .Q(n1583) );
  AO22X1 U35458 ( .IN1(n18400), .IN2(n18367), .IN3(conf0_13_), .IN4(n1687), 
        .Q(n1584) );
  AO22X1 U35459 ( .IN1(n18401), .IN2(n18369), .IN3(conf0_14_), .IN4(n1687), 
        .Q(n1585) );
  AO22X1 U35460 ( .IN1(n18400), .IN2(n18339), .IN3(conf0_15_), .IN4(n1687), 
        .Q(n1586) );
  AO22X1 U35461 ( .IN1(n18337), .IN2(s15_data_o[0]), .IN3(test_so16), .IN4(
        n1692), .Q(n821) );
  AO22X1 U35462 ( .IN1(n18336), .IN2(s15_data_o[1]), .IN3(conf15_1_), .IN4(
        n1692), .Q(n822) );
  AO22X1 U35463 ( .IN1(n18337), .IN2(s15_data_o[2]), .IN3(conf15_2_), .IN4(
        n1692), .Q(n823) );
  AO22X1 U35464 ( .IN1(n18336), .IN2(s15_data_o[3]), .IN3(conf15_3_), .IN4(
        n1692), .Q(n824) );
  AO22X1 U35465 ( .IN1(n18337), .IN2(s15_data_o[4]), .IN3(conf15_4_), .IN4(
        n1692), .Q(n825) );
  AO22X1 U35466 ( .IN1(n18336), .IN2(s15_data_o[5]), .IN3(conf15_5_), .IN4(
        n1692), .Q(n826) );
  AO22X1 U35467 ( .IN1(n18337), .IN2(s15_data_o[6]), .IN3(conf15_6_), .IN4(
        n1692), .Q(n827) );
  AO22X1 U35468 ( .IN1(n18336), .IN2(s15_data_o[7]), .IN3(conf15_7_), .IN4(
        n1692), .Q(n828) );
  AO22X1 U35469 ( .IN1(n18337), .IN2(s15_data_o[8]), .IN3(conf15_8_), .IN4(
        n1692), .Q(n829) );
  AO22X1 U35470 ( .IN1(n18336), .IN2(s15_data_o[9]), .IN3(conf15_9_), .IN4(
        n1692), .Q(n830) );
  AO22X1 U35471 ( .IN1(n18337), .IN2(s15_data_o[10]), .IN3(conf15_10_), .IN4(
        n1692), .Q(n831) );
  AO22X1 U35472 ( .IN1(n18336), .IN2(s15_data_o[11]), .IN3(conf15_11_), .IN4(
        n1692), .Q(n832) );
  AO22X1 U35473 ( .IN1(n18337), .IN2(s15_data_o[12]), .IN3(conf15_12_), .IN4(
        n1692), .Q(n833) );
  AO22X1 U35474 ( .IN1(n18336), .IN2(s15_data_o[13]), .IN3(conf15_13_), .IN4(
        n1692), .Q(n834) );
  AO22X1 U35475 ( .IN1(n18337), .IN2(s15_data_o[14]), .IN3(conf15_14_), .IN4(
        n1692), .Q(n835) );
  AO22X1 U35476 ( .IN1(n18336), .IN2(s15_data_o[15]), .IN3(conf15_15_), .IN4(
        n1692), .Q(n836) );
  AO22X1 U35477 ( .IN1(n18405), .IN2(s15_data_o[0]), .IN3(test_so15), .IN4(
        n1680), .Q(n871) );
  AO22X1 U35478 ( .IN1(n18404), .IN2(s15_data_o[1]), .IN3(conf14_1_), .IN4(
        n1680), .Q(n872) );
  AO22X1 U35479 ( .IN1(n18405), .IN2(s15_data_o[2]), .IN3(conf14_2_), .IN4(
        n1680), .Q(n873) );
  AO22X1 U35480 ( .IN1(n18404), .IN2(s15_data_o[3]), .IN3(conf14_3_), .IN4(
        n1680), .Q(n874) );
  AO22X1 U35481 ( .IN1(n18405), .IN2(s15_data_o[4]), .IN3(conf14_4_), .IN4(
        n1680), .Q(n875) );
  AO22X1 U35482 ( .IN1(n18404), .IN2(s15_data_o[5]), .IN3(conf14_5_), .IN4(
        n1680), .Q(n876) );
  AO22X1 U35483 ( .IN1(n18405), .IN2(s15_data_o[6]), .IN3(conf14_6_), .IN4(
        n1680), .Q(n877) );
  AO22X1 U35484 ( .IN1(n18404), .IN2(s15_data_o[7]), .IN3(conf14_7_), .IN4(
        n1680), .Q(n878) );
  AO22X1 U35485 ( .IN1(n18405), .IN2(s15_data_o[8]), .IN3(conf14_8_), .IN4(
        n1680), .Q(n879) );
  AO22X1 U35486 ( .IN1(n18404), .IN2(s15_data_o[9]), .IN3(conf14_9_), .IN4(
        n1680), .Q(n880) );
  AO22X1 U35487 ( .IN1(n18405), .IN2(s15_data_o[10]), .IN3(conf14_10_), .IN4(
        n1680), .Q(n881) );
  AO22X1 U35488 ( .IN1(n18404), .IN2(s15_data_o[11]), .IN3(conf14_11_), .IN4(
        n1680), .Q(n882) );
  AO22X1 U35489 ( .IN1(n18405), .IN2(s15_data_o[12]), .IN3(conf14_12_), .IN4(
        n1680), .Q(n883) );
  AO22X1 U35490 ( .IN1(n18404), .IN2(s15_data_o[13]), .IN3(conf14_13_), .IN4(
        n1680), .Q(n884) );
  AO22X1 U35491 ( .IN1(n18405), .IN2(s15_data_o[14]), .IN3(conf14_14_), .IN4(
        n1680), .Q(n885) );
  AO22X1 U35492 ( .IN1(n18404), .IN2(s15_data_o[15]), .IN3(conf14_15_), .IN4(
        n1680), .Q(n886) );
  NAND4X0 U35493 ( .IN1(m4s15_cyc), .IN2(n14301), .IN3(n14070), .IN4(n14277), 
        .QN(n14294) );
  NAND3X0 U35494 ( .IN1(m7s15_cyc), .IN2(n19744), .IN3(s15_m7_cyc_r), .QN(
        n17104) );
  NAND3X0 U35495 ( .IN1(m3s15_cyc), .IN2(n19678), .IN3(s15_m3_cyc_r), .QN(
        n17100) );
  AO221X1 U35496 ( .IN1(s7_msel_gnt_p3[2]), .IN2(n17008), .IN3(
        s7_msel_gnt_p2_2_), .IN4(n17009), .IN5(n17010), .Q(n14824) );
  AO22X1 U35497 ( .IN1(s7_msel_gnt_p0_2_), .IN2(n17011), .IN3(
        s7_msel_gnt_p1[2]), .IN4(n17012), .Q(n17010) );
  AO221X1 U35498 ( .IN1(test_so65), .IN2(n16999), .IN3(s6_msel_gnt_p2[2]), 
        .IN4(n17000), .IN5(n17001), .Q(n14819) );
  AO22X1 U35499 ( .IN1(s6_msel_gnt_p0[2]), .IN2(n17002), .IN3(test_so64), 
        .IN4(n17003), .Q(n17001) );
  AO221X1 U35500 ( .IN1(s14_msel_gnt_p3[2]), .IN2(n17072), .IN3(
        s14_msel_gnt_p2_2_), .IN4(n17073), .IN5(n17074), .Q(n14857) );
  AO22X1 U35501 ( .IN1(s14_msel_gnt_p0_2_), .IN2(n17075), .IN3(
        s14_msel_gnt_p1[2]), .IN4(n17076), .Q(n17074) );
  AO221X1 U35502 ( .IN1(s5_msel_gnt_p3_2_), .IN2(n17042), .IN3(
        s5_msel_gnt_p2[2]), .IN4(n17043), .IN5(n17044), .Q(n14842) );
  AO22X1 U35503 ( .IN1(s5_msel_gnt_p0[2]), .IN2(n17045), .IN3(
        s5_msel_gnt_p1_2_), .IN4(n17046), .Q(n17044) );
  AO221X1 U35504 ( .IN1(s4_msel_gnt_p3_2_), .IN2(n17034), .IN3(
        s4_msel_gnt_p2[2]), .IN4(n17035), .IN5(n17036), .Q(n14838) );
  AO22X1 U35505 ( .IN1(s4_msel_gnt_p0[2]), .IN2(n17037), .IN3(
        s4_msel_gnt_p1_2_), .IN4(n17038), .Q(n17036) );
  AO221X1 U35506 ( .IN1(s13_msel_gnt_p3[2]), .IN2(n17065), .IN3(
        s13_msel_gnt_p2_2_), .IN4(n17066), .IN5(n17067), .Q(n14854) );
  AO22X1 U35507 ( .IN1(s13_msel_gnt_p0_2_), .IN2(n17068), .IN3(
        s13_msel_gnt_p1[2]), .IN4(n17069), .Q(n17067) );
  AO221X1 U35508 ( .IN1(test_so88), .IN2(n17135), .IN3(s12_msel_gnt_p2[2]), 
        .IN4(n17136), .IN5(n17137), .Q(n14867) );
  AO22X1 U35509 ( .IN1(s12_msel_gnt_p0[2]), .IN2(n17138), .IN3(test_so87), 
        .IN4(n17139), .Q(n17137) );
  AO221X1 U35510 ( .IN1(s3_msel_gnt_p3[2]), .IN2(n17049), .IN3(test_so53), 
        .IN4(n17050), .IN5(n17051), .Q(n14845) );
  AO22X1 U35511 ( .IN1(test_so52), .IN2(n17052), .IN3(s3_msel_gnt_p1[2]), 
        .IN4(n17053), .Q(n17051) );
  AO221X1 U35512 ( .IN1(s2_msel_gnt_p3[2]), .IN2(n17057), .IN3(
        s2_msel_gnt_p2_2_), .IN4(n17058), .IN5(n17059), .Q(n14849) );
  AO22X1 U35513 ( .IN1(s2_msel_gnt_p0_2_), .IN2(n17060), .IN3(
        s2_msel_gnt_p1[2]), .IN4(n17061), .Q(n17059) );
  AO221X1 U35514 ( .IN1(s11_msel_gnt_p3_2_), .IN2(n17128), .IN3(
        s11_msel_gnt_p2[2]), .IN4(n17129), .IN5(n17130), .Q(n14864) );
  AO22X1 U35515 ( .IN1(s11_msel_gnt_p0[2]), .IN2(n17131), .IN3(
        s11_msel_gnt_p1_2_), .IN4(n17132), .Q(n17130) );
  AO221X1 U35516 ( .IN1(s10_msel_gnt_p3_2_), .IN2(n17142), .IN3(
        s10_msel_gnt_p2[2]), .IN4(n17143), .IN5(n17144), .Q(n14870) );
  AO22X1 U35517 ( .IN1(s10_msel_gnt_p0[2]), .IN2(n17145), .IN3(
        s10_msel_gnt_p1_2_), .IN4(n17146), .Q(n17144) );
  AO221X1 U35518 ( .IN1(s1_msel_gnt_p3[2]), .IN2(n17079), .IN3(
        s1_msel_gnt_p2_2_), .IN4(n17080), .IN5(n17081), .Q(n14860) );
  AO22X1 U35519 ( .IN1(s1_msel_gnt_p0_2_), .IN2(n17082), .IN3(
        s1_msel_gnt_p1[2]), .IN4(n17083), .Q(n17081) );
  AO221X1 U35520 ( .IN1(test_so42), .IN2(n17149), .IN3(s0_msel_gnt_p2[2]), 
        .IN4(n17150), .IN5(n17151), .Q(n14873) );
  AO22X1 U35521 ( .IN1(s0_msel_gnt_p0[2]), .IN2(n17152), .IN3(test_so41), 
        .IN4(n17153), .Q(n17151) );
  AO221X1 U35522 ( .IN1(s8_msel_gnt_p3[2]), .IN2(n17025), .IN3(
        s8_msel_gnt_p2_2_), .IN4(n17026), .IN5(n17027), .Q(n14833) );
  AO22X1 U35523 ( .IN1(s8_msel_gnt_p0_2_), .IN2(n17028), .IN3(
        s8_msel_gnt_p1[2]), .IN4(n17029), .Q(n17027) );
  AO221X1 U35524 ( .IN1(s9_msel_gnt_p3[2]), .IN2(n17016), .IN3(test_so76), 
        .IN4(n17017), .IN5(n17018), .Q(n14828) );
  AO22X1 U35525 ( .IN1(test_so75), .IN2(n17019), .IN3(s9_msel_gnt_p1[2]), 
        .IN4(n17020), .Q(n17018) );
  AO221X1 U35526 ( .IN1(s7_msel_gnt_p3[1]), .IN2(n17008), .IN3(
        s7_msel_gnt_p2_1_), .IN4(n17009), .IN5(n17014), .Q(n14823) );
  AO22X1 U35527 ( .IN1(s7_msel_gnt_p0_1_), .IN2(n17011), .IN3(
        s7_msel_gnt_p1[1]), .IN4(n17012), .Q(n17014) );
  AO221X1 U35528 ( .IN1(s6_msel_gnt_p3_1_), .IN2(n16999), .IN3(
        s6_msel_gnt_p2[1]), .IN4(n17000), .IN5(n17005), .Q(n14818) );
  AO22X1 U35529 ( .IN1(s6_msel_gnt_p0[1]), .IN2(n17002), .IN3(
        s6_msel_gnt_p1_1_), .IN4(n17003), .Q(n17005) );
  AO221X1 U35530 ( .IN1(s14_msel_gnt_p3[1]), .IN2(n17072), .IN3(test_so95), 
        .IN4(n17073), .IN5(n17078), .Q(n14856) );
  AO22X1 U35531 ( .IN1(test_so94), .IN2(n17075), .IN3(s14_msel_gnt_p1[1]), 
        .IN4(n17076), .Q(n17078) );
  AO221X1 U35532 ( .IN1(test_so61), .IN2(n17042), .IN3(s5_msel_gnt_p2[1]), 
        .IN4(n17043), .IN5(n17048), .Q(n14841) );
  AO22X1 U35533 ( .IN1(s5_msel_gnt_p0[1]), .IN2(n17045), .IN3(test_so60), 
        .IN4(n17046), .Q(n17048) );
  AO221X1 U35534 ( .IN1(s4_msel_gnt_p3_1_), .IN2(n17034), .IN3(
        s4_msel_gnt_p2[1]), .IN4(n17035), .IN5(n17040), .Q(n14837) );
  AO22X1 U35535 ( .IN1(s4_msel_gnt_p0[1]), .IN2(n17037), .IN3(
        s4_msel_gnt_p1_1_), .IN4(n17038), .Q(n17040) );
  AO221X1 U35536 ( .IN1(s13_msel_gnt_p3[1]), .IN2(n17065), .IN3(
        s13_msel_gnt_p2_1_), .IN4(n17066), .IN5(n17071), .Q(n14853) );
  AO22X1 U35537 ( .IN1(s13_msel_gnt_p0_1_), .IN2(n17068), .IN3(
        s13_msel_gnt_p1[1]), .IN4(n17069), .Q(n17071) );
  AO221X1 U35538 ( .IN1(s12_msel_gnt_p3_1_), .IN2(n17135), .IN3(
        s12_msel_gnt_p2[1]), .IN4(n17136), .IN5(n17141), .Q(n14866) );
  AO22X1 U35539 ( .IN1(s12_msel_gnt_p0[1]), .IN2(n17138), .IN3(
        s12_msel_gnt_p1_1_), .IN4(n17139), .Q(n17141) );
  AO221X1 U35540 ( .IN1(s3_msel_gnt_p3[1]), .IN2(n17049), .IN3(
        s3_msel_gnt_p2_1_), .IN4(n17050), .IN5(n17055), .Q(n14844) );
  AO22X1 U35541 ( .IN1(s3_msel_gnt_p0_1_), .IN2(n17052), .IN3(
        s3_msel_gnt_p1[1]), .IN4(n17053), .Q(n17055) );
  AO221X1 U35542 ( .IN1(s2_msel_gnt_p3[1]), .IN2(n17057), .IN3(test_so49), 
        .IN4(n17058), .IN5(n17063), .Q(n14848) );
  AO22X1 U35543 ( .IN1(test_so48), .IN2(n17060), .IN3(s2_msel_gnt_p1[1]), 
        .IN4(n17061), .Q(n17063) );
  AO221X1 U35544 ( .IN1(test_so84), .IN2(n17128), .IN3(s11_msel_gnt_p2[1]), 
        .IN4(n17129), .IN5(n17134), .Q(n14863) );
  AO22X1 U35545 ( .IN1(s11_msel_gnt_p0[1]), .IN2(n17131), .IN3(test_so83), 
        .IN4(n17132), .Q(n17134) );
  AO221X1 U35546 ( .IN1(s10_msel_gnt_p3_1_), .IN2(n17142), .IN3(
        s10_msel_gnt_p2[1]), .IN4(n17143), .IN5(n17148), .Q(n14869) );
  AO22X1 U35547 ( .IN1(s10_msel_gnt_p0[1]), .IN2(n17145), .IN3(
        s10_msel_gnt_p1_1_), .IN4(n17146), .Q(n17148) );
  AO221X1 U35548 ( .IN1(s1_msel_gnt_p3[1]), .IN2(n17079), .IN3(
        s1_msel_gnt_p2_1_), .IN4(n17080), .IN5(n17085), .Q(n14859) );
  AO22X1 U35549 ( .IN1(s1_msel_gnt_p0_1_), .IN2(n17082), .IN3(
        s1_msel_gnt_p1[1]), .IN4(n17083), .Q(n17085) );
  AO221X1 U35550 ( .IN1(s0_msel_gnt_p3_1_), .IN2(n17149), .IN3(
        s0_msel_gnt_p2[1]), .IN4(n17150), .IN5(n17155), .Q(n14872) );
  AO22X1 U35551 ( .IN1(s0_msel_gnt_p0[1]), .IN2(n17152), .IN3(
        s0_msel_gnt_p1_1_), .IN4(n17153), .Q(n17155) );
  AO221X1 U35552 ( .IN1(s8_msel_gnt_p3[1]), .IN2(n17025), .IN3(test_so72), 
        .IN4(n17026), .IN5(n17031), .Q(n14832) );
  AO22X1 U35553 ( .IN1(test_so71), .IN2(n17028), .IN3(s8_msel_gnt_p1[1]), 
        .IN4(n17029), .Q(n17031) );
  AO221X1 U35554 ( .IN1(s9_msel_gnt_p3[1]), .IN2(n17016), .IN3(
        s9_msel_gnt_p2_1_), .IN4(n17017), .IN5(n17022), .Q(n14827) );
  AO22X1 U35555 ( .IN1(s9_msel_gnt_p0_1_), .IN2(n17019), .IN3(
        s9_msel_gnt_p1[1]), .IN4(n17020), .Q(n17022) );
  AO221X1 U35556 ( .IN1(s7_msel_gnt_p3[0]), .IN2(n17008), .IN3(test_so68), 
        .IN4(n17009), .IN5(n17013), .Q(n14825) );
  AO22X1 U35557 ( .IN1(test_so67), .IN2(n17011), .IN3(s7_msel_gnt_p1[0]), 
        .IN4(n17012), .Q(n17013) );
  AO221X1 U35558 ( .IN1(s6_msel_gnt_p3_0_), .IN2(n16999), .IN3(
        s6_msel_gnt_p2[0]), .IN4(n17000), .IN5(n17004), .Q(n14820) );
  AO22X1 U35559 ( .IN1(s6_msel_gnt_p0[0]), .IN2(n17002), .IN3(
        s6_msel_gnt_p1_0_), .IN4(n17003), .Q(n17004) );
  AO221X1 U35560 ( .IN1(s14_msel_gnt_p3[0]), .IN2(n17072), .IN3(
        s14_msel_gnt_p2_0_), .IN4(n17073), .IN5(n17077), .Q(n14858) );
  AO22X1 U35561 ( .IN1(s14_msel_gnt_p0_0_), .IN2(n17075), .IN3(
        s14_msel_gnt_p1[0]), .IN4(n17076), .Q(n17077) );
  AO221X1 U35562 ( .IN1(s5_msel_gnt_p3_0_), .IN2(n17042), .IN3(
        s5_msel_gnt_p2[0]), .IN4(n17043), .IN5(n17047), .Q(n14843) );
  AO22X1 U35563 ( .IN1(s5_msel_gnt_p0[0]), .IN2(n17045), .IN3(
        s5_msel_gnt_p1_0_), .IN4(n17046), .Q(n17047) );
  AO221X1 U35564 ( .IN1(test_so57), .IN2(n17034), .IN3(s4_msel_gnt_p2[0]), 
        .IN4(n17035), .IN5(n17039), .Q(n14839) );
  AO22X1 U35565 ( .IN1(s4_msel_gnt_p0[0]), .IN2(n17037), .IN3(test_so56), 
        .IN4(n17038), .Q(n17039) );
  AO221X1 U35566 ( .IN1(s13_msel_gnt_p3[0]), .IN2(n17065), .IN3(test_so91), 
        .IN4(n17066), .IN5(n17070), .Q(n14855) );
  AO22X1 U35567 ( .IN1(test_so90), .IN2(n17068), .IN3(s13_msel_gnt_p1[0]), 
        .IN4(n17069), .Q(n17070) );
  AO221X1 U35568 ( .IN1(s12_msel_gnt_p3_0_), .IN2(n17135), .IN3(
        s12_msel_gnt_p2[0]), .IN4(n17136), .IN5(n17140), .Q(n14868) );
  AO22X1 U35569 ( .IN1(s12_msel_gnt_p0[0]), .IN2(n17138), .IN3(
        s12_msel_gnt_p1_0_), .IN4(n17139), .Q(n17140) );
  AO221X1 U35570 ( .IN1(s3_msel_gnt_p3[0]), .IN2(n17049), .IN3(
        s3_msel_gnt_p2_0_), .IN4(n17050), .IN5(n17054), .Q(n14846) );
  AO22X1 U35571 ( .IN1(s3_msel_gnt_p0_0_), .IN2(n17052), .IN3(
        s3_msel_gnt_p1[0]), .IN4(n17053), .Q(n17054) );
  AO221X1 U35572 ( .IN1(s2_msel_gnt_p3[0]), .IN2(n17057), .IN3(
        s2_msel_gnt_p2_0_), .IN4(n17058), .IN5(n17062), .Q(n14850) );
  AO22X1 U35573 ( .IN1(s2_msel_gnt_p0_0_), .IN2(n17060), .IN3(
        s2_msel_gnt_p1[0]), .IN4(n17061), .Q(n17062) );
  AO221X1 U35574 ( .IN1(s11_msel_gnt_p3_0_), .IN2(n17128), .IN3(
        s11_msel_gnt_p2[0]), .IN4(n17129), .IN5(n17133), .Q(n14865) );
  AO22X1 U35575 ( .IN1(s11_msel_gnt_p0[0]), .IN2(n17131), .IN3(
        s11_msel_gnt_p1_0_), .IN4(n17132), .Q(n17133) );
  AO221X1 U35576 ( .IN1(test_so80), .IN2(n17142), .IN3(s10_msel_gnt_p2[0]), 
        .IN4(n17143), .IN5(n17147), .Q(n14871) );
  AO22X1 U35577 ( .IN1(s10_msel_gnt_p0[0]), .IN2(n17145), .IN3(test_so79), 
        .IN4(n17146), .Q(n17147) );
  AO221X1 U35578 ( .IN1(s1_msel_gnt_p3[0]), .IN2(n17079), .IN3(test_so45), 
        .IN4(n17080), .IN5(n17084), .Q(n14861) );
  AO22X1 U35579 ( .IN1(test_so44), .IN2(n17082), .IN3(s1_msel_gnt_p1[0]), 
        .IN4(n17083), .Q(n17084) );
  AO221X1 U35580 ( .IN1(s0_msel_gnt_p3_0_), .IN2(n17149), .IN3(
        s0_msel_gnt_p2[0]), .IN4(n17150), .IN5(n17154), .Q(n14874) );
  AO22X1 U35581 ( .IN1(s0_msel_gnt_p0[0]), .IN2(n17152), .IN3(
        s0_msel_gnt_p1_0_), .IN4(n17153), .Q(n17154) );
  AO221X1 U35582 ( .IN1(s9_msel_gnt_p3[0]), .IN2(n17016), .IN3(
        s9_msel_gnt_p2_0_), .IN4(n17017), .IN5(n17021), .Q(n14829) );
  AO22X1 U35583 ( .IN1(s9_msel_gnt_p0_0_), .IN2(n17019), .IN3(
        s9_msel_gnt_p1[0]), .IN4(n17020), .Q(n17021) );
  AO221X1 U35584 ( .IN1(s8_msel_gnt_p3[0]), .IN2(n17025), .IN3(
        s8_msel_gnt_p2_0_), .IN4(n17026), .IN5(n17030), .Q(n14834) );
  AO22X1 U35585 ( .IN1(s8_msel_gnt_p0_0_), .IN2(n17028), .IN3(
        s8_msel_gnt_p1[0]), .IN4(n17029), .Q(n17030) );
  NOR2X0 U35586 ( .IN1(m7_addr_i[30]), .IN2(m7_addr_i[29]), .QN(n14830) );
  NOR2X0 U35587 ( .IN1(m6_addr_i[30]), .IN2(m6_addr_i[29]), .QN(n15172) );
  NOR2X0 U35588 ( .IN1(m5_addr_i[30]), .IN2(m5_addr_i[29]), .QN(n15477) );
  NOR2X0 U35589 ( .IN1(m4_addr_i[30]), .IN2(m4_addr_i[29]), .QN(n15782) );
  NOR2X0 U35590 ( .IN1(m3_addr_i[30]), .IN2(m3_addr_i[29]), .QN(n16087) );
  NOR2X0 U35591 ( .IN1(m2_addr_i[30]), .IN2(m2_addr_i[29]), .QN(n16392) );
  NOR2X0 U35592 ( .IN1(m1_addr_i[30]), .IN2(m1_addr_i[29]), .QN(n16697) );
  NOR2X0 U35593 ( .IN1(m0_addr_i[30]), .IN2(m0_addr_i[29]), .QN(n17023) );
  NOR2X0 U35594 ( .IN1(m7_addr_i[31]), .IN2(m7_addr_i[28]), .QN(n14821) );
  NOR2X0 U35595 ( .IN1(m6_addr_i[31]), .IN2(m6_addr_i[28]), .QN(n15169) );
  NOR2X0 U35596 ( .IN1(m5_addr_i[31]), .IN2(m5_addr_i[28]), .QN(n15474) );
  NOR2X0 U35597 ( .IN1(m4_addr_i[31]), .IN2(m4_addr_i[28]), .QN(n15779) );
  NOR2X0 U35598 ( .IN1(m3_addr_i[31]), .IN2(m3_addr_i[28]), .QN(n16084) );
  NOR2X0 U35599 ( .IN1(m2_addr_i[31]), .IN2(m2_addr_i[28]), .QN(n16389) );
  NOR2X0 U35600 ( .IN1(m1_addr_i[31]), .IN2(m1_addr_i[28]), .QN(n16694) );
  NOR2X0 U35601 ( .IN1(m0_addr_i[31]), .IN2(m0_addr_i[28]), .QN(n17006) );
  NOR2X0 U35602 ( .IN1(n2274), .IN2(m7_addr_i[28]), .QN(n14835) );
  NOR2X0 U35603 ( .IN1(n2102), .IN2(m5_addr_i[28]), .QN(n15479) );
  NOR2X0 U35604 ( .IN1(n1930), .IN2(m3_addr_i[28]), .QN(n16089) );
  NOR2X0 U35605 ( .IN1(n1758), .IN2(m1_addr_i[28]), .QN(n16699) );
  NOR2X0 U35606 ( .IN1(n2188), .IN2(m6_addr_i[28]), .QN(n15174) );
  NOR2X0 U35607 ( .IN1(n2016), .IN2(m4_addr_i[28]), .QN(n15784) );
  NOR2X0 U35608 ( .IN1(n1844), .IN2(m2_addr_i[28]), .QN(n16394) );
  NOR2X0 U35609 ( .IN1(n1650), .IN2(m0_addr_i[28]), .QN(n17032) );
  NOR2X0 U35610 ( .IN1(n2277), .IN2(m7_addr_i[31]), .QN(n14826) );
  NOR2X0 U35611 ( .IN1(n2105), .IN2(m5_addr_i[31]), .QN(n15476) );
  NOR2X0 U35612 ( .IN1(n1933), .IN2(m3_addr_i[31]), .QN(n16086) );
  NOR2X0 U35613 ( .IN1(n1761), .IN2(m1_addr_i[31]), .QN(n16696) );
  NOR2X0 U35614 ( .IN1(n2191), .IN2(m6_addr_i[31]), .QN(n15171) );
  NOR2X0 U35615 ( .IN1(n2019), .IN2(m4_addr_i[31]), .QN(n15781) );
  NOR2X0 U35616 ( .IN1(n1847), .IN2(m2_addr_i[31]), .QN(n16391) );
  NOR2X0 U35617 ( .IN1(n1657), .IN2(m0_addr_i[31]), .QN(n17015) );
  NOR2X0 U35618 ( .IN1(n2276), .IN2(m7_addr_i[30]), .QN(n14847) );
  NOR2X0 U35619 ( .IN1(n2104), .IN2(m5_addr_i[30]), .QN(n15482) );
  NOR2X0 U35620 ( .IN1(n1932), .IN2(m3_addr_i[30]), .QN(n16092) );
  NOR2X0 U35621 ( .IN1(n1760), .IN2(m1_addr_i[30]), .QN(n16702) );
  NOR2X0 U35622 ( .IN1(n2275), .IN2(m7_addr_i[29]), .QN(n14840) );
  NOR2X0 U35623 ( .IN1(n2103), .IN2(m5_addr_i[29]), .QN(n15481) );
  NOR2X0 U35624 ( .IN1(n1931), .IN2(m3_addr_i[29]), .QN(n16091) );
  NOR2X0 U35625 ( .IN1(n1759), .IN2(m1_addr_i[29]), .QN(n16701) );
  NOR2X0 U35626 ( .IN1(n2190), .IN2(m6_addr_i[30]), .QN(n15177) );
  NOR2X0 U35627 ( .IN1(n2018), .IN2(m4_addr_i[30]), .QN(n15787) );
  NOR2X0 U35628 ( .IN1(n1846), .IN2(m2_addr_i[30]), .QN(n16397) );
  NOR2X0 U35629 ( .IN1(n1656), .IN2(m0_addr_i[30]), .QN(n17056) );
  NOR2X0 U35630 ( .IN1(n2189), .IN2(m6_addr_i[29]), .QN(n15176) );
  NOR2X0 U35631 ( .IN1(n2017), .IN2(m4_addr_i[29]), .QN(n15786) );
  NOR2X0 U35632 ( .IN1(n1845), .IN2(m2_addr_i[29]), .QN(n16396) );
  NOR2X0 U35633 ( .IN1(n1655), .IN2(m0_addr_i[29]), .QN(n17041) );
  ISOLANDX1 U35634 ( .D(m6s7_cyc), .ISO(n13662), .Q(n13677) );
  ISOLANDX1 U35635 ( .D(m6s6_cyc), .ISO(n13353), .Q(n13368) );
  ISOLANDX1 U35636 ( .D(m6s14_cyc), .ISO(n11187), .Q(n11202) );
  ISOLANDX1 U35637 ( .D(m6s5_cyc), .ISO(n13044), .Q(n13059) );
  ISOLANDX1 U35638 ( .D(m6s4_cyc), .ISO(n12735), .Q(n12750) );
  ISOLANDX1 U35639 ( .D(m6s13_cyc), .ISO(n10878), .Q(n10893) );
  ISOLANDX1 U35640 ( .D(m6s12_cyc), .ISO(n10568), .Q(n10583) );
  ISOLANDX1 U35641 ( .D(test_so31), .ISO(n12426), .Q(n12441) );
  ISOLANDX1 U35642 ( .D(m6s2_cyc), .ISO(n12117), .Q(n12132) );
  ISOLANDX1 U35643 ( .D(m6s11_cyc), .ISO(n10259), .Q(n10274) );
  ISOLANDX1 U35644 ( .D(m6s10_cyc), .ISO(n9949), .Q(n9964) );
  ISOLANDX1 U35645 ( .D(m6s1_cyc), .ISO(n11807), .Q(n11822) );
  ISOLANDX1 U35646 ( .D(m6s0_cyc), .ISO(n11497), .Q(n11512) );
  ISOLANDX1 U35647 ( .D(test_so32), .ISO(n9639), .Q(n9654) );
  ISOLANDX1 U35648 ( .D(m6s8_cyc), .ISO(n9328), .Q(n9343) );
  INVX0 U35649 ( .IN(m7_addr_i[2]), .QN(n2303) );
  INVX0 U35650 ( .IN(m5_addr_i[2]), .QN(n2131) );
  INVX0 U35651 ( .IN(m3_addr_i[2]), .QN(n1959) );
  INVX0 U35652 ( .IN(m1_addr_i[2]), .QN(n1787) );
  INVX0 U35653 ( .IN(m7_addr_i[3]), .QN(n2302) );
  INVX0 U35654 ( .IN(m5_addr_i[3]), .QN(n2130) );
  INVX0 U35655 ( .IN(m3_addr_i[3]), .QN(n1958) );
  INVX0 U35656 ( .IN(m1_addr_i[3]), .QN(n1786) );
  INVX0 U35657 ( .IN(m7_addr_i[4]), .QN(n2301) );
  INVX0 U35658 ( .IN(m5_addr_i[4]), .QN(n2129) );
  INVX0 U35659 ( .IN(m3_addr_i[4]), .QN(n1957) );
  INVX0 U35660 ( .IN(m1_addr_i[4]), .QN(n1785) );
  INVX0 U35661 ( .IN(m7_addr_i[5]), .QN(n2300) );
  INVX0 U35662 ( .IN(m5_addr_i[5]), .QN(n2128) );
  INVX0 U35663 ( .IN(m3_addr_i[5]), .QN(n1956) );
  INVX0 U35664 ( .IN(m1_addr_i[5]), .QN(n1784) );
  INVX0 U35665 ( .IN(m6_addr_i[2]), .QN(n2217) );
  INVX0 U35666 ( .IN(m4_addr_i[2]), .QN(n2045) );
  INVX0 U35667 ( .IN(m2_addr_i[2]), .QN(n1873) );
  INVX0 U35668 ( .IN(m0_addr_i[2]), .QN(n1701) );
  INVX0 U35669 ( .IN(m6_addr_i[3]), .QN(n2216) );
  INVX0 U35670 ( .IN(m4_addr_i[3]), .QN(n2044) );
  INVX0 U35671 ( .IN(m2_addr_i[3]), .QN(n1872) );
  INVX0 U35672 ( .IN(m0_addr_i[3]), .QN(n1699) );
  INVX0 U35673 ( .IN(m6_addr_i[4]), .QN(n2215) );
  INVX0 U35674 ( .IN(m4_addr_i[4]), .QN(n2043) );
  INVX0 U35675 ( .IN(m2_addr_i[4]), .QN(n1871) );
  INVX0 U35676 ( .IN(m0_addr_i[4]), .QN(n1697) );
  INVX0 U35677 ( .IN(m6_addr_i[5]), .QN(n2214) );
  INVX0 U35678 ( .IN(m4_addr_i[5]), .QN(n2042) );
  INVX0 U35679 ( .IN(m2_addr_i[5]), .QN(n1870) );
  INVX0 U35680 ( .IN(m0_addr_i[5]), .QN(n1696) );
  NOR2X0 U35681 ( .IN1(n21016), .IN2(s7_next), .QN(n13627) );
  NOR2X0 U35682 ( .IN1(n21015), .IN2(s6_next), .QN(n13318) );
  NOR2X0 U35683 ( .IN1(n21008), .IN2(s14_next), .QN(n11152) );
  NOR2X0 U35684 ( .IN1(n21014), .IN2(s5_next), .QN(n13009) );
  NOR2X0 U35685 ( .IN1(n21013), .IN2(s4_next), .QN(n12700) );
  NOR2X0 U35686 ( .IN1(n21007), .IN2(s13_next), .QN(n10843) );
  NOR2X0 U35687 ( .IN1(n21006), .IN2(s12_next), .QN(n10533) );
  NOR2X0 U35688 ( .IN1(n21012), .IN2(test_so54), .QN(n12391) );
  NOR2X0 U35689 ( .IN1(n21011), .IN2(s2_next), .QN(n12082) );
  NOR2X0 U35690 ( .IN1(n21005), .IN2(s11_next), .QN(n10224) );
  NOR2X0 U35691 ( .IN1(n21004), .IN2(s10_next), .QN(n9914) );
  NOR2X0 U35692 ( .IN1(n21010), .IN2(s1_next), .QN(n11772) );
  NOR2X0 U35693 ( .IN1(n21009), .IN2(s0_next), .QN(n11462) );
  NOR2X0 U35694 ( .IN1(n21003), .IN2(test_so77), .QN(n9604) );
  NOR2X0 U35695 ( .IN1(n21002), .IN2(s8_next), .QN(n9293) );
  NOR2X0 U35696 ( .IN1(n21017), .IN2(test_so100), .QN(n14270) );
  NOR2X0 U35697 ( .IN1(n3853), .IN2(test_so69), .QN(n17009) );
  NOR2X0 U35698 ( .IN1(n3808), .IN2(s6_msel_pri_out_0_), .QN(n17000) );
  NOR2X0 U35699 ( .IN1(n4168), .IN2(s14_msel_pri_out_0_), .QN(n17073) );
  NOR2X0 U35700 ( .IN1(n3763), .IN2(s5_msel_pri_out_0_), .QN(n17043) );
  NOR2X0 U35701 ( .IN1(n3718), .IN2(s4_msel_pri_out_0_), .QN(n17035) );
  NOR2X0 U35702 ( .IN1(n4123), .IN2(test_so92), .QN(n17066) );
  NOR2X0 U35703 ( .IN1(n4078), .IN2(s12_msel_pri_out_0_), .QN(n17136) );
  NOR2X0 U35704 ( .IN1(n3673), .IN2(s3_msel_pri_out_0_), .QN(n17050) );
  NOR2X0 U35705 ( .IN1(n3628), .IN2(s2_msel_pri_out_0_), .QN(n17058) );
  NOR2X0 U35706 ( .IN1(n4033), .IN2(s11_msel_pri_out_0_), .QN(n17129) );
  NOR2X0 U35707 ( .IN1(n3988), .IN2(s10_msel_pri_out_0_), .QN(n17143) );
  NOR2X0 U35708 ( .IN1(n3583), .IN2(test_so46), .QN(n17080) );
  NOR2X0 U35709 ( .IN1(n3538), .IN2(s0_msel_pri_out_0_), .QN(n17150) );
  NOR2X0 U35710 ( .IN1(n3898), .IN2(s8_msel_pri_out_0_), .QN(n17026) );
  NOR2X0 U35711 ( .IN1(n3943), .IN2(s9_msel_pri_out_0_), .QN(n17017) );
  NOR2X0 U35712 ( .IN1(n3853), .IN2(n3852), .QN(n17008) );
  NOR2X0 U35713 ( .IN1(n3808), .IN2(n3807), .QN(n16999) );
  NOR2X0 U35714 ( .IN1(n4168), .IN2(n4167), .QN(n17072) );
  NOR2X0 U35715 ( .IN1(n3763), .IN2(n3762), .QN(n17042) );
  NOR2X0 U35716 ( .IN1(n3718), .IN2(n3717), .QN(n17034) );
  NOR2X0 U35717 ( .IN1(n4123), .IN2(n4122), .QN(n17065) );
  NOR2X0 U35718 ( .IN1(n4078), .IN2(n4077), .QN(n17135) );
  NOR2X0 U35719 ( .IN1(n3673), .IN2(n3672), .QN(n17049) );
  NOR2X0 U35720 ( .IN1(n3628), .IN2(n3627), .QN(n17057) );
  NOR2X0 U35721 ( .IN1(n4033), .IN2(n4032), .QN(n17128) );
  NOR2X0 U35722 ( .IN1(n3988), .IN2(n3987), .QN(n17142) );
  NOR2X0 U35723 ( .IN1(n3583), .IN2(n3582), .QN(n17079) );
  NOR2X0 U35724 ( .IN1(n3538), .IN2(n3537), .QN(n17149) );
  NOR2X0 U35725 ( .IN1(n3898), .IN2(n3897), .QN(n17025) );
  NOR2X0 U35726 ( .IN1(n3943), .IN2(n3942), .QN(n17016) );
  NOR2X0 U35727 ( .IN1(test_so69), .IN2(s7_msel_pri_out_1_), .QN(n17011) );
  NOR2X0 U35728 ( .IN1(s6_msel_pri_out_0_), .IN2(s6_msel_pri_out_1_), .QN(
        n17002) );
  NOR2X0 U35729 ( .IN1(s14_msel_pri_out_0_), .IN2(test_so96), .QN(n17075) );
  NOR2X0 U35730 ( .IN1(s5_msel_pri_out_0_), .IN2(s5_msel_pri_out_1_), .QN(
        n17045) );
  NOR2X0 U35731 ( .IN1(s4_msel_pri_out_0_), .IN2(s4_msel_pri_out_1_), .QN(
        n17037) );
  NOR2X0 U35732 ( .IN1(test_so92), .IN2(s13_msel_pri_out_1_), .QN(n17068) );
  NOR2X0 U35733 ( .IN1(s12_msel_pri_out_0_), .IN2(s12_msel_pri_out_1_), .QN(
        n17138) );
  NOR2X0 U35734 ( .IN1(s3_msel_pri_out_0_), .IN2(s3_msel_pri_out_1_), .QN(
        n17052) );
  NOR2X0 U35735 ( .IN1(s2_msel_pri_out_0_), .IN2(test_so50), .QN(n17060) );
  NOR2X0 U35736 ( .IN1(s11_msel_pri_out_0_), .IN2(s11_msel_pri_out_1_), .QN(
        n17131) );
  NOR2X0 U35737 ( .IN1(s10_msel_pri_out_0_), .IN2(s10_msel_pri_out_1_), .QN(
        n17145) );
  NOR2X0 U35738 ( .IN1(test_so46), .IN2(s1_msel_pri_out_1_), .QN(n17082) );
  NOR2X0 U35739 ( .IN1(s0_msel_pri_out_0_), .IN2(s0_msel_pri_out_1_), .QN(
        n17152) );
  NOR2X0 U35740 ( .IN1(s8_msel_pri_out_0_), .IN2(test_so73), .QN(n17028) );
  NOR2X0 U35741 ( .IN1(s9_msel_pri_out_0_), .IN2(s9_msel_pri_out_1_), .QN(
        n17019) );
  INVX0 U35742 ( .IN(rst_i), .QN(n21089) );
  INVX0 U35743 ( .IN(rst_i), .QN(n21088) );
  NOR2X0 U35744 ( .IN1(n3852), .IN2(s7_msel_pri_out_1_), .QN(n17012) );
  NOR2X0 U35745 ( .IN1(n3807), .IN2(s6_msel_pri_out_1_), .QN(n17003) );
  NOR2X0 U35746 ( .IN1(n4167), .IN2(test_so96), .QN(n17076) );
  NOR2X0 U35747 ( .IN1(n3762), .IN2(s5_msel_pri_out_1_), .QN(n17046) );
  NOR2X0 U35748 ( .IN1(n3717), .IN2(s4_msel_pri_out_1_), .QN(n17038) );
  NOR2X0 U35749 ( .IN1(n4122), .IN2(s13_msel_pri_out_1_), .QN(n17069) );
  NOR2X0 U35750 ( .IN1(n4077), .IN2(s12_msel_pri_out_1_), .QN(n17139) );
  NOR2X0 U35751 ( .IN1(n3672), .IN2(s3_msel_pri_out_1_), .QN(n17053) );
  NOR2X0 U35752 ( .IN1(n3627), .IN2(test_so50), .QN(n17061) );
  NOR2X0 U35753 ( .IN1(n4032), .IN2(s11_msel_pri_out_1_), .QN(n17132) );
  NOR2X0 U35754 ( .IN1(n3987), .IN2(s10_msel_pri_out_1_), .QN(n17146) );
  NOR2X0 U35755 ( .IN1(n3582), .IN2(s1_msel_pri_out_1_), .QN(n17083) );
  NOR2X0 U35756 ( .IN1(n3537), .IN2(s0_msel_pri_out_1_), .QN(n17153) );
  NOR2X0 U35757 ( .IN1(n3897), .IN2(test_so73), .QN(n17029) );
  NOR2X0 U35758 ( .IN1(n3942), .IN2(s9_msel_pri_out_1_), .QN(n17020) );
  NAND2X0 U35759 ( .IN1(conf7_13_), .IN2(n18029), .QN(n13662) );
  NAND2X0 U35760 ( .IN1(conf6_13_), .IN2(n18197), .QN(n13353) );
  NAND2X0 U35761 ( .IN1(conf14_13_), .IN2(n18198), .QN(n11187) );
  NAND2X0 U35762 ( .IN1(conf5_13_), .IN2(n18045), .QN(n13044) );
  NAND2X0 U35763 ( .IN1(conf4_13_), .IN2(n18213), .QN(n12735) );
  NAND2X0 U35764 ( .IN1(conf13_13_), .IN2(n18046), .QN(n10878) );
  NAND2X0 U35765 ( .IN1(conf12_13_), .IN2(n18214), .QN(n10568) );
  NAND2X0 U35766 ( .IN1(conf3_13_), .IN2(n18030), .QN(n12426) );
  NAND2X0 U35767 ( .IN1(conf2_13_), .IN2(n18199), .QN(n12117) );
  NAND2X0 U35768 ( .IN1(conf11_13_), .IN2(n18047), .QN(n10259) );
  NAND2X0 U35769 ( .IN1(conf10_13_), .IN2(n18215), .QN(n9949) );
  NAND2X0 U35770 ( .IN1(conf1_13_), .IN2(n18048), .QN(n11807) );
  NAND2X0 U35771 ( .IN1(conf0_13_), .IN2(n18216), .QN(n11497) );
  NAND2X0 U35772 ( .IN1(conf9_13_), .IN2(n18031), .QN(n9639) );
  NAND2X0 U35773 ( .IN1(conf8_13_), .IN2(n18200), .QN(n9328) );
  NAND2X0 U35774 ( .IN1(conf15_9_), .IN2(n18150), .QN(n14301) );
  NAND3X0 U35775 ( .IN1(m7s7_cyc), .IN2(n20666), .IN3(s7_m7_cyc_r), .QN(n14419) );
  NAND3X0 U35776 ( .IN1(test_so24), .IN2(n20600), .IN3(s7_m3_cyc_r), .QN(
        n14415) );
  NAND3X0 U35777 ( .IN1(m7s6_cyc), .IN2(n20534), .IN3(test_so63), .QN(n14429)
         );
  NAND3X0 U35778 ( .IN1(m3s6_cyc), .IN2(n20468), .IN3(s6_m3_cyc_r), .QN(n14425) );
  NAND3X0 U35779 ( .IN1(m7s14_cyc), .IN2(n19612), .IN3(s14_m7_cyc_r), .QN(
        n14349) );
  NAND3X0 U35780 ( .IN1(test_so25), .IN2(n19546), .IN3(test_so93), .QN(n14345)
         );
  NAND3X0 U35781 ( .IN1(test_so34), .IN2(n20402), .IN3(s5_m7_cyc_r), .QN(
        n14439) );
  NAND3X0 U35782 ( .IN1(m3s5_cyc), .IN2(n20336), .IN3(s5_m3_cyc_r), .QN(n14435) );
  NAND3X0 U35783 ( .IN1(m7s4_cyc), .IN2(n20270), .IN3(s4_m7_cyc_r), .QN(n14449) );
  NAND3X0 U35784 ( .IN1(m3s4_cyc), .IN2(n20204), .IN3(s4_m3_cyc_r), .QN(n14445) );
  NAND3X0 U35785 ( .IN1(m7s13_cyc), .IN2(n19480), .IN3(s13_m7_cyc_r), .QN(
        n14359) );
  NAND3X0 U35786 ( .IN1(m3s13_cyc), .IN2(n19414), .IN3(s13_m3_cyc_r), .QN(
        n14355) );
  NAND3X0 U35787 ( .IN1(m7s12_cyc), .IN2(n19348), .IN3(test_so86), .QN(n14369)
         );
  NAND3X0 U35788 ( .IN1(m3s12_cyc), .IN2(n19282), .IN3(s12_m3_cyc_r), .QN(
        n14365) );
  NAND3X0 U35789 ( .IN1(m7s3_cyc), .IN2(n20138), .IN3(s3_m7_cyc_r), .QN(n14459) );
  NAND3X0 U35790 ( .IN1(m3s3_cyc), .IN2(n20073), .IN3(s3_m3_cyc_r), .QN(n14455) );
  NAND3X0 U35791 ( .IN1(m7s2_cyc), .IN2(n20007), .IN3(s2_m7_cyc_r), .QN(n14469) );
  NAND3X0 U35792 ( .IN1(m3s2_cyc), .IN2(n19942), .IN3(test_so47), .QN(n14465)
         );
  NAND3X0 U35793 ( .IN1(test_so35), .IN2(n19216), .IN3(s11_m7_cyc_r), .QN(
        n14379) );
  NAND3X0 U35794 ( .IN1(m3s11_cyc), .IN2(n19150), .IN3(s11_m3_cyc_r), .QN(
        n14375) );
  NAND3X0 U35795 ( .IN1(m7s10_cyc), .IN2(n19084), .IN3(s10_m7_cyc_r), .QN(
        n14389) );
  NAND3X0 U35796 ( .IN1(m3s10_cyc), .IN2(n19018), .IN3(s10_m3_cyc_r), .QN(
        n14385) );
  NAND3X0 U35797 ( .IN1(m7s1_cyc), .IN2(n19876), .IN3(s1_m7_cyc_r), .QN(n14479) );
  NAND3X0 U35798 ( .IN1(m3s1_cyc), .IN2(n19810), .IN3(s1_m3_cyc_r), .QN(n14475) );
  NAND3X0 U35799 ( .IN1(m7s0_cyc), .IN2(n18952), .IN3(test_so40), .QN(n14489)
         );
  NAND3X0 U35800 ( .IN1(test_so23), .IN2(n18886), .IN3(s0_m3_cyc_r), .QN(
        n14485) );
  NAND3X0 U35801 ( .IN1(m7s9_cyc), .IN2(n20870), .IN3(s9_m7_cyc_r), .QN(n14399) );
  NAND3X0 U35802 ( .IN1(m3s9_cyc), .IN2(n20834), .IN3(s9_m3_cyc_r), .QN(n14395) );
  NAND3X0 U35803 ( .IN1(m7s8_cyc), .IN2(n20798), .IN3(s8_m7_cyc_r), .QN(n14409) );
  NAND3X0 U35804 ( .IN1(m3s8_cyc), .IN2(n20732), .IN3(test_so70), .QN(n14405)
         );
  NAND3X0 U35805 ( .IN1(m6s7_cyc), .IN2(n20657), .IN3(s7_m6_cyc_r), .QN(n14418) );
  NAND3X0 U35806 ( .IN1(m2s7_cyc), .IN2(n20591), .IN3(test_so66), .QN(n14414)
         );
  NAND3X0 U35807 ( .IN1(m6s6_cyc), .IN2(n20525), .IN3(s6_m6_cyc_r), .QN(n14428) );
  NAND3X0 U35808 ( .IN1(m2s6_cyc), .IN2(n20459), .IN3(s6_m2_cyc_r), .QN(n14424) );
  NAND3X0 U35809 ( .IN1(m6s14_cyc), .IN2(n19603), .IN3(s14_m6_cyc_r), .QN(
        n14348) );
  NAND3X0 U35810 ( .IN1(m2s14_cyc), .IN2(n19537), .IN3(s14_m2_cyc_r), .QN(
        n14344) );
  NAND3X0 U35811 ( .IN1(m6s5_cyc), .IN2(n20393), .IN3(test_so59), .QN(n14438)
         );
  NAND3X0 U35812 ( .IN1(m2s5_cyc), .IN2(n20327), .IN3(s5_m2_cyc_r), .QN(n14434) );
  NAND3X0 U35813 ( .IN1(m6s4_cyc), .IN2(n20261), .IN3(s4_m6_cyc_r), .QN(n14448) );
  NAND3X0 U35814 ( .IN1(m2s4_cyc), .IN2(n20195), .IN3(s4_m2_cyc_r), .QN(n14444) );
  NAND3X0 U35815 ( .IN1(m6s13_cyc), .IN2(n19471), .IN3(s13_m6_cyc_r), .QN(
        n14358) );
  NAND3X0 U35816 ( .IN1(m2s13_cyc), .IN2(n19405), .IN3(test_so89), .QN(n14354)
         );
  NAND3X0 U35817 ( .IN1(m6s12_cyc), .IN2(n19339), .IN3(s12_m6_cyc_r), .QN(
        n14368) );
  NAND3X0 U35818 ( .IN1(m2s12_cyc), .IN2(n19273), .IN3(s12_m2_cyc_r), .QN(
        n14364) );
  NAND3X0 U35819 ( .IN1(test_so31), .IN2(n20129), .IN3(s3_m6_cyc_r), .QN(
        n14458) );
  NAND3X0 U35820 ( .IN1(m2s3_cyc), .IN2(n17915), .IN3(s3_m2_cyc_r), .QN(n14454) );
  NAND3X0 U35821 ( .IN1(m6s2_cyc), .IN2(n19998), .IN3(s2_m6_cyc_r), .QN(n14468) );
  NAND3X0 U35822 ( .IN1(test_so21), .IN2(n17916), .IN3(s2_m2_cyc_r), .QN(
        n14464) );
  NAND3X0 U35823 ( .IN1(m6s11_cyc), .IN2(n19207), .IN3(test_so82), .QN(n14378)
         );
  NAND3X0 U35824 ( .IN1(m2s11_cyc), .IN2(n19141), .IN3(s11_m2_cyc_r), .QN(
        n14374) );
  NAND3X0 U35825 ( .IN1(m6s10_cyc), .IN2(n19075), .IN3(s10_m6_cyc_r), .QN(
        n14388) );
  NAND3X0 U35826 ( .IN1(m2s10_cyc), .IN2(n17906), .IN3(s10_m2_cyc_r), .QN(
        n14384) );
  NAND3X0 U35827 ( .IN1(m6s1_cyc), .IN2(n19867), .IN3(s1_m6_cyc_r), .QN(n14478) );
  NAND3X0 U35828 ( .IN1(m2s1_cyc), .IN2(n17917), .IN3(test_so43), .QN(n14474)
         );
  NAND3X0 U35829 ( .IN1(m6s0_cyc), .IN2(n18943), .IN3(s0_m6_cyc_r), .QN(n14488) );
  NAND3X0 U35830 ( .IN1(m2s0_cyc), .IN2(n17918), .IN3(s0_m2_cyc_r), .QN(n14484) );
  NAND3X0 U35831 ( .IN1(test_so32), .IN2(n20861), .IN3(s9_m6_cyc_r), .QN(
        n14398) );
  NAND3X0 U35832 ( .IN1(test_so22), .IN2(n20825), .IN3(s9_m2_cyc_r), .QN(
        n14394) );
  NAND3X0 U35833 ( .IN1(m6s8_cyc), .IN2(n20789), .IN3(s8_m6_cyc_r), .QN(n14408) );
  NAND3X0 U35834 ( .IN1(m2s8_cyc), .IN2(n17908), .IN3(s8_m2_cyc_r), .QN(n14404) );
  NAND3X0 U35835 ( .IN1(m1s9_cyc), .IN2(n20816), .IN3(s9_m1_cyc_r), .QN(n14393) );
  NAND3X0 U35836 ( .IN1(m0s7_cyc), .IN2(n20557), .IN3(s7_m0_cyc_r), .QN(n14412) );
  NAND3X0 U35837 ( .IN1(test_so17), .IN2(n20425), .IN3(s6_m0_cyc_r), .QN(
        n14422) );
  NAND3X0 U35838 ( .IN1(m0s14_cyc), .IN2(n19504), .IN3(s14_m0_cyc_r), .QN(
        n14342) );
  NAND3X0 U35839 ( .IN1(m0s5_cyc), .IN2(n20293), .IN3(test_so58), .QN(n14432)
         );
  NAND3X0 U35840 ( .IN1(m0s4_cyc), .IN2(n20162), .IN3(s4_m0_cyc_r), .QN(n14442) );
  NAND3X0 U35841 ( .IN1(test_so18), .IN2(n19372), .IN3(s13_m0_cyc_r), .QN(
        n14352) );
  NAND3X0 U35842 ( .IN1(m0s12_cyc), .IN2(n19240), .IN3(s12_m0_cyc_r), .QN(
        n14362) );
  NAND3X0 U35843 ( .IN1(m0s3_cyc), .IN2(n20031), .IN3(s3_m0_cyc_r), .QN(n14452) );
  NAND3X0 U35844 ( .IN1(m0s2_cyc), .IN2(n19900), .IN3(s2_m0_cyc_r), .QN(n14462) );
  NAND3X0 U35845 ( .IN1(m0s11_cyc), .IN2(n19108), .IN3(test_so81), .QN(n14372)
         );
  NAND3X0 U35846 ( .IN1(m0s10_cyc), .IN2(n18976), .IN3(s10_m0_cyc_r), .QN(
        n14382) );
  NAND3X0 U35847 ( .IN1(m0s1_cyc), .IN2(n19768), .IN3(s1_m0_cyc_r), .QN(n14472) );
  NAND3X0 U35848 ( .IN1(m0s0_cyc), .IN2(n18844), .IN3(s0_m0_cyc_r), .QN(n14482) );
  NAND3X0 U35849 ( .IN1(m0s8_cyc), .IN2(n20690), .IN3(s8_m0_cyc_r), .QN(n14402) );
  ISOLANDX1 U35850 ( .D(m7_cyc_i), .ISO(m7_stb_i), .Q(n14324) );
  ISOLANDX1 U35851 ( .D(m6_cyc_i), .ISO(m6_stb_i), .Q(n14326) );
  ISOLANDX1 U35852 ( .D(m4_cyc_i), .ISO(m4_stb_i), .Q(n14330) );
  ISOLANDX1 U35853 ( .D(m3_cyc_i), .ISO(m3_stb_i), .Q(n14332) );
  ISOLANDX1 U35854 ( .D(m2_cyc_i), .ISO(m2_stb_i), .Q(n14334) );
  ISOLANDX1 U35855 ( .D(m1_cyc_i), .ISO(m1_stb_i), .Q(n14336) );
  ISOLANDX1 U35856 ( .D(m0_cyc_i), .ISO(m0_stb_i), .Q(n14338) );
  ISOLANDX1 U35857 ( .D(m5_cyc_i), .ISO(m5_stb_i), .Q(n14328) );
  ISOLANDX1 U35858 ( .D(m7_cyc_i), .ISO(n14324), .Q(n14325) );
  ISOLANDX1 U35859 ( .D(m6_cyc_i), .ISO(n14326), .Q(n14327) );
  ISOLANDX1 U35860 ( .D(m4_cyc_i), .ISO(n14330), .Q(n14331) );
  ISOLANDX1 U35861 ( .D(m3_cyc_i), .ISO(n14332), .Q(n14333) );
  ISOLANDX1 U35862 ( .D(m2_cyc_i), .ISO(n14334), .Q(n14335) );
  ISOLANDX1 U35863 ( .D(m1_cyc_i), .ISO(n14336), .Q(n14337) );
  ISOLANDX1 U35864 ( .D(m0_cyc_i), .ISO(n14338), .Q(n14339) );
  ISOLANDX1 U35865 ( .D(m5_cyc_i), .ISO(n14328), .Q(n14329) );
  NAND3X0 U35866 ( .IN1(conf7_13_), .IN2(m6s7_cyc), .IN3(conf7_12_), .QN(
        n13883) );
  NAND3X0 U35867 ( .IN1(conf6_13_), .IN2(m6s6_cyc), .IN3(conf6_12_), .QN(
        n13574) );
  NAND3X0 U35868 ( .IN1(conf14_13_), .IN2(m6s14_cyc), .IN3(conf14_12_), .QN(
        n11408) );
  NAND3X0 U35869 ( .IN1(conf5_13_), .IN2(m6s5_cyc), .IN3(conf5_12_), .QN(
        n13265) );
  NAND3X0 U35870 ( .IN1(conf4_13_), .IN2(m6s4_cyc), .IN3(conf4_12_), .QN(
        n12956) );
  NAND3X0 U35871 ( .IN1(conf13_13_), .IN2(m6s13_cyc), .IN3(conf13_12_), .QN(
        n11099) );
  NAND3X0 U35872 ( .IN1(conf12_13_), .IN2(m6s12_cyc), .IN3(conf12_12_), .QN(
        n10789) );
  NAND3X0 U35873 ( .IN1(conf3_13_), .IN2(test_so31), .IN3(conf3_12_), .QN(
        n12647) );
  NAND3X0 U35874 ( .IN1(conf2_13_), .IN2(m6s2_cyc), .IN3(conf2_12_), .QN(
        n12338) );
  NAND3X0 U35875 ( .IN1(conf11_13_), .IN2(m6s11_cyc), .IN3(conf11_12_), .QN(
        n10480) );
  NAND3X0 U35876 ( .IN1(conf10_13_), .IN2(m6s10_cyc), .IN3(conf10_12_), .QN(
        n10170) );
  NAND3X0 U35877 ( .IN1(conf1_13_), .IN2(m6s1_cyc), .IN3(conf1_12_), .QN(
        n12028) );
  NAND3X0 U35878 ( .IN1(conf0_13_), .IN2(m6s0_cyc), .IN3(conf0_12_), .QN(
        n11718) );
  NAND3X0 U35879 ( .IN1(conf9_13_), .IN2(test_so32), .IN3(conf9_12_), .QN(
        n9860) );
  NAND3X0 U35880 ( .IN1(conf8_13_), .IN2(m6s8_cyc), .IN3(conf8_12_), .QN(n9549) );
  NAND3X0 U35881 ( .IN1(conf15_13_), .IN2(test_so33), .IN3(conf15_12_), .QN(
        n14157) );
  NAND3X0 U35882 ( .IN1(conf7_7_), .IN2(test_so24), .IN3(conf7_6_), .QN(n13888) );
  NAND3X0 U35883 ( .IN1(conf6_7_), .IN2(m3s6_cyc), .IN3(conf6_6_), .QN(n13579)
         );
  NAND3X0 U35884 ( .IN1(conf14_7_), .IN2(test_so25), .IN3(conf14_6_), .QN(
        n11413) );
  NAND3X0 U35885 ( .IN1(conf5_7_), .IN2(m3s5_cyc), .IN3(conf5_6_), .QN(n13270)
         );
  NAND3X0 U35886 ( .IN1(conf4_7_), .IN2(m3s4_cyc), .IN3(conf4_6_), .QN(n12961)
         );
  NAND3X0 U35887 ( .IN1(conf13_7_), .IN2(m3s13_cyc), .IN3(conf13_6_), .QN(
        n11104) );
  NAND3X0 U35888 ( .IN1(conf12_7_), .IN2(m3s12_cyc), .IN3(conf12_6_), .QN(
        n10794) );
  NAND3X0 U35889 ( .IN1(conf3_7_), .IN2(m3s3_cyc), .IN3(conf3_6_), .QN(n12652)
         );
  NAND3X0 U35890 ( .IN1(conf2_7_), .IN2(m3s2_cyc), .IN3(conf2_6_), .QN(n12343)
         );
  NAND3X0 U35891 ( .IN1(conf11_7_), .IN2(m3s11_cyc), .IN3(conf11_6_), .QN(
        n10485) );
  NAND3X0 U35892 ( .IN1(conf10_7_), .IN2(m3s10_cyc), .IN3(conf10_6_), .QN(
        n10175) );
  NAND3X0 U35893 ( .IN1(conf1_7_), .IN2(m3s1_cyc), .IN3(conf1_6_), .QN(n12033)
         );
  NAND3X0 U35894 ( .IN1(conf0_7_), .IN2(test_so23), .IN3(conf0_6_), .QN(n11723) );
  NAND3X0 U35895 ( .IN1(conf9_7_), .IN2(m3s9_cyc), .IN3(conf9_6_), .QN(n9865)
         );
  NAND3X0 U35896 ( .IN1(conf8_7_), .IN2(m3s8_cyc), .IN3(conf8_6_), .QN(n9554)
         );
  NAND3X0 U35897 ( .IN1(conf15_7_), .IN2(m3s15_cyc), .IN3(conf15_6_), .QN(
        n14162) );
  NAND3X0 U35898 ( .IN1(n3883), .IN2(n3885), .IN3(s7_msel_gnt_p3[1]), .QN(
        n13901) );
  NAND3X0 U35899 ( .IN1(n3838), .IN2(n3840), .IN3(s6_msel_gnt_p3_1_), .QN(
        n13592) );
  NAND3X0 U35900 ( .IN1(n4198), .IN2(n4200), .IN3(s14_msel_gnt_p3[1]), .QN(
        n11426) );
  NAND3X0 U35901 ( .IN1(n3793), .IN2(n3795), .IN3(test_so61), .QN(n13283) );
  NAND3X0 U35902 ( .IN1(n3748), .IN2(n3750), .IN3(s4_msel_gnt_p3_1_), .QN(
        n12974) );
  NAND3X0 U35903 ( .IN1(n4153), .IN2(n4155), .IN3(s13_msel_gnt_p3[1]), .QN(
        n11117) );
  NAND3X0 U35904 ( .IN1(n4108), .IN2(n4110), .IN3(s12_msel_gnt_p3_1_), .QN(
        n10807) );
  NAND3X0 U35905 ( .IN1(n3703), .IN2(n3705), .IN3(s3_msel_gnt_p3[1]), .QN(
        n12665) );
  NAND3X0 U35906 ( .IN1(n3658), .IN2(n3660), .IN3(s2_msel_gnt_p3[1]), .QN(
        n12356) );
  NAND3X0 U35907 ( .IN1(n4063), .IN2(n4065), .IN3(test_so84), .QN(n10498) );
  NAND3X0 U35908 ( .IN1(n4018), .IN2(n4020), .IN3(s10_msel_gnt_p3_1_), .QN(
        n10188) );
  NAND3X0 U35909 ( .IN1(n3613), .IN2(n3615), .IN3(s1_msel_gnt_p3[1]), .QN(
        n12046) );
  NAND3X0 U35910 ( .IN1(n3568), .IN2(n3570), .IN3(s0_msel_gnt_p3_1_), .QN(
        n11736) );
  NAND3X0 U35911 ( .IN1(n3973), .IN2(n3975), .IN3(s9_msel_gnt_p3[1]), .QN(
        n9878) );
  NAND3X0 U35912 ( .IN1(n3928), .IN2(n3930), .IN3(s8_msel_gnt_p3[1]), .QN(
        n9567) );
  NAND3X0 U35913 ( .IN1(n4227), .IN2(n4229), .IN3(s15_msel_gnt_p1[1]), .QN(
        n13967) );
  NAND3X0 U35914 ( .IN1(n4243), .IN2(n4245), .IN3(s15_msel_gnt_p3[1]), .QN(
        n14175) );
  NAND3X0 U35915 ( .IN1(n4235), .IN2(n4237), .IN3(s15_msel_gnt_p2_1_), .QN(
        n14107) );
  NAND3X0 U35916 ( .IN1(n3867), .IN2(n3869), .IN3(s7_msel_gnt_p1[1]), .QN(
        n13834) );
  NAND3X0 U35917 ( .IN1(n3875), .IN2(n3877), .IN3(s7_msel_gnt_p2_1_), .QN(
        n13707) );
  NAND3X0 U35918 ( .IN1(n3822), .IN2(n3824), .IN3(s6_msel_gnt_p1_1_), .QN(
        n13525) );
  NAND3X0 U35919 ( .IN1(n3830), .IN2(n3832), .IN3(s6_msel_gnt_p2[1]), .QN(
        n13398) );
  NAND3X0 U35920 ( .IN1(n4182), .IN2(n4184), .IN3(s14_msel_gnt_p1[1]), .QN(
        n11359) );
  NAND3X0 U35921 ( .IN1(n4190), .IN2(n4192), .IN3(test_so95), .QN(n11232) );
  NAND3X0 U35922 ( .IN1(n3777), .IN2(n3779), .IN3(test_so60), .QN(n13216) );
  NAND3X0 U35923 ( .IN1(n3785), .IN2(n3787), .IN3(s5_msel_gnt_p2[1]), .QN(
        n13089) );
  NAND3X0 U35924 ( .IN1(n3732), .IN2(n3734), .IN3(s4_msel_gnt_p1_1_), .QN(
        n12907) );
  NAND3X0 U35925 ( .IN1(n3740), .IN2(n3742), .IN3(s4_msel_gnt_p2[1]), .QN(
        n12780) );
  NAND3X0 U35926 ( .IN1(n4137), .IN2(n4139), .IN3(s13_msel_gnt_p1[1]), .QN(
        n11050) );
  NAND3X0 U35927 ( .IN1(n4145), .IN2(n4147), .IN3(s13_msel_gnt_p2_1_), .QN(
        n10923) );
  NAND3X0 U35928 ( .IN1(n4092), .IN2(n4094), .IN3(s12_msel_gnt_p1_1_), .QN(
        n10740) );
  NAND3X0 U35929 ( .IN1(n4100), .IN2(n4102), .IN3(s12_msel_gnt_p2[1]), .QN(
        n10613) );
  NAND3X0 U35930 ( .IN1(n3687), .IN2(n3689), .IN3(s3_msel_gnt_p1[1]), .QN(
        n12598) );
  NAND3X0 U35931 ( .IN1(n3695), .IN2(n3697), .IN3(s3_msel_gnt_p2_1_), .QN(
        n12471) );
  NAND3X0 U35932 ( .IN1(n3642), .IN2(n3644), .IN3(s2_msel_gnt_p1[1]), .QN(
        n12289) );
  NAND3X0 U35933 ( .IN1(n3650), .IN2(n3652), .IN3(test_so49), .QN(n12162) );
  NAND3X0 U35934 ( .IN1(n4047), .IN2(n4049), .IN3(test_so83), .QN(n10431) );
  NAND3X0 U35935 ( .IN1(n4055), .IN2(n4057), .IN3(s11_msel_gnt_p2[1]), .QN(
        n10304) );
  NAND3X0 U35936 ( .IN1(n4002), .IN2(n4004), .IN3(s10_msel_gnt_p1_1_), .QN(
        n10121) );
  NAND3X0 U35937 ( .IN1(n4010), .IN2(n4012), .IN3(s10_msel_gnt_p2[1]), .QN(
        n9994) );
  NAND3X0 U35938 ( .IN1(n3597), .IN2(n3599), .IN3(s1_msel_gnt_p1[1]), .QN(
        n11979) );
  NAND3X0 U35939 ( .IN1(n3605), .IN2(n3607), .IN3(s1_msel_gnt_p2_1_), .QN(
        n11852) );
  NAND3X0 U35940 ( .IN1(n3552), .IN2(n3554), .IN3(s0_msel_gnt_p1_1_), .QN(
        n11669) );
  NAND3X0 U35941 ( .IN1(n3560), .IN2(n3562), .IN3(s0_msel_gnt_p2[1]), .QN(
        n11542) );
  NAND3X0 U35942 ( .IN1(n3957), .IN2(n3959), .IN3(s9_msel_gnt_p1[1]), .QN(
        n9811) );
  NAND3X0 U35943 ( .IN1(n3965), .IN2(n3967), .IN3(s9_msel_gnt_p2_1_), .QN(
        n9684) );
  NAND3X0 U35944 ( .IN1(n3912), .IN2(n3914), .IN3(s8_msel_gnt_p1[1]), .QN(
        n9500) );
  NAND3X0 U35945 ( .IN1(n3920), .IN2(n3922), .IN3(test_so72), .QN(n9373) );
  ISOLANDX1 U35946 ( .D(m2s7_cyc), .ISO(n13646), .Q(n13673) );
  ISOLANDX1 U35947 ( .D(m2s6_cyc), .ISO(n13337), .Q(n13364) );
  ISOLANDX1 U35948 ( .D(m2s14_cyc), .ISO(n11171), .Q(n11198) );
  ISOLANDX1 U35949 ( .D(m2s5_cyc), .ISO(n13028), .Q(n13055) );
  ISOLANDX1 U35950 ( .D(m2s4_cyc), .ISO(n12719), .Q(n12746) );
  ISOLANDX1 U35951 ( .D(m2s13_cyc), .ISO(n10862), .Q(n10889) );
  ISOLANDX1 U35952 ( .D(m2s12_cyc), .ISO(n10552), .Q(n10579) );
  ISOLANDX1 U35953 ( .D(m2s3_cyc), .ISO(n12410), .Q(n12437) );
  ISOLANDX1 U35954 ( .D(test_so21), .ISO(n12101), .Q(n12128) );
  ISOLANDX1 U35955 ( .D(m2s11_cyc), .ISO(n10243), .Q(n10270) );
  ISOLANDX1 U35956 ( .D(m2s10_cyc), .ISO(n9933), .Q(n9960) );
  ISOLANDX1 U35957 ( .D(m2s1_cyc), .ISO(n11791), .Q(n11818) );
  ISOLANDX1 U35958 ( .D(m2s0_cyc), .ISO(n11481), .Q(n11508) );
  ISOLANDX1 U35959 ( .D(test_so22), .ISO(n9623), .Q(n9650) );
  ISOLANDX1 U35960 ( .D(m2s8_cyc), .ISO(n9312), .Q(n9339) );
  ISOLANDX1 U35961 ( .D(m2s15_cyc), .ISO(n14291), .Q(n14105) );
  NAND3X0 U35962 ( .IN1(conf7_3_), .IN2(m1s7_cyc), .IN3(conf7_2_), .QN(n13907)
         );
  NAND3X0 U35963 ( .IN1(conf6_3_), .IN2(m1s6_cyc), .IN3(conf6_2_), .QN(n13598)
         );
  NAND3X0 U35964 ( .IN1(conf14_3_), .IN2(m1s14_cyc), .IN3(conf14_2_), .QN(
        n11432) );
  NAND3X0 U35965 ( .IN1(conf5_3_), .IN2(m1s5_cyc), .IN3(conf5_2_), .QN(n13289)
         );
  NAND3X0 U35966 ( .IN1(conf4_3_), .IN2(test_so19), .IN3(conf4_2_), .QN(n12980) );
  NAND3X0 U35967 ( .IN1(conf13_3_), .IN2(m1s13_cyc), .IN3(conf13_2_), .QN(
        n11123) );
  NAND3X0 U35968 ( .IN1(conf12_3_), .IN2(m1s12_cyc), .IN3(conf12_2_), .QN(
        n10813) );
  NAND3X0 U35969 ( .IN1(conf3_3_), .IN2(m1s3_cyc), .IN3(conf3_2_), .QN(n12671)
         );
  NAND3X0 U35970 ( .IN1(conf2_3_), .IN2(m1s2_cyc), .IN3(conf2_2_), .QN(n12362)
         );
  NAND3X0 U35971 ( .IN1(conf11_3_), .IN2(test_so20), .IN3(conf11_2_), .QN(
        n10504) );
  NAND3X0 U35972 ( .IN1(conf10_3_), .IN2(m1s10_cyc), .IN3(conf10_2_), .QN(
        n10194) );
  NAND3X0 U35973 ( .IN1(conf1_3_), .IN2(m1s1_cyc), .IN3(conf1_2_), .QN(n12052)
         );
  NAND3X0 U35974 ( .IN1(conf0_3_), .IN2(m1s0_cyc), .IN3(conf0_2_), .QN(n11742)
         );
  NAND3X0 U35975 ( .IN1(conf9_3_), .IN2(m1s9_cyc), .IN3(conf9_2_), .QN(n9884)
         );
  NAND3X0 U35976 ( .IN1(conf8_3_), .IN2(m1s8_cyc), .IN3(conf8_2_), .QN(n9573)
         );
  NAND3X0 U35977 ( .IN1(conf15_3_), .IN2(m1s15_cyc), .IN3(conf15_2_), .QN(
        n14181) );
  NAND3X0 U35978 ( .IN1(s7_msel_gnt_p0_2_), .IN2(n3859), .IN3(
        s7_msel_gnt_p0_1_), .QN(n13758) );
  NAND3X0 U35979 ( .IN1(s6_msel_gnt_p0[2]), .IN2(n3814), .IN3(
        s6_msel_gnt_p0[1]), .QN(n13449) );
  NAND3X0 U35980 ( .IN1(s14_msel_gnt_p0_2_), .IN2(n4174), .IN3(test_so94), 
        .QN(n11283) );
  NAND3X0 U35981 ( .IN1(s5_msel_gnt_p0[2]), .IN2(n3769), .IN3(
        s5_msel_gnt_p0[1]), .QN(n13140) );
  NAND3X0 U35982 ( .IN1(s4_msel_gnt_p0[2]), .IN2(n3724), .IN3(
        s4_msel_gnt_p0[1]), .QN(n12831) );
  NAND3X0 U35983 ( .IN1(s13_msel_gnt_p0_2_), .IN2(n4129), .IN3(
        s13_msel_gnt_p0_1_), .QN(n10974) );
  NAND3X0 U35984 ( .IN1(s12_msel_gnt_p0[2]), .IN2(n4084), .IN3(
        s12_msel_gnt_p0[1]), .QN(n10664) );
  NAND3X0 U35985 ( .IN1(test_so52), .IN2(n3679), .IN3(s3_msel_gnt_p0_1_), .QN(
        n12522) );
  NAND3X0 U35986 ( .IN1(s2_msel_gnt_p0_2_), .IN2(n3634), .IN3(test_so48), .QN(
        n12213) );
  NAND3X0 U35987 ( .IN1(s11_msel_gnt_p0[2]), .IN2(n4039), .IN3(
        s11_msel_gnt_p0[1]), .QN(n10355) );
  NAND3X0 U35988 ( .IN1(s10_msel_gnt_p0[2]), .IN2(n3994), .IN3(
        s10_msel_gnt_p0[1]), .QN(n10045) );
  NAND3X0 U35989 ( .IN1(s1_msel_gnt_p0_2_), .IN2(n3589), .IN3(
        s1_msel_gnt_p0_1_), .QN(n11903) );
  NAND3X0 U35990 ( .IN1(s0_msel_gnt_p0[2]), .IN2(n3544), .IN3(
        s0_msel_gnt_p0[1]), .QN(n11593) );
  NAND3X0 U35991 ( .IN1(test_so75), .IN2(n3949), .IN3(s9_msel_gnt_p0_1_), .QN(
        n9735) );
  NAND3X0 U35992 ( .IN1(s8_msel_gnt_p0_2_), .IN2(n3904), .IN3(test_so71), .QN(
        n9424) );
  NAND3X0 U35993 ( .IN1(test_so98), .IN2(n4219), .IN3(s15_msel_gnt_p0_1_), 
        .QN(n14022) );
  ISOLANDX1 U35994 ( .D(m2s7_cyc), .ISO(n13645), .Q(n13832) );
  ISOLANDX1 U35995 ( .D(m2s6_cyc), .ISO(n13336), .Q(n13523) );
  ISOLANDX1 U35996 ( .D(m2s14_cyc), .ISO(n11170), .Q(n11357) );
  ISOLANDX1 U35997 ( .D(m2s5_cyc), .ISO(n13027), .Q(n13214) );
  ISOLANDX1 U35998 ( .D(m2s4_cyc), .ISO(n12718), .Q(n12905) );
  ISOLANDX1 U35999 ( .D(m2s13_cyc), .ISO(n10861), .Q(n11048) );
  ISOLANDX1 U36000 ( .D(m2s12_cyc), .ISO(n10551), .Q(n10738) );
  ISOLANDX1 U36001 ( .D(m2s3_cyc), .ISO(n12409), .Q(n12596) );
  ISOLANDX1 U36002 ( .D(test_so21), .ISO(n12100), .Q(n12287) );
  ISOLANDX1 U36003 ( .D(m2s11_cyc), .ISO(n10242), .Q(n10429) );
  ISOLANDX1 U36004 ( .D(m2s10_cyc), .ISO(n9932), .Q(n10119) );
  ISOLANDX1 U36005 ( .D(m2s1_cyc), .ISO(n11790), .Q(n11977) );
  ISOLANDX1 U36006 ( .D(m2s0_cyc), .ISO(n11480), .Q(n11667) );
  ISOLANDX1 U36007 ( .D(test_so22), .ISO(n9622), .Q(n9809) );
  ISOLANDX1 U36008 ( .D(m2s8_cyc), .ISO(n9311), .Q(n9498) );
  ISOLANDX1 U36009 ( .D(m2s15_cyc), .ISO(n14279), .Q(n13965) );
  ISOLANDX1 U36010 ( .D(m3s15_cyc), .ISO(n14290), .Q(n14090) );
  ISOLANDX1 U36011 ( .D(test_so24), .ISO(n13643), .Q(n13674) );
  ISOLANDX1 U36012 ( .D(m3s6_cyc), .ISO(n13334), .Q(n13365) );
  ISOLANDX1 U36013 ( .D(test_so25), .ISO(n11168), .Q(n11199) );
  ISOLANDX1 U36014 ( .D(m3s5_cyc), .ISO(n13025), .Q(n13056) );
  ISOLANDX1 U36015 ( .D(m3s4_cyc), .ISO(n12716), .Q(n12747) );
  ISOLANDX1 U36016 ( .D(m3s13_cyc), .ISO(n10859), .Q(n10890) );
  ISOLANDX1 U36017 ( .D(m3s12_cyc), .ISO(n10549), .Q(n10580) );
  ISOLANDX1 U36018 ( .D(m3s3_cyc), .ISO(n12407), .Q(n12438) );
  ISOLANDX1 U36019 ( .D(m3s2_cyc), .ISO(n12098), .Q(n12129) );
  ISOLANDX1 U36020 ( .D(m3s11_cyc), .ISO(n10240), .Q(n10271) );
  ISOLANDX1 U36021 ( .D(m3s10_cyc), .ISO(n9930), .Q(n9961) );
  ISOLANDX1 U36022 ( .D(m3s1_cyc), .ISO(n11788), .Q(n11819) );
  ISOLANDX1 U36023 ( .D(test_so23), .ISO(n11478), .Q(n11509) );
  ISOLANDX1 U36024 ( .D(m3s9_cyc), .ISO(n9620), .Q(n9651) );
  ISOLANDX1 U36025 ( .D(m3s8_cyc), .ISO(n9309), .Q(n9340) );
  NAND3X0 U36026 ( .IN1(conf7_5_), .IN2(m2s7_cyc), .IN3(conf7_4_), .QN(n13894)
         );
  NAND3X0 U36027 ( .IN1(conf6_5_), .IN2(m2s6_cyc), .IN3(conf6_4_), .QN(n13585)
         );
  NAND3X0 U36028 ( .IN1(conf14_5_), .IN2(m2s14_cyc), .IN3(conf14_4_), .QN(
        n11419) );
  NAND3X0 U36029 ( .IN1(conf5_5_), .IN2(m2s5_cyc), .IN3(conf5_4_), .QN(n13276)
         );
  NAND3X0 U36030 ( .IN1(conf4_5_), .IN2(m2s4_cyc), .IN3(conf4_4_), .QN(n12967)
         );
  NAND3X0 U36031 ( .IN1(conf13_5_), .IN2(m2s13_cyc), .IN3(conf13_4_), .QN(
        n11110) );
  NAND3X0 U36032 ( .IN1(conf12_5_), .IN2(m2s12_cyc), .IN3(conf12_4_), .QN(
        n10800) );
  NAND3X0 U36033 ( .IN1(conf3_5_), .IN2(m2s3_cyc), .IN3(conf3_4_), .QN(n12658)
         );
  NAND3X0 U36034 ( .IN1(conf2_5_), .IN2(test_so21), .IN3(conf2_4_), .QN(n12349) );
  NAND3X0 U36035 ( .IN1(conf11_5_), .IN2(m2s11_cyc), .IN3(conf11_4_), .QN(
        n10491) );
  NAND3X0 U36036 ( .IN1(conf10_5_), .IN2(m2s10_cyc), .IN3(conf10_4_), .QN(
        n10181) );
  NAND3X0 U36037 ( .IN1(conf1_5_), .IN2(m2s1_cyc), .IN3(conf1_4_), .QN(n12039)
         );
  NAND3X0 U36038 ( .IN1(conf0_5_), .IN2(m2s0_cyc), .IN3(conf0_4_), .QN(n11729)
         );
  NAND3X0 U36039 ( .IN1(conf9_5_), .IN2(test_so22), .IN3(conf9_4_), .QN(n9871)
         );
  NAND3X0 U36040 ( .IN1(conf8_5_), .IN2(m2s8_cyc), .IN3(conf8_4_), .QN(n9560)
         );
  NAND3X0 U36041 ( .IN1(conf15_5_), .IN2(m2s15_cyc), .IN3(conf15_4_), .QN(
        n14168) );
  NAND3X0 U36042 ( .IN1(s7_msel_gnt_p3[1]), .IN2(n3885), .IN3(
        s7_msel_gnt_p3[0]), .QN(n13885) );
  NAND3X0 U36043 ( .IN1(s6_msel_gnt_p3_1_), .IN2(n3840), .IN3(
        s6_msel_gnt_p3_0_), .QN(n13576) );
  NAND3X0 U36044 ( .IN1(s14_msel_gnt_p3[1]), .IN2(n4200), .IN3(
        s14_msel_gnt_p3[0]), .QN(n11410) );
  NAND3X0 U36045 ( .IN1(test_so61), .IN2(n3795), .IN3(s5_msel_gnt_p3_0_), .QN(
        n13267) );
  NAND3X0 U36046 ( .IN1(s4_msel_gnt_p3_1_), .IN2(n3750), .IN3(test_so57), .QN(
        n12958) );
  NAND3X0 U36047 ( .IN1(s13_msel_gnt_p3[1]), .IN2(n4155), .IN3(
        s13_msel_gnt_p3[0]), .QN(n11101) );
  NAND3X0 U36048 ( .IN1(s12_msel_gnt_p3_1_), .IN2(n4110), .IN3(
        s12_msel_gnt_p3_0_), .QN(n10791) );
  NAND3X0 U36049 ( .IN1(s3_msel_gnt_p3[1]), .IN2(n3705), .IN3(
        s3_msel_gnt_p3[0]), .QN(n12649) );
  NAND3X0 U36050 ( .IN1(s2_msel_gnt_p3[1]), .IN2(n3660), .IN3(
        s2_msel_gnt_p3[0]), .QN(n12340) );
  NAND3X0 U36051 ( .IN1(test_so84), .IN2(n4065), .IN3(s11_msel_gnt_p3_0_), 
        .QN(n10482) );
  NAND3X0 U36052 ( .IN1(s10_msel_gnt_p3_1_), .IN2(n4020), .IN3(test_so80), 
        .QN(n10172) );
  NAND3X0 U36053 ( .IN1(s1_msel_gnt_p3[1]), .IN2(n3615), .IN3(
        s1_msel_gnt_p3[0]), .QN(n12030) );
  NAND3X0 U36054 ( .IN1(s0_msel_gnt_p3_1_), .IN2(n3570), .IN3(
        s0_msel_gnt_p3_0_), .QN(n11720) );
  NAND3X0 U36055 ( .IN1(s9_msel_gnt_p3[1]), .IN2(n3975), .IN3(
        s9_msel_gnt_p3[0]), .QN(n9862) );
  NAND3X0 U36056 ( .IN1(s8_msel_gnt_p3[1]), .IN2(n3930), .IN3(
        s8_msel_gnt_p3[0]), .QN(n9551) );
  NAND3X0 U36057 ( .IN1(s15_msel_gnt_p1[1]), .IN2(n4229), .IN3(
        s15_msel_gnt_p1[0]), .QN(n13948) );
  NAND3X0 U36058 ( .IN1(s15_msel_gnt_p3[1]), .IN2(n4245), .IN3(
        s15_msel_gnt_p3[0]), .QN(n14159) );
  NAND3X0 U36059 ( .IN1(s15_msel_gnt_p2_1_), .IN2(n4237), .IN3(
        s15_msel_gnt_p2_0_), .QN(n14088) );
  NAND3X0 U36060 ( .IN1(s7_msel_gnt_p1[1]), .IN2(n3869), .IN3(
        s7_msel_gnt_p1[0]), .QN(n13816) );
  NAND3X0 U36061 ( .IN1(s7_msel_gnt_p2_1_), .IN2(n3877), .IN3(test_so68), .QN(
        n13691) );
  NAND3X0 U36062 ( .IN1(s6_msel_gnt_p1_1_), .IN2(n3824), .IN3(
        s6_msel_gnt_p1_0_), .QN(n13507) );
  NAND3X0 U36063 ( .IN1(s6_msel_gnt_p2[1]), .IN2(n3832), .IN3(
        s6_msel_gnt_p2[0]), .QN(n13382) );
  NAND3X0 U36064 ( .IN1(s14_msel_gnt_p1[1]), .IN2(n4184), .IN3(
        s14_msel_gnt_p1[0]), .QN(n11341) );
  NAND3X0 U36065 ( .IN1(test_so95), .IN2(n4192), .IN3(s14_msel_gnt_p2_0_), 
        .QN(n11216) );
  NAND3X0 U36066 ( .IN1(test_so60), .IN2(n3779), .IN3(s5_msel_gnt_p1_0_), .QN(
        n13198) );
  NAND3X0 U36067 ( .IN1(s5_msel_gnt_p2[1]), .IN2(n3787), .IN3(
        s5_msel_gnt_p2[0]), .QN(n13073) );
  NAND3X0 U36068 ( .IN1(s4_msel_gnt_p1_1_), .IN2(n3734), .IN3(test_so56), .QN(
        n12889) );
  NAND3X0 U36069 ( .IN1(s4_msel_gnt_p2[1]), .IN2(n3742), .IN3(
        s4_msel_gnt_p2[0]), .QN(n12764) );
  NAND3X0 U36070 ( .IN1(s13_msel_gnt_p1[1]), .IN2(n4139), .IN3(
        s13_msel_gnt_p1[0]), .QN(n11032) );
  NAND3X0 U36071 ( .IN1(s13_msel_gnt_p2_1_), .IN2(n4147), .IN3(test_so91), 
        .QN(n10907) );
  NAND3X0 U36072 ( .IN1(s12_msel_gnt_p1_1_), .IN2(n4094), .IN3(
        s12_msel_gnt_p1_0_), .QN(n10722) );
  NAND3X0 U36073 ( .IN1(s12_msel_gnt_p2[1]), .IN2(n4102), .IN3(
        s12_msel_gnt_p2[0]), .QN(n10597) );
  NAND3X0 U36074 ( .IN1(s3_msel_gnt_p1[1]), .IN2(n3689), .IN3(
        s3_msel_gnt_p1[0]), .QN(n12580) );
  NAND3X0 U36075 ( .IN1(s3_msel_gnt_p2_1_), .IN2(n3697), .IN3(
        s3_msel_gnt_p2_0_), .QN(n12455) );
  NAND3X0 U36076 ( .IN1(s2_msel_gnt_p1[1]), .IN2(n3644), .IN3(
        s2_msel_gnt_p1[0]), .QN(n12271) );
  NAND3X0 U36077 ( .IN1(test_so49), .IN2(n3652), .IN3(s2_msel_gnt_p2_0_), .QN(
        n12146) );
  NAND3X0 U36078 ( .IN1(test_so83), .IN2(n4049), .IN3(s11_msel_gnt_p1_0_), 
        .QN(n10413) );
  NAND3X0 U36079 ( .IN1(s11_msel_gnt_p2[1]), .IN2(n4057), .IN3(
        s11_msel_gnt_p2[0]), .QN(n10288) );
  NAND3X0 U36080 ( .IN1(s10_msel_gnt_p1_1_), .IN2(n4004), .IN3(test_so79), 
        .QN(n10103) );
  NAND3X0 U36081 ( .IN1(s10_msel_gnt_p2[1]), .IN2(n4012), .IN3(
        s10_msel_gnt_p2[0]), .QN(n9978) );
  NAND3X0 U36082 ( .IN1(s1_msel_gnt_p1[1]), .IN2(n3599), .IN3(
        s1_msel_gnt_p1[0]), .QN(n11961) );
  NAND3X0 U36083 ( .IN1(s1_msel_gnt_p2_1_), .IN2(n3607), .IN3(test_so45), .QN(
        n11836) );
  NAND3X0 U36084 ( .IN1(s0_msel_gnt_p1_1_), .IN2(n3554), .IN3(
        s0_msel_gnt_p1_0_), .QN(n11651) );
  NAND3X0 U36085 ( .IN1(s0_msel_gnt_p2[1]), .IN2(n3562), .IN3(
        s0_msel_gnt_p2[0]), .QN(n11526) );
  NAND3X0 U36086 ( .IN1(s9_msel_gnt_p1[1]), .IN2(n3959), .IN3(
        s9_msel_gnt_p1[0]), .QN(n9793) );
  NAND3X0 U36087 ( .IN1(s9_msel_gnt_p2_1_), .IN2(n3967), .IN3(
        s9_msel_gnt_p2_0_), .QN(n9668) );
  NAND3X0 U36088 ( .IN1(s8_msel_gnt_p1[1]), .IN2(n3914), .IN3(
        s8_msel_gnt_p1[0]), .QN(n9482) );
  NAND3X0 U36089 ( .IN1(test_so72), .IN2(n3922), .IN3(s8_msel_gnt_p2_0_), .QN(
        n9357) );
  ISOLANDX1 U36090 ( .D(m7s7_cyc), .ISO(n13659), .Q(n13678) );
  ISOLANDX1 U36091 ( .D(m7s6_cyc), .ISO(n13350), .Q(n13369) );
  ISOLANDX1 U36092 ( .D(m7s14_cyc), .ISO(n11184), .Q(n11203) );
  ISOLANDX1 U36093 ( .D(test_so34), .ISO(n13041), .Q(n13060) );
  ISOLANDX1 U36094 ( .D(m7s4_cyc), .ISO(n12732), .Q(n12751) );
  ISOLANDX1 U36095 ( .D(m7s13_cyc), .ISO(n10875), .Q(n10894) );
  ISOLANDX1 U36096 ( .D(m7s12_cyc), .ISO(n10565), .Q(n10584) );
  ISOLANDX1 U36097 ( .D(m7s3_cyc), .ISO(n12423), .Q(n12442) );
  ISOLANDX1 U36098 ( .D(m7s2_cyc), .ISO(n12114), .Q(n12133) );
  ISOLANDX1 U36099 ( .D(test_so35), .ISO(n10256), .Q(n10275) );
  ISOLANDX1 U36100 ( .D(m7s10_cyc), .ISO(n9946), .Q(n9965) );
  ISOLANDX1 U36101 ( .D(m7s1_cyc), .ISO(n11804), .Q(n11823) );
  ISOLANDX1 U36102 ( .D(m7s0_cyc), .ISO(n11494), .Q(n11513) );
  ISOLANDX1 U36103 ( .D(m7s9_cyc), .ISO(n9636), .Q(n9655) );
  ISOLANDX1 U36104 ( .D(m7s8_cyc), .ISO(n9325), .Q(n9344) );
  NAND3X0 U36105 ( .IN1(s6_msel_gnt_p0[2]), .IN2(n3815), .IN3(
        s6_msel_gnt_p0[0]), .QN(n13448) );
  NAND3X0 U36106 ( .IN1(s13_msel_gnt_p0_2_), .IN2(n4130), .IN3(test_so90), 
        .QN(n10973) );
  NAND3X0 U36107 ( .IN1(s11_msel_gnt_p0[2]), .IN2(n4040), .IN3(
        s11_msel_gnt_p0[0]), .QN(n10354) );
  NAND3X0 U36108 ( .IN1(test_so75), .IN2(n3950), .IN3(s9_msel_gnt_p0_0_), .QN(
        n9734) );
  NAND3X0 U36109 ( .IN1(s7_msel_gnt_p0_2_), .IN2(n3860), .IN3(test_so67), .QN(
        n13757) );
  NAND3X0 U36110 ( .IN1(s14_msel_gnt_p0_2_), .IN2(n4175), .IN3(
        s14_msel_gnt_p0_0_), .QN(n11282) );
  NAND3X0 U36111 ( .IN1(s5_msel_gnt_p0[2]), .IN2(n3770), .IN3(
        s5_msel_gnt_p0[0]), .QN(n13139) );
  NAND3X0 U36112 ( .IN1(s4_msel_gnt_p0[2]), .IN2(n3725), .IN3(
        s4_msel_gnt_p0[0]), .QN(n12830) );
  NAND3X0 U36113 ( .IN1(s12_msel_gnt_p0[2]), .IN2(n4085), .IN3(
        s12_msel_gnt_p0[0]), .QN(n10663) );
  NAND3X0 U36114 ( .IN1(test_so52), .IN2(n3680), .IN3(s3_msel_gnt_p0_0_), .QN(
        n12521) );
  NAND3X0 U36115 ( .IN1(s2_msel_gnt_p0_2_), .IN2(n3635), .IN3(
        s2_msel_gnt_p0_0_), .QN(n12212) );
  NAND3X0 U36116 ( .IN1(s10_msel_gnt_p0[2]), .IN2(n3995), .IN3(
        s10_msel_gnt_p0[0]), .QN(n10044) );
  NAND3X0 U36117 ( .IN1(s1_msel_gnt_p0_2_), .IN2(n3590), .IN3(test_so44), .QN(
        n11902) );
  NAND3X0 U36118 ( .IN1(s0_msel_gnt_p0[2]), .IN2(n3545), .IN3(
        s0_msel_gnt_p0[0]), .QN(n11592) );
  NAND3X0 U36119 ( .IN1(s8_msel_gnt_p0_2_), .IN2(n3905), .IN3(
        s8_msel_gnt_p0_0_), .QN(n9423) );
  NAND3X0 U36120 ( .IN1(test_so98), .IN2(n4220), .IN3(s15_msel_gnt_p0_0_), 
        .QN(n14021) );
  NAND3X0 U36121 ( .IN1(conf7_1_), .IN2(m0s7_cyc), .IN3(test_so8), .QN(n13928)
         );
  NAND3X0 U36122 ( .IN1(conf6_1_), .IN2(test_so17), .IN3(test_so7), .QN(n13619) );
  NAND3X0 U36123 ( .IN1(conf14_1_), .IN2(m0s14_cyc), .IN3(test_so15), .QN(
        n11453) );
  NAND3X0 U36124 ( .IN1(conf5_1_), .IN2(m0s5_cyc), .IN3(test_so6), .QN(n13310)
         );
  NAND3X0 U36125 ( .IN1(conf4_1_), .IN2(m0s4_cyc), .IN3(test_so5), .QN(n13001)
         );
  NAND3X0 U36126 ( .IN1(conf13_1_), .IN2(test_so18), .IN3(test_so14), .QN(
        n11144) );
  NAND3X0 U36127 ( .IN1(conf12_1_), .IN2(m0s12_cyc), .IN3(test_so13), .QN(
        n10834) );
  NAND3X0 U36128 ( .IN1(conf3_1_), .IN2(m0s3_cyc), .IN3(test_so4), .QN(n12692)
         );
  NAND3X0 U36129 ( .IN1(conf2_1_), .IN2(m0s2_cyc), .IN3(test_so3), .QN(n12383)
         );
  NAND3X0 U36130 ( .IN1(conf11_1_), .IN2(m0s11_cyc), .IN3(test_so12), .QN(
        n10525) );
  NAND3X0 U36131 ( .IN1(conf10_1_), .IN2(m0s10_cyc), .IN3(test_so11), .QN(
        n10215) );
  NAND3X0 U36132 ( .IN1(conf1_1_), .IN2(m0s1_cyc), .IN3(test_so2), .QN(n12073)
         );
  NAND3X0 U36133 ( .IN1(conf0_1_), .IN2(m0s0_cyc), .IN3(test_so1), .QN(n11763)
         );
  NAND3X0 U36134 ( .IN1(conf9_1_), .IN2(m0s9_cyc), .IN3(test_so10), .QN(n9905)
         );
  NAND3X0 U36135 ( .IN1(conf8_1_), .IN2(m0s8_cyc), .IN3(test_so9), .QN(n9594)
         );
  NAND3X0 U36136 ( .IN1(conf15_1_), .IN2(m0s15_cyc), .IN3(test_so16), .QN(
        n14202) );
  ISOLANDX1 U36137 ( .D(m1s7_cyc), .ISO(n13649), .Q(n13675) );
  ISOLANDX1 U36138 ( .D(m1s6_cyc), .ISO(n13340), .Q(n13366) );
  ISOLANDX1 U36139 ( .D(m1s14_cyc), .ISO(n11174), .Q(n11200) );
  ISOLANDX1 U36140 ( .D(m1s5_cyc), .ISO(n13031), .Q(n13057) );
  ISOLANDX1 U36141 ( .D(test_so19), .ISO(n12722), .Q(n12748) );
  ISOLANDX1 U36142 ( .D(m1s13_cyc), .ISO(n10865), .Q(n10891) );
  ISOLANDX1 U36143 ( .D(m1s12_cyc), .ISO(n10555), .Q(n10581) );
  ISOLANDX1 U36144 ( .D(m1s3_cyc), .ISO(n12413), .Q(n12439) );
  ISOLANDX1 U36145 ( .D(m1s2_cyc), .ISO(n12104), .Q(n12130) );
  ISOLANDX1 U36146 ( .D(test_so20), .ISO(n10246), .Q(n10272) );
  ISOLANDX1 U36147 ( .D(m1s10_cyc), .ISO(n9936), .Q(n9962) );
  ISOLANDX1 U36148 ( .D(m1s1_cyc), .ISO(n11794), .Q(n11820) );
  ISOLANDX1 U36149 ( .D(m1s0_cyc), .ISO(n11484), .Q(n11510) );
  ISOLANDX1 U36150 ( .D(m1s9_cyc), .ISO(n9626), .Q(n9652) );
  ISOLANDX1 U36151 ( .D(m1s8_cyc), .ISO(n9315), .Q(n9341) );
  ISOLANDX1 U36152 ( .D(m1s15_cyc), .ISO(n14292), .Q(n14108) );
  ISOLANDX1 U36153 ( .D(m6s7_cyc), .ISO(n13661), .Q(n13838) );
  ISOLANDX1 U36154 ( .D(m6s6_cyc), .ISO(n13352), .Q(n13529) );
  ISOLANDX1 U36155 ( .D(m6s14_cyc), .ISO(n11186), .Q(n11363) );
  ISOLANDX1 U36156 ( .D(m6s5_cyc), .ISO(n13043), .Q(n13220) );
  ISOLANDX1 U36157 ( .D(m6s4_cyc), .ISO(n12734), .Q(n12911) );
  ISOLANDX1 U36158 ( .D(m6s13_cyc), .ISO(n10877), .Q(n11054) );
  ISOLANDX1 U36159 ( .D(m6s12_cyc), .ISO(n10567), .Q(n10744) );
  ISOLANDX1 U36160 ( .D(test_so31), .ISO(n12425), .Q(n12602) );
  ISOLANDX1 U36161 ( .D(m6s2_cyc), .ISO(n12116), .Q(n12293) );
  ISOLANDX1 U36162 ( .D(m6s11_cyc), .ISO(n10258), .Q(n10435) );
  ISOLANDX1 U36163 ( .D(m6s10_cyc), .ISO(n9948), .Q(n10125) );
  ISOLANDX1 U36164 ( .D(m6s1_cyc), .ISO(n11806), .Q(n11983) );
  ISOLANDX1 U36165 ( .D(m6s0_cyc), .ISO(n11496), .Q(n11673) );
  ISOLANDX1 U36166 ( .D(test_so32), .ISO(n9638), .Q(n9815) );
  ISOLANDX1 U36167 ( .D(m6s8_cyc), .ISO(n9327), .Q(n9504) );
  ISOLANDX1 U36168 ( .D(m7s15_cyc), .ISO(n14298), .Q(n14127) );
  ISOLANDX1 U36169 ( .D(test_so33), .ISO(n14283), .Q(n13971) );
  ISOLANDX1 U36170 ( .D(test_so33), .ISO(n14299), .Q(n14111) );
  ISOLANDX1 U36171 ( .D(test_so24), .ISO(n13642), .Q(n13818) );
  ISOLANDX1 U36172 ( .D(m3s6_cyc), .ISO(n13333), .Q(n13509) );
  ISOLANDX1 U36173 ( .D(test_so25), .ISO(n11167), .Q(n11343) );
  ISOLANDX1 U36174 ( .D(m3s5_cyc), .ISO(n13024), .Q(n13200) );
  ISOLANDX1 U36175 ( .D(m3s4_cyc), .ISO(n12715), .Q(n12891) );
  ISOLANDX1 U36176 ( .D(m3s13_cyc), .ISO(n10858), .Q(n11034) );
  ISOLANDX1 U36177 ( .D(m3s12_cyc), .ISO(n10548), .Q(n10724) );
  ISOLANDX1 U36178 ( .D(m3s3_cyc), .ISO(n12406), .Q(n12582) );
  ISOLANDX1 U36179 ( .D(m3s2_cyc), .ISO(n12097), .Q(n12273) );
  ISOLANDX1 U36180 ( .D(m3s11_cyc), .ISO(n10239), .Q(n10415) );
  ISOLANDX1 U36181 ( .D(m3s10_cyc), .ISO(n9929), .Q(n10105) );
  ISOLANDX1 U36182 ( .D(m3s1_cyc), .ISO(n11787), .Q(n11963) );
  ISOLANDX1 U36183 ( .D(test_so23), .ISO(n11477), .Q(n11653) );
  ISOLANDX1 U36184 ( .D(m3s9_cyc), .ISO(n9619), .Q(n9795) );
  ISOLANDX1 U36185 ( .D(m3s8_cyc), .ISO(n9308), .Q(n9484) );
  ISOLANDX1 U36186 ( .D(m3s15_cyc), .ISO(n14276), .Q(n13950) );
  ISOLANDX1 U36187 ( .D(m6s7_cyc), .ISO(n13660), .Q(n13775) );
  ISOLANDX1 U36188 ( .D(m6s6_cyc), .ISO(n13351), .Q(n13466) );
  ISOLANDX1 U36189 ( .D(m6s14_cyc), .ISO(n11185), .Q(n11300) );
  ISOLANDX1 U36190 ( .D(m6s5_cyc), .ISO(n13042), .Q(n13157) );
  ISOLANDX1 U36191 ( .D(m6s4_cyc), .ISO(n12733), .Q(n12848) );
  ISOLANDX1 U36192 ( .D(m6s13_cyc), .ISO(n10876), .Q(n10991) );
  ISOLANDX1 U36193 ( .D(m6s12_cyc), .ISO(n10566), .Q(n10681) );
  ISOLANDX1 U36194 ( .D(test_so31), .ISO(n12424), .Q(n12539) );
  ISOLANDX1 U36195 ( .D(m6s2_cyc), .ISO(n12115), .Q(n12230) );
  ISOLANDX1 U36196 ( .D(m6s11_cyc), .ISO(n10257), .Q(n10372) );
  ISOLANDX1 U36197 ( .D(m6s10_cyc), .ISO(n9947), .Q(n10062) );
  ISOLANDX1 U36198 ( .D(m6s1_cyc), .ISO(n11805), .Q(n11920) );
  ISOLANDX1 U36199 ( .D(m6s0_cyc), .ISO(n11495), .Q(n11610) );
  ISOLANDX1 U36200 ( .D(test_so32), .ISO(n9637), .Q(n9752) );
  ISOLANDX1 U36201 ( .D(m6s8_cyc), .ISO(n9326), .Q(n9441) );
  ISOLANDX1 U36202 ( .D(test_so33), .ISO(n14068), .Q(n14039) );
  ISOLANDX1 U36203 ( .D(m0s15_cyc), .ISO(n14293), .Q(n14120) );
  NAND3X0 U36204 ( .IN1(conf7_15_), .IN2(m7s7_cyc), .IN3(conf7_14_), .QN(
        n13876) );
  NAND3X0 U36205 ( .IN1(conf6_15_), .IN2(m7s6_cyc), .IN3(conf6_14_), .QN(
        n13567) );
  NAND3X0 U36206 ( .IN1(conf14_15_), .IN2(m7s14_cyc), .IN3(conf14_14_), .QN(
        n11401) );
  NAND3X0 U36207 ( .IN1(conf5_15_), .IN2(test_so34), .IN3(conf5_14_), .QN(
        n13258) );
  NAND3X0 U36208 ( .IN1(conf4_15_), .IN2(m7s4_cyc), .IN3(conf4_14_), .QN(
        n12949) );
  NAND3X0 U36209 ( .IN1(conf13_15_), .IN2(m7s13_cyc), .IN3(conf13_14_), .QN(
        n11092) );
  NAND3X0 U36210 ( .IN1(conf12_15_), .IN2(m7s12_cyc), .IN3(conf12_14_), .QN(
        n10782) );
  NAND3X0 U36211 ( .IN1(conf3_15_), .IN2(m7s3_cyc), .IN3(conf3_14_), .QN(
        n12640) );
  NAND3X0 U36212 ( .IN1(conf2_15_), .IN2(m7s2_cyc), .IN3(conf2_14_), .QN(
        n12331) );
  NAND3X0 U36213 ( .IN1(conf11_15_), .IN2(test_so35), .IN3(conf11_14_), .QN(
        n10473) );
  NAND3X0 U36214 ( .IN1(conf10_15_), .IN2(m7s10_cyc), .IN3(conf10_14_), .QN(
        n10163) );
  NAND3X0 U36215 ( .IN1(conf1_15_), .IN2(m7s1_cyc), .IN3(conf1_14_), .QN(
        n12021) );
  NAND3X0 U36216 ( .IN1(conf0_15_), .IN2(m7s0_cyc), .IN3(conf0_14_), .QN(
        n11711) );
  NAND3X0 U36217 ( .IN1(conf9_15_), .IN2(m7s9_cyc), .IN3(conf9_14_), .QN(n9853) );
  NAND3X0 U36218 ( .IN1(conf8_15_), .IN2(m7s8_cyc), .IN3(conf8_14_), .QN(n9542) );
  NAND3X0 U36219 ( .IN1(conf15_15_), .IN2(m7s15_cyc), .IN3(conf15_14_), .QN(
        n14150) );
  ISOLANDX1 U36220 ( .D(m1s7_cyc), .ISO(n13648), .Q(n13835) );
  ISOLANDX1 U36221 ( .D(m1s6_cyc), .ISO(n13339), .Q(n13526) );
  ISOLANDX1 U36222 ( .D(m1s14_cyc), .ISO(n11173), .Q(n11360) );
  ISOLANDX1 U36223 ( .D(m1s5_cyc), .ISO(n13030), .Q(n13217) );
  ISOLANDX1 U36224 ( .D(test_so19), .ISO(n12721), .Q(n12908) );
  ISOLANDX1 U36225 ( .D(m1s13_cyc), .ISO(n10864), .Q(n11051) );
  ISOLANDX1 U36226 ( .D(m1s12_cyc), .ISO(n10554), .Q(n10741) );
  ISOLANDX1 U36227 ( .D(m1s3_cyc), .ISO(n12412), .Q(n12599) );
  ISOLANDX1 U36228 ( .D(m1s2_cyc), .ISO(n12103), .Q(n12290) );
  ISOLANDX1 U36229 ( .D(test_so20), .ISO(n10245), .Q(n10432) );
  ISOLANDX1 U36230 ( .D(m1s10_cyc), .ISO(n9935), .Q(n10122) );
  ISOLANDX1 U36231 ( .D(m1s1_cyc), .ISO(n11793), .Q(n11980) );
  ISOLANDX1 U36232 ( .D(m1s0_cyc), .ISO(n11483), .Q(n11670) );
  ISOLANDX1 U36233 ( .D(m1s9_cyc), .ISO(n9625), .Q(n9812) );
  ISOLANDX1 U36234 ( .D(m1s8_cyc), .ISO(n9314), .Q(n9501) );
  ISOLANDX1 U36235 ( .D(m1s15_cyc), .ISO(n14278), .Q(n13968) );
  NAND3X0 U36236 ( .IN1(n3814), .IN2(n3815), .IN3(s6_msel_gnt_p0[2]), .QN(
        n13473) );
  NAND3X0 U36237 ( .IN1(n4129), .IN2(n4130), .IN3(s13_msel_gnt_p0_2_), .QN(
        n10998) );
  NAND3X0 U36238 ( .IN1(n4039), .IN2(n4040), .IN3(s11_msel_gnt_p0[2]), .QN(
        n10379) );
  NAND3X0 U36239 ( .IN1(n3949), .IN2(n3950), .IN3(test_so75), .QN(n9759) );
  NAND3X0 U36240 ( .IN1(n3859), .IN2(n3860), .IN3(s7_msel_gnt_p0_2_), .QN(
        n13782) );
  NAND3X0 U36241 ( .IN1(n4174), .IN2(n4175), .IN3(s14_msel_gnt_p0_2_), .QN(
        n11307) );
  NAND3X0 U36242 ( .IN1(n3769), .IN2(n3770), .IN3(s5_msel_gnt_p0[2]), .QN(
        n13164) );
  NAND3X0 U36243 ( .IN1(n3724), .IN2(n3725), .IN3(s4_msel_gnt_p0[2]), .QN(
        n12855) );
  NAND3X0 U36244 ( .IN1(n4084), .IN2(n4085), .IN3(s12_msel_gnt_p0[2]), .QN(
        n10688) );
  NAND3X0 U36245 ( .IN1(n3679), .IN2(n3680), .IN3(test_so52), .QN(n12546) );
  NAND3X0 U36246 ( .IN1(n3634), .IN2(n3635), .IN3(s2_msel_gnt_p0_2_), .QN(
        n12237) );
  NAND3X0 U36247 ( .IN1(n3994), .IN2(n3995), .IN3(s10_msel_gnt_p0[2]), .QN(
        n10069) );
  NAND3X0 U36248 ( .IN1(n3589), .IN2(n3590), .IN3(s1_msel_gnt_p0_2_), .QN(
        n11927) );
  NAND3X0 U36249 ( .IN1(n3544), .IN2(n3545), .IN3(s0_msel_gnt_p0[2]), .QN(
        n11617) );
  NAND3X0 U36250 ( .IN1(n3904), .IN2(n3905), .IN3(s8_msel_gnt_p0_2_), .QN(
        n9448) );
  NAND3X0 U36251 ( .IN1(n4219), .IN2(n4220), .IN3(test_so98), .QN(n14046) );
  NAND3X0 U36252 ( .IN1(n3867), .IN2(n3868), .IN3(s7_msel_gnt_p1[2]), .QN(
        n13844) );
  NAND3X0 U36253 ( .IN1(n3875), .IN2(n3876), .IN3(s7_msel_gnt_p2_2_), .QN(
        n13715) );
  NAND3X0 U36254 ( .IN1(n3822), .IN2(n3823), .IN3(test_so64), .QN(n13535) );
  NAND3X0 U36255 ( .IN1(n3830), .IN2(n3831), .IN3(s6_msel_gnt_p2[2]), .QN(
        n13406) );
  NAND3X0 U36256 ( .IN1(n4182), .IN2(n4183), .IN3(s14_msel_gnt_p1[2]), .QN(
        n11369) );
  NAND3X0 U36257 ( .IN1(n4190), .IN2(n4191), .IN3(s14_msel_gnt_p2_2_), .QN(
        n11240) );
  NAND3X0 U36258 ( .IN1(n3777), .IN2(n3778), .IN3(s5_msel_gnt_p1_2_), .QN(
        n13226) );
  NAND3X0 U36259 ( .IN1(n3785), .IN2(n3786), .IN3(s5_msel_gnt_p2[2]), .QN(
        n13097) );
  NAND3X0 U36260 ( .IN1(n3732), .IN2(n3733), .IN3(s4_msel_gnt_p1_2_), .QN(
        n12917) );
  NAND3X0 U36261 ( .IN1(n3740), .IN2(n3741), .IN3(s4_msel_gnt_p2[2]), .QN(
        n12788) );
  NAND3X0 U36262 ( .IN1(n4137), .IN2(n4138), .IN3(s13_msel_gnt_p1[2]), .QN(
        n11060) );
  NAND3X0 U36263 ( .IN1(n4145), .IN2(n4146), .IN3(s13_msel_gnt_p2_2_), .QN(
        n10931) );
  NAND3X0 U36264 ( .IN1(n4092), .IN2(n4093), .IN3(test_so87), .QN(n10750) );
  NAND3X0 U36265 ( .IN1(n4100), .IN2(n4101), .IN3(s12_msel_gnt_p2[2]), .QN(
        n10621) );
  NAND3X0 U36266 ( .IN1(n3687), .IN2(n3688), .IN3(s3_msel_gnt_p1[2]), .QN(
        n12608) );
  NAND3X0 U36267 ( .IN1(n3695), .IN2(n3696), .IN3(test_so53), .QN(n12479) );
  NAND3X0 U36268 ( .IN1(n3642), .IN2(n3643), .IN3(s2_msel_gnt_p1[2]), .QN(
        n12299) );
  NAND3X0 U36269 ( .IN1(n3650), .IN2(n3651), .IN3(s2_msel_gnt_p2_2_), .QN(
        n12170) );
  NAND3X0 U36270 ( .IN1(n4047), .IN2(n4048), .IN3(s11_msel_gnt_p1_2_), .QN(
        n10441) );
  NAND3X0 U36271 ( .IN1(n4055), .IN2(n4056), .IN3(s11_msel_gnt_p2[2]), .QN(
        n10312) );
  NAND3X0 U36272 ( .IN1(n4002), .IN2(n4003), .IN3(s10_msel_gnt_p1_2_), .QN(
        n10131) );
  NAND3X0 U36273 ( .IN1(n4010), .IN2(n4011), .IN3(s10_msel_gnt_p2[2]), .QN(
        n10002) );
  NAND3X0 U36274 ( .IN1(n3597), .IN2(n3598), .IN3(s1_msel_gnt_p1[2]), .QN(
        n11989) );
  NAND3X0 U36275 ( .IN1(n3605), .IN2(n3606), .IN3(s1_msel_gnt_p2_2_), .QN(
        n11860) );
  NAND3X0 U36276 ( .IN1(n3552), .IN2(n3553), .IN3(test_so41), .QN(n11679) );
  NAND3X0 U36277 ( .IN1(n3560), .IN2(n3561), .IN3(s0_msel_gnt_p2[2]), .QN(
        n11550) );
  NAND3X0 U36278 ( .IN1(n3957), .IN2(n3958), .IN3(s9_msel_gnt_p1[2]), .QN(
        n9821) );
  NAND3X0 U36279 ( .IN1(n3965), .IN2(n3966), .IN3(test_so76), .QN(n9692) );
  NAND3X0 U36280 ( .IN1(n3912), .IN2(n3913), .IN3(s8_msel_gnt_p1[2]), .QN(
        n9510) );
  NAND3X0 U36281 ( .IN1(n3920), .IN2(n3921), .IN3(s8_msel_gnt_p2_2_), .QN(
        n9381) );
  NAND3X0 U36282 ( .IN1(n4227), .IN2(n4228), .IN3(s15_msel_gnt_p1[2]), .QN(
        n13977) );
  NAND3X0 U36283 ( .IN1(n4235), .IN2(n4236), .IN3(test_so99), .QN(n14117) );
  NAND3X0 U36284 ( .IN1(n3883), .IN2(n3884), .IN3(s7_msel_gnt_p3[2]), .QN(
        n13911) );
  NAND3X0 U36285 ( .IN1(n3838), .IN2(n3839), .IN3(test_so65), .QN(n13602) );
  NAND3X0 U36286 ( .IN1(n4198), .IN2(n4199), .IN3(s14_msel_gnt_p3[2]), .QN(
        n11436) );
  NAND3X0 U36287 ( .IN1(n3793), .IN2(n3794), .IN3(s5_msel_gnt_p3_2_), .QN(
        n13293) );
  NAND3X0 U36288 ( .IN1(n3748), .IN2(n3749), .IN3(s4_msel_gnt_p3_2_), .QN(
        n12984) );
  NAND3X0 U36289 ( .IN1(n4153), .IN2(n4154), .IN3(s13_msel_gnt_p3[2]), .QN(
        n11127) );
  NAND3X0 U36290 ( .IN1(n4108), .IN2(n4109), .IN3(test_so88), .QN(n10817) );
  NAND3X0 U36291 ( .IN1(n3703), .IN2(n3704), .IN3(s3_msel_gnt_p3[2]), .QN(
        n12675) );
  NAND3X0 U36292 ( .IN1(n3658), .IN2(n3659), .IN3(s2_msel_gnt_p3[2]), .QN(
        n12366) );
  NAND3X0 U36293 ( .IN1(n4063), .IN2(n4064), .IN3(s11_msel_gnt_p3_2_), .QN(
        n10508) );
  NAND3X0 U36294 ( .IN1(n4018), .IN2(n4019), .IN3(s10_msel_gnt_p3_2_), .QN(
        n10198) );
  NAND3X0 U36295 ( .IN1(n3613), .IN2(n3614), .IN3(s1_msel_gnt_p3[2]), .QN(
        n12056) );
  NAND3X0 U36296 ( .IN1(n3568), .IN2(n3569), .IN3(test_so42), .QN(n11746) );
  NAND3X0 U36297 ( .IN1(n3973), .IN2(n3974), .IN3(s9_msel_gnt_p3[2]), .QN(
        n9888) );
  NAND3X0 U36298 ( .IN1(n3928), .IN2(n3929), .IN3(s8_msel_gnt_p3[2]), .QN(
        n9577) );
  NAND3X0 U36299 ( .IN1(n4243), .IN2(n4244), .IN3(s15_msel_gnt_p3[2]), .QN(
        n14185) );
  NAND3X0 U36300 ( .IN1(s7_msel_gnt_p3[2]), .IN2(n3883), .IN3(
        s7_msel_gnt_p3[1]), .QN(n13917) );
  NAND3X0 U36301 ( .IN1(s7_msel_gnt_p2_2_), .IN2(n3875), .IN3(
        s7_msel_gnt_p2_1_), .QN(n13720) );
  NAND3X0 U36302 ( .IN1(test_so65), .IN2(n3838), .IN3(s6_msel_gnt_p3_1_), .QN(
        n13608) );
  NAND3X0 U36303 ( .IN1(s6_msel_gnt_p2[2]), .IN2(n3830), .IN3(
        s6_msel_gnt_p2[1]), .QN(n13411) );
  NAND3X0 U36304 ( .IN1(s14_msel_gnt_p3[2]), .IN2(n4198), .IN3(
        s14_msel_gnt_p3[1]), .QN(n11442) );
  NAND3X0 U36305 ( .IN1(s14_msel_gnt_p2_2_), .IN2(n4190), .IN3(test_so95), 
        .QN(n11245) );
  NAND3X0 U36306 ( .IN1(s5_msel_gnt_p3_2_), .IN2(n3793), .IN3(test_so61), .QN(
        n13299) );
  NAND3X0 U36307 ( .IN1(s5_msel_gnt_p2[2]), .IN2(n3785), .IN3(
        s5_msel_gnt_p2[1]), .QN(n13102) );
  NAND3X0 U36308 ( .IN1(s4_msel_gnt_p3_2_), .IN2(n3748), .IN3(
        s4_msel_gnt_p3_1_), .QN(n12990) );
  NAND3X0 U36309 ( .IN1(s4_msel_gnt_p2[2]), .IN2(n3740), .IN3(
        s4_msel_gnt_p2[1]), .QN(n12793) );
  NAND3X0 U36310 ( .IN1(s13_msel_gnt_p3[2]), .IN2(n4153), .IN3(
        s13_msel_gnt_p3[1]), .QN(n11133) );
  NAND3X0 U36311 ( .IN1(s13_msel_gnt_p2_2_), .IN2(n4145), .IN3(
        s13_msel_gnt_p2_1_), .QN(n10936) );
  NAND3X0 U36312 ( .IN1(test_so88), .IN2(n4108), .IN3(s12_msel_gnt_p3_1_), 
        .QN(n10823) );
  NAND3X0 U36313 ( .IN1(s12_msel_gnt_p2[2]), .IN2(n4100), .IN3(
        s12_msel_gnt_p2[1]), .QN(n10626) );
  NAND3X0 U36314 ( .IN1(s3_msel_gnt_p3[2]), .IN2(n3703), .IN3(
        s3_msel_gnt_p3[1]), .QN(n12681) );
  NAND3X0 U36315 ( .IN1(test_so53), .IN2(n3695), .IN3(s3_msel_gnt_p2_1_), .QN(
        n12484) );
  NAND3X0 U36316 ( .IN1(s2_msel_gnt_p3[2]), .IN2(n3658), .IN3(
        s2_msel_gnt_p3[1]), .QN(n12372) );
  NAND3X0 U36317 ( .IN1(s2_msel_gnt_p2_2_), .IN2(n3650), .IN3(test_so49), .QN(
        n12175) );
  NAND3X0 U36318 ( .IN1(s11_msel_gnt_p3_2_), .IN2(n4063), .IN3(test_so84), 
        .QN(n10514) );
  NAND3X0 U36319 ( .IN1(s11_msel_gnt_p2[2]), .IN2(n4055), .IN3(
        s11_msel_gnt_p2[1]), .QN(n10317) );
  NAND3X0 U36320 ( .IN1(s10_msel_gnt_p3_2_), .IN2(n4018), .IN3(
        s10_msel_gnt_p3_1_), .QN(n10204) );
  NAND3X0 U36321 ( .IN1(s10_msel_gnt_p2[2]), .IN2(n4010), .IN3(
        s10_msel_gnt_p2[1]), .QN(n10007) );
  NAND3X0 U36322 ( .IN1(s1_msel_gnt_p3[2]), .IN2(n3613), .IN3(
        s1_msel_gnt_p3[1]), .QN(n12062) );
  NAND3X0 U36323 ( .IN1(s1_msel_gnt_p2_2_), .IN2(n3605), .IN3(
        s1_msel_gnt_p2_1_), .QN(n11865) );
  NAND3X0 U36324 ( .IN1(test_so42), .IN2(n3568), .IN3(s0_msel_gnt_p3_1_), .QN(
        n11752) );
  NAND3X0 U36325 ( .IN1(s0_msel_gnt_p2[2]), .IN2(n3560), .IN3(
        s0_msel_gnt_p2[1]), .QN(n11555) );
  NAND3X0 U36326 ( .IN1(s9_msel_gnt_p3[2]), .IN2(n3973), .IN3(
        s9_msel_gnt_p3[1]), .QN(n9894) );
  NAND3X0 U36327 ( .IN1(test_so76), .IN2(n3965), .IN3(s9_msel_gnt_p2_1_), .QN(
        n9697) );
  NAND3X0 U36328 ( .IN1(s8_msel_gnt_p3[2]), .IN2(n3928), .IN3(
        s8_msel_gnt_p3[1]), .QN(n9583) );
  NAND3X0 U36329 ( .IN1(s8_msel_gnt_p2_2_), .IN2(n3920), .IN3(test_so72), .QN(
        n9386) );
  NAND3X0 U36330 ( .IN1(s15_msel_gnt_p3[2]), .IN2(n4243), .IN3(
        s15_msel_gnt_p3[1]), .QN(n14191) );
  NAND3X0 U36331 ( .IN1(test_so99), .IN2(n4235), .IN3(s15_msel_gnt_p2_1_), 
        .QN(n14123) );
  NAND3X0 U36332 ( .IN1(s7_msel_gnt_p1[2]), .IN2(n3867), .IN3(
        s7_msel_gnt_p1[1]), .QN(n13850) );
  NAND3X0 U36333 ( .IN1(test_so64), .IN2(n3822), .IN3(s6_msel_gnt_p1_1_), .QN(
        n13541) );
  NAND3X0 U36334 ( .IN1(s14_msel_gnt_p1[2]), .IN2(n4182), .IN3(
        s14_msel_gnt_p1[1]), .QN(n11375) );
  NAND3X0 U36335 ( .IN1(s5_msel_gnt_p1_2_), .IN2(n3777), .IN3(test_so60), .QN(
        n13232) );
  NAND3X0 U36336 ( .IN1(s4_msel_gnt_p1_2_), .IN2(n3732), .IN3(
        s4_msel_gnt_p1_1_), .QN(n12923) );
  NAND3X0 U36337 ( .IN1(s13_msel_gnt_p1[2]), .IN2(n4137), .IN3(
        s13_msel_gnt_p1[1]), .QN(n11066) );
  NAND3X0 U36338 ( .IN1(test_so87), .IN2(n4092), .IN3(s12_msel_gnt_p1_1_), 
        .QN(n10756) );
  NAND3X0 U36339 ( .IN1(s3_msel_gnt_p1[2]), .IN2(n3687), .IN3(
        s3_msel_gnt_p1[1]), .QN(n12614) );
  NAND3X0 U36340 ( .IN1(s2_msel_gnt_p1[2]), .IN2(n3642), .IN3(
        s2_msel_gnt_p1[1]), .QN(n12305) );
  NAND3X0 U36341 ( .IN1(s11_msel_gnt_p1_2_), .IN2(n4047), .IN3(test_so83), 
        .QN(n10447) );
  NAND3X0 U36342 ( .IN1(s10_msel_gnt_p1_2_), .IN2(n4002), .IN3(
        s10_msel_gnt_p1_1_), .QN(n10137) );
  NAND3X0 U36343 ( .IN1(s1_msel_gnt_p1[2]), .IN2(n3597), .IN3(
        s1_msel_gnt_p1[1]), .QN(n11995) );
  NAND3X0 U36344 ( .IN1(test_so41), .IN2(n3552), .IN3(s0_msel_gnt_p1_1_), .QN(
        n11685) );
  NAND3X0 U36345 ( .IN1(s9_msel_gnt_p1[2]), .IN2(n3957), .IN3(
        s9_msel_gnt_p1[1]), .QN(n9827) );
  NAND3X0 U36346 ( .IN1(s8_msel_gnt_p1[2]), .IN2(n3912), .IN3(
        s8_msel_gnt_p1[1]), .QN(n9516) );
  NAND3X0 U36347 ( .IN1(s15_msel_gnt_p1[2]), .IN2(n4227), .IN3(
        s15_msel_gnt_p1[1]), .QN(n13983) );
  INVX0 U36348 ( .IN(m7_data_i[0]), .QN(n2257) );
  INVX0 U36349 ( .IN(m7_data_i[1]), .QN(n2256) );
  INVX0 U36350 ( .IN(m7_data_i[2]), .QN(n2255) );
  INVX0 U36351 ( .IN(m7_data_i[3]), .QN(n2254) );
  INVX0 U36352 ( .IN(m7_data_i[4]), .QN(n2253) );
  INVX0 U36353 ( .IN(m7_data_i[5]), .QN(n2252) );
  INVX0 U36354 ( .IN(m7_data_i[6]), .QN(n2251) );
  INVX0 U36355 ( .IN(m7_data_i[7]), .QN(n2250) );
  INVX0 U36356 ( .IN(m7_data_i[8]), .QN(n2249) );
  INVX0 U36357 ( .IN(m7_data_i[9]), .QN(n2248) );
  INVX0 U36358 ( .IN(m7_data_i[10]), .QN(n2247) );
  INVX0 U36359 ( .IN(m7_data_i[11]), .QN(n2246) );
  INVX0 U36360 ( .IN(m7_data_i[12]), .QN(n2245) );
  INVX0 U36361 ( .IN(m7_data_i[13]), .QN(n2244) );
  INVX0 U36362 ( .IN(m7_data_i[14]), .QN(n2243) );
  INVX0 U36363 ( .IN(m7_data_i[15]), .QN(n2242) );
  INVX0 U36364 ( .IN(m7_we_i), .QN(n2310) );
  INVX0 U36365 ( .IN(m5_we_i), .QN(n2138) );
  INVX0 U36366 ( .IN(m3_we_i), .QN(n1966) );
  INVX0 U36367 ( .IN(m1_we_i), .QN(n1794) );
  INVX0 U36368 ( .IN(m7_sel_i[0]), .QN(n2309) );
  INVX0 U36369 ( .IN(m5_sel_i[0]), .QN(n2137) );
  INVX0 U36370 ( .IN(m3_sel_i[0]), .QN(n1965) );
  INVX0 U36371 ( .IN(m1_sel_i[0]), .QN(n1793) );
  INVX0 U36372 ( .IN(m7_sel_i[1]), .QN(n2308) );
  INVX0 U36373 ( .IN(m5_sel_i[1]), .QN(n2136) );
  INVX0 U36374 ( .IN(m3_sel_i[1]), .QN(n1964) );
  INVX0 U36375 ( .IN(m1_sel_i[1]), .QN(n1792) );
  INVX0 U36376 ( .IN(m7_sel_i[2]), .QN(n2307) );
  INVX0 U36377 ( .IN(m5_sel_i[2]), .QN(n2135) );
  INVX0 U36378 ( .IN(m3_sel_i[2]), .QN(n1963) );
  INVX0 U36379 ( .IN(m1_sel_i[2]), .QN(n1791) );
  INVX0 U36380 ( .IN(m7_sel_i[3]), .QN(n2306) );
  INVX0 U36381 ( .IN(m5_sel_i[3]), .QN(n2134) );
  INVX0 U36382 ( .IN(m3_sel_i[3]), .QN(n1962) );
  INVX0 U36383 ( .IN(m1_sel_i[3]), .QN(n1790) );
  INVX0 U36384 ( .IN(m7_addr_i[0]), .QN(n2305) );
  INVX0 U36385 ( .IN(m5_addr_i[0]), .QN(n2133) );
  INVX0 U36386 ( .IN(m3_addr_i[0]), .QN(n1961) );
  INVX0 U36387 ( .IN(m1_addr_i[0]), .QN(n1789) );
  INVX0 U36388 ( .IN(m7_addr_i[1]), .QN(n2304) );
  INVX0 U36389 ( .IN(m5_addr_i[1]), .QN(n2132) );
  INVX0 U36390 ( .IN(m3_addr_i[1]), .QN(n1960) );
  INVX0 U36391 ( .IN(m1_addr_i[1]), .QN(n1788) );
  INVX0 U36392 ( .IN(m7_addr_i[6]), .QN(n2299) );
  INVX0 U36393 ( .IN(m5_addr_i[6]), .QN(n2127) );
  INVX0 U36394 ( .IN(m3_addr_i[6]), .QN(n1955) );
  INVX0 U36395 ( .IN(m1_addr_i[6]), .QN(n1783) );
  INVX0 U36396 ( .IN(m7_addr_i[7]), .QN(n2298) );
  INVX0 U36397 ( .IN(m5_addr_i[7]), .QN(n2126) );
  INVX0 U36398 ( .IN(m3_addr_i[7]), .QN(n1954) );
  INVX0 U36399 ( .IN(m1_addr_i[7]), .QN(n1782) );
  INVX0 U36400 ( .IN(m7_addr_i[8]), .QN(n2297) );
  INVX0 U36401 ( .IN(m5_addr_i[8]), .QN(n2125) );
  INVX0 U36402 ( .IN(m3_addr_i[8]), .QN(n1953) );
  INVX0 U36403 ( .IN(m1_addr_i[8]), .QN(n1781) );
  INVX0 U36404 ( .IN(m7_addr_i[9]), .QN(n2296) );
  INVX0 U36405 ( .IN(m5_addr_i[9]), .QN(n2124) );
  INVX0 U36406 ( .IN(m3_addr_i[9]), .QN(n1952) );
  INVX0 U36407 ( .IN(m1_addr_i[9]), .QN(n1780) );
  INVX0 U36408 ( .IN(m7_addr_i[10]), .QN(n2295) );
  INVX0 U36409 ( .IN(m5_addr_i[10]), .QN(n2123) );
  INVX0 U36410 ( .IN(m3_addr_i[10]), .QN(n1951) );
  INVX0 U36411 ( .IN(m1_addr_i[10]), .QN(n1779) );
  INVX0 U36412 ( .IN(m7_addr_i[11]), .QN(n2294) );
  INVX0 U36413 ( .IN(m5_addr_i[11]), .QN(n2122) );
  INVX0 U36414 ( .IN(m3_addr_i[11]), .QN(n1950) );
  INVX0 U36415 ( .IN(m1_addr_i[11]), .QN(n1778) );
  INVX0 U36416 ( .IN(m7_addr_i[12]), .QN(n2293) );
  INVX0 U36417 ( .IN(m5_addr_i[12]), .QN(n2121) );
  INVX0 U36418 ( .IN(m3_addr_i[12]), .QN(n1949) );
  INVX0 U36419 ( .IN(m1_addr_i[12]), .QN(n1777) );
  INVX0 U36420 ( .IN(m7_addr_i[13]), .QN(n2292) );
  INVX0 U36421 ( .IN(m5_addr_i[13]), .QN(n2120) );
  INVX0 U36422 ( .IN(m3_addr_i[13]), .QN(n1948) );
  INVX0 U36423 ( .IN(m1_addr_i[13]), .QN(n1776) );
  INVX0 U36424 ( .IN(m7_addr_i[14]), .QN(n2291) );
  INVX0 U36425 ( .IN(m5_addr_i[14]), .QN(n2119) );
  INVX0 U36426 ( .IN(m3_addr_i[14]), .QN(n1947) );
  INVX0 U36427 ( .IN(m1_addr_i[14]), .QN(n1775) );
  INVX0 U36428 ( .IN(m7_addr_i[15]), .QN(n2290) );
  INVX0 U36429 ( .IN(m5_addr_i[15]), .QN(n2118) );
  INVX0 U36430 ( .IN(m3_addr_i[15]), .QN(n1946) );
  INVX0 U36431 ( .IN(m1_addr_i[15]), .QN(n1774) );
  INVX0 U36432 ( .IN(m7_addr_i[16]), .QN(n2289) );
  INVX0 U36433 ( .IN(m5_addr_i[16]), .QN(n2117) );
  INVX0 U36434 ( .IN(m3_addr_i[16]), .QN(n1945) );
  INVX0 U36435 ( .IN(m1_addr_i[16]), .QN(n1773) );
  INVX0 U36436 ( .IN(m7_addr_i[17]), .QN(n2288) );
  INVX0 U36437 ( .IN(m5_addr_i[17]), .QN(n2116) );
  INVX0 U36438 ( .IN(m3_addr_i[17]), .QN(n1944) );
  INVX0 U36439 ( .IN(m1_addr_i[17]), .QN(n1772) );
  INVX0 U36440 ( .IN(m7_addr_i[18]), .QN(n2287) );
  INVX0 U36441 ( .IN(m5_addr_i[18]), .QN(n2115) );
  INVX0 U36442 ( .IN(m3_addr_i[18]), .QN(n1943) );
  INVX0 U36443 ( .IN(m1_addr_i[18]), .QN(n1771) );
  INVX0 U36444 ( .IN(m7_addr_i[19]), .QN(n2286) );
  INVX0 U36445 ( .IN(m5_addr_i[19]), .QN(n2114) );
  INVX0 U36446 ( .IN(m3_addr_i[19]), .QN(n1942) );
  INVX0 U36447 ( .IN(m1_addr_i[19]), .QN(n1770) );
  INVX0 U36448 ( .IN(m7_addr_i[20]), .QN(n2285) );
  INVX0 U36449 ( .IN(m5_addr_i[20]), .QN(n2113) );
  INVX0 U36450 ( .IN(m3_addr_i[20]), .QN(n1941) );
  INVX0 U36451 ( .IN(m1_addr_i[20]), .QN(n1769) );
  INVX0 U36452 ( .IN(m7_addr_i[21]), .QN(n2284) );
  INVX0 U36453 ( .IN(m5_addr_i[21]), .QN(n2112) );
  INVX0 U36454 ( .IN(m3_addr_i[21]), .QN(n1940) );
  INVX0 U36455 ( .IN(m1_addr_i[21]), .QN(n1768) );
  INVX0 U36456 ( .IN(m7_addr_i[22]), .QN(n2283) );
  INVX0 U36457 ( .IN(m5_addr_i[22]), .QN(n2111) );
  INVX0 U36458 ( .IN(m3_addr_i[22]), .QN(n1939) );
  INVX0 U36459 ( .IN(m1_addr_i[22]), .QN(n1767) );
  INVX0 U36460 ( .IN(m7_addr_i[23]), .QN(n2282) );
  INVX0 U36461 ( .IN(m5_addr_i[23]), .QN(n2110) );
  INVX0 U36462 ( .IN(m3_addr_i[23]), .QN(n1938) );
  INVX0 U36463 ( .IN(m1_addr_i[23]), .QN(n1766) );
  INVX0 U36464 ( .IN(m5_data_i[0]), .QN(n2085) );
  INVX0 U36465 ( .IN(m3_data_i[0]), .QN(n1913) );
  INVX0 U36466 ( .IN(m1_data_i[0]), .QN(n1741) );
  INVX0 U36467 ( .IN(m5_data_i[1]), .QN(n2084) );
  INVX0 U36468 ( .IN(m3_data_i[1]), .QN(n1912) );
  INVX0 U36469 ( .IN(m1_data_i[1]), .QN(n1740) );
  INVX0 U36470 ( .IN(m5_data_i[2]), .QN(n2083) );
  INVX0 U36471 ( .IN(m3_data_i[2]), .QN(n1911) );
  INVX0 U36472 ( .IN(m1_data_i[2]), .QN(n1739) );
  INVX0 U36473 ( .IN(m5_data_i[3]), .QN(n2082) );
  INVX0 U36474 ( .IN(m3_data_i[3]), .QN(n1910) );
  INVX0 U36475 ( .IN(m1_data_i[3]), .QN(n1738) );
  INVX0 U36476 ( .IN(m5_data_i[4]), .QN(n2081) );
  INVX0 U36477 ( .IN(m3_data_i[4]), .QN(n1909) );
  INVX0 U36478 ( .IN(m1_data_i[4]), .QN(n1737) );
  INVX0 U36479 ( .IN(m5_data_i[5]), .QN(n2080) );
  INVX0 U36480 ( .IN(m3_data_i[5]), .QN(n1908) );
  INVX0 U36481 ( .IN(m1_data_i[5]), .QN(n1736) );
  INVX0 U36482 ( .IN(m5_data_i[6]), .QN(n2079) );
  INVX0 U36483 ( .IN(m3_data_i[6]), .QN(n1907) );
  INVX0 U36484 ( .IN(m1_data_i[6]), .QN(n1735) );
  INVX0 U36485 ( .IN(m5_data_i[7]), .QN(n2078) );
  INVX0 U36486 ( .IN(m3_data_i[7]), .QN(n1906) );
  INVX0 U36487 ( .IN(m1_data_i[7]), .QN(n1734) );
  INVX0 U36488 ( .IN(m5_data_i[8]), .QN(n2077) );
  INVX0 U36489 ( .IN(m3_data_i[8]), .QN(n1905) );
  INVX0 U36490 ( .IN(m1_data_i[8]), .QN(n1733) );
  INVX0 U36491 ( .IN(m5_data_i[9]), .QN(n2076) );
  INVX0 U36492 ( .IN(m3_data_i[9]), .QN(n1904) );
  INVX0 U36493 ( .IN(m1_data_i[9]), .QN(n1732) );
  INVX0 U36494 ( .IN(m5_data_i[10]), .QN(n2075) );
  INVX0 U36495 ( .IN(m3_data_i[10]), .QN(n1903) );
  INVX0 U36496 ( .IN(m1_data_i[10]), .QN(n1731) );
  INVX0 U36497 ( .IN(m5_data_i[11]), .QN(n2074) );
  INVX0 U36498 ( .IN(m3_data_i[11]), .QN(n1902) );
  INVX0 U36499 ( .IN(m1_data_i[11]), .QN(n1730) );
  INVX0 U36500 ( .IN(m5_data_i[12]), .QN(n2073) );
  INVX0 U36501 ( .IN(m3_data_i[12]), .QN(n1901) );
  INVX0 U36502 ( .IN(m1_data_i[12]), .QN(n1729) );
  INVX0 U36503 ( .IN(m5_data_i[13]), .QN(n2072) );
  INVX0 U36504 ( .IN(m3_data_i[13]), .QN(n1900) );
  INVX0 U36505 ( .IN(m1_data_i[13]), .QN(n1728) );
  INVX0 U36506 ( .IN(m5_data_i[14]), .QN(n2071) );
  INVX0 U36507 ( .IN(m3_data_i[14]), .QN(n1899) );
  INVX0 U36508 ( .IN(m1_data_i[14]), .QN(n1727) );
  INVX0 U36509 ( .IN(m5_data_i[15]), .QN(n2070) );
  INVX0 U36510 ( .IN(m3_data_i[15]), .QN(n1898) );
  INVX0 U36511 ( .IN(m1_data_i[15]), .QN(n1726) );
  INVX0 U36512 ( .IN(m7_data_i[16]), .QN(n2241) );
  INVX0 U36513 ( .IN(m5_data_i[16]), .QN(n2069) );
  INVX0 U36514 ( .IN(m3_data_i[16]), .QN(n1897) );
  INVX0 U36515 ( .IN(m1_data_i[16]), .QN(n1725) );
  INVX0 U36516 ( .IN(m7_data_i[17]), .QN(n2240) );
  INVX0 U36517 ( .IN(m5_data_i[17]), .QN(n2068) );
  INVX0 U36518 ( .IN(m3_data_i[17]), .QN(n1896) );
  INVX0 U36519 ( .IN(m1_data_i[17]), .QN(n1724) );
  INVX0 U36520 ( .IN(m7_data_i[18]), .QN(n2239) );
  INVX0 U36521 ( .IN(m5_data_i[18]), .QN(n2067) );
  INVX0 U36522 ( .IN(m3_data_i[18]), .QN(n1895) );
  INVX0 U36523 ( .IN(m1_data_i[18]), .QN(n1723) );
  INVX0 U36524 ( .IN(m7_data_i[19]), .QN(n2238) );
  INVX0 U36525 ( .IN(m5_data_i[19]), .QN(n2066) );
  INVX0 U36526 ( .IN(m3_data_i[19]), .QN(n1894) );
  INVX0 U36527 ( .IN(m1_data_i[19]), .QN(n1722) );
  INVX0 U36528 ( .IN(m7_data_i[20]), .QN(n2237) );
  INVX0 U36529 ( .IN(m5_data_i[20]), .QN(n2065) );
  INVX0 U36530 ( .IN(m3_data_i[20]), .QN(n1893) );
  INVX0 U36531 ( .IN(m1_data_i[20]), .QN(n1721) );
  INVX0 U36532 ( .IN(m7_data_i[21]), .QN(n2236) );
  INVX0 U36533 ( .IN(m5_data_i[21]), .QN(n2064) );
  INVX0 U36534 ( .IN(m3_data_i[21]), .QN(n1892) );
  INVX0 U36535 ( .IN(m1_data_i[21]), .QN(n1720) );
  INVX0 U36536 ( .IN(m7_data_i[22]), .QN(n2235) );
  INVX0 U36537 ( .IN(m5_data_i[22]), .QN(n2063) );
  INVX0 U36538 ( .IN(m3_data_i[22]), .QN(n1891) );
  INVX0 U36539 ( .IN(m1_data_i[22]), .QN(n1719) );
  INVX0 U36540 ( .IN(m7_data_i[23]), .QN(n2234) );
  INVX0 U36541 ( .IN(m5_data_i[23]), .QN(n2062) );
  INVX0 U36542 ( .IN(m3_data_i[23]), .QN(n1890) );
  INVX0 U36543 ( .IN(m1_data_i[23]), .QN(n1718) );
  INVX0 U36544 ( .IN(m7_data_i[24]), .QN(n2233) );
  INVX0 U36545 ( .IN(m5_data_i[24]), .QN(n2061) );
  INVX0 U36546 ( .IN(m3_data_i[24]), .QN(n1889) );
  INVX0 U36547 ( .IN(m1_data_i[24]), .QN(n1717) );
  INVX0 U36548 ( .IN(m7_data_i[25]), .QN(n2232) );
  INVX0 U36549 ( .IN(m5_data_i[25]), .QN(n2060) );
  INVX0 U36550 ( .IN(m3_data_i[25]), .QN(n1888) );
  INVX0 U36551 ( .IN(m1_data_i[25]), .QN(n1716) );
  INVX0 U36552 ( .IN(m7_data_i[26]), .QN(n2231) );
  INVX0 U36553 ( .IN(m5_data_i[26]), .QN(n2059) );
  INVX0 U36554 ( .IN(m3_data_i[26]), .QN(n1887) );
  INVX0 U36555 ( .IN(m1_data_i[26]), .QN(n1715) );
  INVX0 U36556 ( .IN(m7_data_i[27]), .QN(n2230) );
  INVX0 U36557 ( .IN(m5_data_i[27]), .QN(n2058) );
  INVX0 U36558 ( .IN(m3_data_i[27]), .QN(n1886) );
  INVX0 U36559 ( .IN(m1_data_i[27]), .QN(n1714) );
  INVX0 U36560 ( .IN(m7_data_i[28]), .QN(n2229) );
  INVX0 U36561 ( .IN(m5_data_i[28]), .QN(n2057) );
  INVX0 U36562 ( .IN(m3_data_i[28]), .QN(n1885) );
  INVX0 U36563 ( .IN(m1_data_i[28]), .QN(n1713) );
  INVX0 U36564 ( .IN(m7_data_i[29]), .QN(n2228) );
  INVX0 U36565 ( .IN(m5_data_i[29]), .QN(n2056) );
  INVX0 U36566 ( .IN(m3_data_i[29]), .QN(n1884) );
  INVX0 U36567 ( .IN(m1_data_i[29]), .QN(n1712) );
  INVX0 U36568 ( .IN(m7_data_i[30]), .QN(n2227) );
  INVX0 U36569 ( .IN(m5_data_i[30]), .QN(n2055) );
  INVX0 U36570 ( .IN(m3_data_i[30]), .QN(n1883) );
  INVX0 U36571 ( .IN(m1_data_i[30]), .QN(n1711) );
  INVX0 U36572 ( .IN(m7_data_i[31]), .QN(n2226) );
  INVX0 U36573 ( .IN(m5_data_i[31]), .QN(n2054) );
  INVX0 U36574 ( .IN(m3_data_i[31]), .QN(n1882) );
  INVX0 U36575 ( .IN(m1_data_i[31]), .QN(n1710) );
  ISOLANDX1 U36576 ( .D(m0s7_cyc), .ISO(n13652), .Q(n13676) );
  ISOLANDX1 U36577 ( .D(test_so17), .ISO(n13343), .Q(n13367) );
  ISOLANDX1 U36578 ( .D(m0s14_cyc), .ISO(n11177), .Q(n11201) );
  ISOLANDX1 U36579 ( .D(m0s5_cyc), .ISO(n13034), .Q(n13058) );
  ISOLANDX1 U36580 ( .D(m0s4_cyc), .ISO(n12725), .Q(n12749) );
  ISOLANDX1 U36581 ( .D(test_so18), .ISO(n10868), .Q(n10892) );
  ISOLANDX1 U36582 ( .D(m0s12_cyc), .ISO(n10558), .Q(n10582) );
  ISOLANDX1 U36583 ( .D(m0s3_cyc), .ISO(n12416), .Q(n12440) );
  ISOLANDX1 U36584 ( .D(m0s2_cyc), .ISO(n12107), .Q(n12131) );
  ISOLANDX1 U36585 ( .D(m0s11_cyc), .ISO(n10249), .Q(n10273) );
  ISOLANDX1 U36586 ( .D(m0s10_cyc), .ISO(n9939), .Q(n9963) );
  ISOLANDX1 U36587 ( .D(m0s1_cyc), .ISO(n11797), .Q(n11821) );
  ISOLANDX1 U36588 ( .D(m0s0_cyc), .ISO(n11487), .Q(n11511) );
  ISOLANDX1 U36589 ( .D(m0s9_cyc), .ISO(n9629), .Q(n9653) );
  ISOLANDX1 U36590 ( .D(m0s8_cyc), .ISO(n9318), .Q(n9342) );
  ISOLANDX1 U36591 ( .D(m7s7_cyc), .ISO(n13658), .Q(n13854) );
  ISOLANDX1 U36592 ( .D(m7s6_cyc), .ISO(n13349), .Q(n13545) );
  ISOLANDX1 U36593 ( .D(m7s14_cyc), .ISO(n11183), .Q(n11379) );
  ISOLANDX1 U36594 ( .D(test_so34), .ISO(n13040), .Q(n13236) );
  ISOLANDX1 U36595 ( .D(m7s4_cyc), .ISO(n12731), .Q(n12927) );
  ISOLANDX1 U36596 ( .D(m7s13_cyc), .ISO(n10874), .Q(n11070) );
  ISOLANDX1 U36597 ( .D(m7s12_cyc), .ISO(n10564), .Q(n10760) );
  ISOLANDX1 U36598 ( .D(m7s3_cyc), .ISO(n12422), .Q(n12618) );
  ISOLANDX1 U36599 ( .D(m7s2_cyc), .ISO(n12113), .Q(n12309) );
  ISOLANDX1 U36600 ( .D(test_so35), .ISO(n10255), .Q(n10451) );
  ISOLANDX1 U36601 ( .D(m7s10_cyc), .ISO(n9945), .Q(n10141) );
  ISOLANDX1 U36602 ( .D(m7s1_cyc), .ISO(n11803), .Q(n11999) );
  ISOLANDX1 U36603 ( .D(m7s0_cyc), .ISO(n11493), .Q(n11689) );
  ISOLANDX1 U36604 ( .D(m7s9_cyc), .ISO(n9635), .Q(n9831) );
  ISOLANDX1 U36605 ( .D(m7s8_cyc), .ISO(n9324), .Q(n9520) );
  ISOLANDX1 U36606 ( .D(m7s15_cyc), .ISO(n14280), .Q(n13987) );
  ISOLANDX1 U36607 ( .D(m7s7_cyc), .ISO(n13657), .Q(n13791) );
  ISOLANDX1 U36608 ( .D(m7s6_cyc), .ISO(n13348), .Q(n13482) );
  ISOLANDX1 U36609 ( .D(m7s14_cyc), .ISO(n11182), .Q(n11316) );
  ISOLANDX1 U36610 ( .D(test_so34), .ISO(n13039), .Q(n13173) );
  ISOLANDX1 U36611 ( .D(m7s4_cyc), .ISO(n12730), .Q(n12864) );
  ISOLANDX1 U36612 ( .D(m7s13_cyc), .ISO(n10873), .Q(n11007) );
  ISOLANDX1 U36613 ( .D(m7s12_cyc), .ISO(n10563), .Q(n10697) );
  ISOLANDX1 U36614 ( .D(m7s3_cyc), .ISO(n12421), .Q(n12555) );
  ISOLANDX1 U36615 ( .D(m7s2_cyc), .ISO(n12112), .Q(n12246) );
  ISOLANDX1 U36616 ( .D(test_so35), .ISO(n10254), .Q(n10388) );
  ISOLANDX1 U36617 ( .D(m7s10_cyc), .ISO(n9944), .Q(n10078) );
  ISOLANDX1 U36618 ( .D(m7s1_cyc), .ISO(n11802), .Q(n11936) );
  ISOLANDX1 U36619 ( .D(m7s0_cyc), .ISO(n11492), .Q(n11626) );
  ISOLANDX1 U36620 ( .D(m7s9_cyc), .ISO(n9634), .Q(n9768) );
  ISOLANDX1 U36621 ( .D(m7s8_cyc), .ISO(n9323), .Q(n9457) );
  ISOLANDX1 U36622 ( .D(m7s15_cyc), .ISO(n14069), .Q(n14055) );
  INVX0 U36623 ( .IN(m6_data_i[0]), .QN(n2171) );
  INVX0 U36624 ( .IN(m6_data_i[1]), .QN(n2170) );
  INVX0 U36625 ( .IN(m6_data_i[2]), .QN(n2169) );
  INVX0 U36626 ( .IN(m6_data_i[3]), .QN(n2168) );
  INVX0 U36627 ( .IN(m6_data_i[4]), .QN(n2167) );
  INVX0 U36628 ( .IN(m6_data_i[5]), .QN(n2166) );
  INVX0 U36629 ( .IN(m6_data_i[6]), .QN(n2165) );
  INVX0 U36630 ( .IN(m6_data_i[7]), .QN(n2164) );
  INVX0 U36631 ( .IN(m6_data_i[8]), .QN(n2163) );
  INVX0 U36632 ( .IN(m6_data_i[9]), .QN(n2162) );
  INVX0 U36633 ( .IN(m6_data_i[10]), .QN(n2161) );
  INVX0 U36634 ( .IN(m6_data_i[11]), .QN(n2160) );
  INVX0 U36635 ( .IN(m6_data_i[12]), .QN(n2159) );
  INVX0 U36636 ( .IN(m6_data_i[13]), .QN(n2158) );
  INVX0 U36637 ( .IN(m6_data_i[14]), .QN(n2157) );
  INVX0 U36638 ( .IN(m6_data_i[15]), .QN(n2156) );
  INVX0 U36639 ( .IN(m6_we_i), .QN(n2224) );
  INVX0 U36640 ( .IN(m4_we_i), .QN(n2052) );
  INVX0 U36641 ( .IN(m2_we_i), .QN(n1880) );
  INVX0 U36642 ( .IN(m0_we_i), .QN(n1708) );
  INVX0 U36643 ( .IN(m6_sel_i[0]), .QN(n2223) );
  INVX0 U36644 ( .IN(m4_sel_i[0]), .QN(n2051) );
  INVX0 U36645 ( .IN(m2_sel_i[0]), .QN(n1879) );
  INVX0 U36646 ( .IN(m0_sel_i[0]), .QN(n1707) );
  INVX0 U36647 ( .IN(m6_sel_i[1]), .QN(n2222) );
  INVX0 U36648 ( .IN(m4_sel_i[1]), .QN(n2050) );
  INVX0 U36649 ( .IN(m2_sel_i[1]), .QN(n1878) );
  INVX0 U36650 ( .IN(m0_sel_i[1]), .QN(n1706) );
  INVX0 U36651 ( .IN(m6_sel_i[2]), .QN(n2221) );
  INVX0 U36652 ( .IN(m4_sel_i[2]), .QN(n2049) );
  INVX0 U36653 ( .IN(m2_sel_i[2]), .QN(n1877) );
  INVX0 U36654 ( .IN(m0_sel_i[2]), .QN(n1705) );
  INVX0 U36655 ( .IN(m6_sel_i[3]), .QN(n2220) );
  INVX0 U36656 ( .IN(m4_sel_i[3]), .QN(n2048) );
  INVX0 U36657 ( .IN(m2_sel_i[3]), .QN(n1876) );
  INVX0 U36658 ( .IN(m0_sel_i[3]), .QN(n1704) );
  INVX0 U36659 ( .IN(m6_addr_i[0]), .QN(n2219) );
  INVX0 U36660 ( .IN(m4_addr_i[0]), .QN(n2047) );
  INVX0 U36661 ( .IN(m2_addr_i[0]), .QN(n1875) );
  INVX0 U36662 ( .IN(m0_addr_i[0]), .QN(n1703) );
  INVX0 U36663 ( .IN(m6_addr_i[1]), .QN(n2218) );
  INVX0 U36664 ( .IN(m4_addr_i[1]), .QN(n2046) );
  INVX0 U36665 ( .IN(m2_addr_i[1]), .QN(n1874) );
  INVX0 U36666 ( .IN(m0_addr_i[1]), .QN(n1702) );
  INVX0 U36667 ( .IN(m6_addr_i[6]), .QN(n2213) );
  INVX0 U36668 ( .IN(m4_addr_i[6]), .QN(n2041) );
  INVX0 U36669 ( .IN(m2_addr_i[6]), .QN(n1869) );
  INVX0 U36670 ( .IN(m0_addr_i[6]), .QN(n1679) );
  INVX0 U36671 ( .IN(m6_addr_i[7]), .QN(n2212) );
  INVX0 U36672 ( .IN(m4_addr_i[7]), .QN(n2040) );
  INVX0 U36673 ( .IN(m2_addr_i[7]), .QN(n1868) );
  INVX0 U36674 ( .IN(m0_addr_i[7]), .QN(n1678) );
  INVX0 U36675 ( .IN(m6_addr_i[8]), .QN(n2211) );
  INVX0 U36676 ( .IN(m4_addr_i[8]), .QN(n2039) );
  INVX0 U36677 ( .IN(m2_addr_i[8]), .QN(n1867) );
  INVX0 U36678 ( .IN(m0_addr_i[8]), .QN(n1677) );
  INVX0 U36679 ( .IN(m6_addr_i[9]), .QN(n2210) );
  INVX0 U36680 ( .IN(m4_addr_i[9]), .QN(n2038) );
  INVX0 U36681 ( .IN(m2_addr_i[9]), .QN(n1866) );
  INVX0 U36682 ( .IN(m0_addr_i[9]), .QN(n1676) );
  INVX0 U36683 ( .IN(m6_addr_i[10]), .QN(n2209) );
  INVX0 U36684 ( .IN(m4_addr_i[10]), .QN(n2037) );
  INVX0 U36685 ( .IN(m2_addr_i[10]), .QN(n1865) );
  INVX0 U36686 ( .IN(m0_addr_i[10]), .QN(n1675) );
  INVX0 U36687 ( .IN(m6_addr_i[11]), .QN(n2208) );
  INVX0 U36688 ( .IN(m4_addr_i[11]), .QN(n2036) );
  INVX0 U36689 ( .IN(m2_addr_i[11]), .QN(n1864) );
  INVX0 U36690 ( .IN(m0_addr_i[11]), .QN(n1674) );
  INVX0 U36691 ( .IN(m6_addr_i[12]), .QN(n2207) );
  INVX0 U36692 ( .IN(m4_addr_i[12]), .QN(n2035) );
  INVX0 U36693 ( .IN(m2_addr_i[12]), .QN(n1863) );
  INVX0 U36694 ( .IN(m0_addr_i[12]), .QN(n1673) );
  INVX0 U36695 ( .IN(m6_addr_i[13]), .QN(n2206) );
  INVX0 U36696 ( .IN(m4_addr_i[13]), .QN(n2034) );
  INVX0 U36697 ( .IN(m2_addr_i[13]), .QN(n1862) );
  INVX0 U36698 ( .IN(m0_addr_i[13]), .QN(n1672) );
  INVX0 U36699 ( .IN(m6_addr_i[14]), .QN(n2205) );
  INVX0 U36700 ( .IN(m4_addr_i[14]), .QN(n2033) );
  INVX0 U36701 ( .IN(m2_addr_i[14]), .QN(n1861) );
  INVX0 U36702 ( .IN(m0_addr_i[14]), .QN(n1671) );
  INVX0 U36703 ( .IN(m6_addr_i[15]), .QN(n2204) );
  INVX0 U36704 ( .IN(m4_addr_i[15]), .QN(n2032) );
  INVX0 U36705 ( .IN(m2_addr_i[15]), .QN(n1860) );
  INVX0 U36706 ( .IN(m0_addr_i[15]), .QN(n1670) );
  INVX0 U36707 ( .IN(m6_addr_i[16]), .QN(n2203) );
  INVX0 U36708 ( .IN(m4_addr_i[16]), .QN(n2031) );
  INVX0 U36709 ( .IN(m2_addr_i[16]), .QN(n1859) );
  INVX0 U36710 ( .IN(m0_addr_i[16]), .QN(n1669) );
  INVX0 U36711 ( .IN(m6_addr_i[17]), .QN(n2202) );
  INVX0 U36712 ( .IN(m4_addr_i[17]), .QN(n2030) );
  INVX0 U36713 ( .IN(m2_addr_i[17]), .QN(n1858) );
  INVX0 U36714 ( .IN(m0_addr_i[17]), .QN(n1668) );
  INVX0 U36715 ( .IN(m6_addr_i[18]), .QN(n2201) );
  INVX0 U36716 ( .IN(m4_addr_i[18]), .QN(n2029) );
  INVX0 U36717 ( .IN(m2_addr_i[18]), .QN(n1857) );
  INVX0 U36718 ( .IN(m0_addr_i[18]), .QN(n1667) );
  INVX0 U36719 ( .IN(m6_addr_i[19]), .QN(n2200) );
  INVX0 U36720 ( .IN(m4_addr_i[19]), .QN(n2028) );
  INVX0 U36721 ( .IN(m2_addr_i[19]), .QN(n1856) );
  INVX0 U36722 ( .IN(m0_addr_i[19]), .QN(n1666) );
  INVX0 U36723 ( .IN(m6_addr_i[20]), .QN(n2199) );
  INVX0 U36724 ( .IN(m4_addr_i[20]), .QN(n2027) );
  INVX0 U36725 ( .IN(m2_addr_i[20]), .QN(n1855) );
  INVX0 U36726 ( .IN(m0_addr_i[20]), .QN(n1665) );
  INVX0 U36727 ( .IN(m6_addr_i[21]), .QN(n2198) );
  INVX0 U36728 ( .IN(m4_addr_i[21]), .QN(n2026) );
  INVX0 U36729 ( .IN(m2_addr_i[21]), .QN(n1854) );
  INVX0 U36730 ( .IN(m0_addr_i[21]), .QN(n1664) );
  INVX0 U36731 ( .IN(m6_addr_i[22]), .QN(n2197) );
  INVX0 U36732 ( .IN(m4_addr_i[22]), .QN(n2025) );
  INVX0 U36733 ( .IN(m2_addr_i[22]), .QN(n1853) );
  INVX0 U36734 ( .IN(m0_addr_i[22]), .QN(n1663) );
  INVX0 U36735 ( .IN(m6_addr_i[23]), .QN(n2196) );
  INVX0 U36736 ( .IN(m4_addr_i[23]), .QN(n2024) );
  INVX0 U36737 ( .IN(m2_addr_i[23]), .QN(n1852) );
  INVX0 U36738 ( .IN(m0_addr_i[23]), .QN(n1662) );
  INVX0 U36739 ( .IN(m4_data_i[0]), .QN(n1999) );
  INVX0 U36740 ( .IN(m2_data_i[0]), .QN(n1827) );
  INVX0 U36741 ( .IN(m0_data_i[0]), .QN(n1636) );
  INVX0 U36742 ( .IN(m4_data_i[1]), .QN(n1998) );
  INVX0 U36743 ( .IN(m2_data_i[1]), .QN(n1826) );
  INVX0 U36744 ( .IN(m0_data_i[1]), .QN(n1635) );
  INVX0 U36745 ( .IN(m4_data_i[2]), .QN(n1997) );
  INVX0 U36746 ( .IN(m2_data_i[2]), .QN(n1825) );
  INVX0 U36747 ( .IN(m0_data_i[2]), .QN(n1634) );
  INVX0 U36748 ( .IN(m4_data_i[3]), .QN(n1996) );
  INVX0 U36749 ( .IN(m2_data_i[3]), .QN(n1824) );
  INVX0 U36750 ( .IN(m0_data_i[3]), .QN(n1633) );
  INVX0 U36751 ( .IN(m4_data_i[4]), .QN(n1995) );
  INVX0 U36752 ( .IN(m2_data_i[4]), .QN(n1823) );
  INVX0 U36753 ( .IN(m0_data_i[4]), .QN(n1632) );
  INVX0 U36754 ( .IN(m4_data_i[5]), .QN(n1994) );
  INVX0 U36755 ( .IN(m2_data_i[5]), .QN(n1822) );
  INVX0 U36756 ( .IN(m0_data_i[5]), .QN(n1631) );
  INVX0 U36757 ( .IN(m4_data_i[6]), .QN(n1993) );
  INVX0 U36758 ( .IN(m2_data_i[6]), .QN(n1821) );
  INVX0 U36759 ( .IN(m0_data_i[6]), .QN(n1630) );
  INVX0 U36760 ( .IN(m4_data_i[7]), .QN(n1992) );
  INVX0 U36761 ( .IN(m2_data_i[7]), .QN(n1820) );
  INVX0 U36762 ( .IN(m0_data_i[7]), .QN(n1629) );
  INVX0 U36763 ( .IN(m4_data_i[8]), .QN(n1991) );
  INVX0 U36764 ( .IN(m2_data_i[8]), .QN(n1819) );
  INVX0 U36765 ( .IN(m0_data_i[8]), .QN(n1628) );
  INVX0 U36766 ( .IN(m4_data_i[9]), .QN(n1990) );
  INVX0 U36767 ( .IN(m2_data_i[9]), .QN(n1818) );
  INVX0 U36768 ( .IN(m0_data_i[9]), .QN(n1627) );
  INVX0 U36769 ( .IN(m4_data_i[10]), .QN(n1989) );
  INVX0 U36770 ( .IN(m2_data_i[10]), .QN(n1817) );
  INVX0 U36771 ( .IN(m0_data_i[10]), .QN(n1626) );
  INVX0 U36772 ( .IN(m4_data_i[11]), .QN(n1988) );
  INVX0 U36773 ( .IN(m2_data_i[11]), .QN(n1816) );
  INVX0 U36774 ( .IN(m0_data_i[11]), .QN(n1625) );
  INVX0 U36775 ( .IN(m4_data_i[12]), .QN(n1987) );
  INVX0 U36776 ( .IN(m2_data_i[12]), .QN(n1815) );
  INVX0 U36777 ( .IN(m0_data_i[12]), .QN(n1624) );
  INVX0 U36778 ( .IN(m4_data_i[13]), .QN(n1986) );
  INVX0 U36779 ( .IN(m2_data_i[13]), .QN(n1814) );
  INVX0 U36780 ( .IN(m0_data_i[13]), .QN(n1623) );
  INVX0 U36781 ( .IN(m4_data_i[14]), .QN(n1985) );
  INVX0 U36782 ( .IN(m2_data_i[14]), .QN(n1813) );
  INVX0 U36783 ( .IN(m0_data_i[14]), .QN(n1622) );
  INVX0 U36784 ( .IN(m4_data_i[15]), .QN(n1984) );
  INVX0 U36785 ( .IN(m2_data_i[15]), .QN(n1812) );
  INVX0 U36786 ( .IN(m0_data_i[15]), .QN(n1621) );
  INVX0 U36787 ( .IN(m6_data_i[16]), .QN(n2155) );
  INVX0 U36788 ( .IN(m4_data_i[16]), .QN(n1983) );
  INVX0 U36789 ( .IN(m2_data_i[16]), .QN(n1811) );
  INVX0 U36790 ( .IN(m0_data_i[16]), .QN(n1620) );
  INVX0 U36791 ( .IN(m6_data_i[17]), .QN(n2154) );
  INVX0 U36792 ( .IN(m4_data_i[17]), .QN(n1982) );
  INVX0 U36793 ( .IN(m2_data_i[17]), .QN(n1810) );
  INVX0 U36794 ( .IN(m0_data_i[17]), .QN(n1619) );
  INVX0 U36795 ( .IN(m6_data_i[18]), .QN(n2153) );
  INVX0 U36796 ( .IN(m4_data_i[18]), .QN(n1981) );
  INVX0 U36797 ( .IN(m2_data_i[18]), .QN(n1809) );
  INVX0 U36798 ( .IN(m0_data_i[18]), .QN(n1618) );
  INVX0 U36799 ( .IN(m6_data_i[19]), .QN(n2152) );
  INVX0 U36800 ( .IN(m4_data_i[19]), .QN(n1980) );
  INVX0 U36801 ( .IN(m2_data_i[19]), .QN(n1808) );
  INVX0 U36802 ( .IN(m0_data_i[19]), .QN(n1617) );
  INVX0 U36803 ( .IN(m6_data_i[20]), .QN(n2151) );
  INVX0 U36804 ( .IN(m4_data_i[20]), .QN(n1979) );
  INVX0 U36805 ( .IN(m2_data_i[20]), .QN(n1807) );
  INVX0 U36806 ( .IN(m0_data_i[20]), .QN(n1616) );
  INVX0 U36807 ( .IN(m6_data_i[21]), .QN(n2150) );
  INVX0 U36808 ( .IN(m4_data_i[21]), .QN(n1978) );
  INVX0 U36809 ( .IN(m2_data_i[21]), .QN(n1806) );
  INVX0 U36810 ( .IN(m0_data_i[21]), .QN(n1615) );
  INVX0 U36811 ( .IN(m6_data_i[22]), .QN(n2149) );
  INVX0 U36812 ( .IN(m4_data_i[22]), .QN(n1977) );
  INVX0 U36813 ( .IN(m2_data_i[22]), .QN(n1805) );
  INVX0 U36814 ( .IN(m0_data_i[22]), .QN(n1614) );
  INVX0 U36815 ( .IN(m6_data_i[23]), .QN(n2148) );
  INVX0 U36816 ( .IN(m4_data_i[23]), .QN(n1976) );
  INVX0 U36817 ( .IN(m2_data_i[23]), .QN(n1804) );
  INVX0 U36818 ( .IN(m0_data_i[23]), .QN(n1613) );
  INVX0 U36819 ( .IN(m6_data_i[24]), .QN(n2147) );
  INVX0 U36820 ( .IN(m4_data_i[24]), .QN(n1975) );
  INVX0 U36821 ( .IN(m2_data_i[24]), .QN(n1803) );
  INVX0 U36822 ( .IN(m0_data_i[24]), .QN(n1612) );
  INVX0 U36823 ( .IN(m6_data_i[25]), .QN(n2146) );
  INVX0 U36824 ( .IN(m4_data_i[25]), .QN(n1974) );
  INVX0 U36825 ( .IN(m2_data_i[25]), .QN(n1802) );
  INVX0 U36826 ( .IN(m0_data_i[25]), .QN(n1611) );
  INVX0 U36827 ( .IN(m6_data_i[26]), .QN(n2145) );
  INVX0 U36828 ( .IN(m4_data_i[26]), .QN(n1973) );
  INVX0 U36829 ( .IN(m2_data_i[26]), .QN(n1801) );
  INVX0 U36830 ( .IN(m0_data_i[26]), .QN(n1610) );
  INVX0 U36831 ( .IN(m6_data_i[27]), .QN(n2144) );
  INVX0 U36832 ( .IN(m4_data_i[27]), .QN(n1972) );
  INVX0 U36833 ( .IN(m2_data_i[27]), .QN(n1800) );
  INVX0 U36834 ( .IN(m0_data_i[27]), .QN(n1609) );
  INVX0 U36835 ( .IN(m6_data_i[28]), .QN(n2143) );
  INVX0 U36836 ( .IN(m4_data_i[28]), .QN(n1971) );
  INVX0 U36837 ( .IN(m2_data_i[28]), .QN(n1799) );
  INVX0 U36838 ( .IN(m0_data_i[28]), .QN(n1608) );
  INVX0 U36839 ( .IN(m6_data_i[29]), .QN(n2142) );
  INVX0 U36840 ( .IN(m4_data_i[29]), .QN(n1970) );
  INVX0 U36841 ( .IN(m2_data_i[29]), .QN(n1798) );
  INVX0 U36842 ( .IN(m0_data_i[29]), .QN(n1607) );
  INVX0 U36843 ( .IN(m6_data_i[30]), .QN(n2141) );
  INVX0 U36844 ( .IN(m4_data_i[30]), .QN(n1969) );
  INVX0 U36845 ( .IN(m2_data_i[30]), .QN(n1797) );
  INVX0 U36846 ( .IN(m0_data_i[30]), .QN(n1606) );
  INVX0 U36847 ( .IN(m6_data_i[31]), .QN(n2140) );
  INVX0 U36848 ( .IN(m4_data_i[31]), .QN(n1968) );
  INVX0 U36849 ( .IN(m2_data_i[31]), .QN(n1796) );
  INVX0 U36850 ( .IN(m0_data_i[31]), .QN(n1605) );
  NAND3X0 U36851 ( .IN1(s7_msel_gnt_p2_2_), .IN2(n3876), .IN3(test_so68), .QN(
        n13732) );
  NAND3X0 U36852 ( .IN1(s6_msel_gnt_p2[2]), .IN2(n3831), .IN3(
        s6_msel_gnt_p2[0]), .QN(n13423) );
  NAND3X0 U36853 ( .IN1(s14_msel_gnt_p2_2_), .IN2(n4191), .IN3(
        s14_msel_gnt_p2_0_), .QN(n11257) );
  NAND3X0 U36854 ( .IN1(s5_msel_gnt_p2[2]), .IN2(n3786), .IN3(
        s5_msel_gnt_p2[0]), .QN(n13114) );
  NAND3X0 U36855 ( .IN1(s4_msel_gnt_p2[2]), .IN2(n3741), .IN3(
        s4_msel_gnt_p2[0]), .QN(n12805) );
  NAND3X0 U36856 ( .IN1(s13_msel_gnt_p2_2_), .IN2(n4146), .IN3(test_so91), 
        .QN(n10948) );
  NAND3X0 U36857 ( .IN1(s12_msel_gnt_p2[2]), .IN2(n4101), .IN3(
        s12_msel_gnt_p2[0]), .QN(n10638) );
  NAND3X0 U36858 ( .IN1(test_so53), .IN2(n3696), .IN3(s3_msel_gnt_p2_0_), .QN(
        n12496) );
  NAND3X0 U36859 ( .IN1(s2_msel_gnt_p2_2_), .IN2(n3651), .IN3(
        s2_msel_gnt_p2_0_), .QN(n12187) );
  NAND3X0 U36860 ( .IN1(s11_msel_gnt_p2[2]), .IN2(n4056), .IN3(
        s11_msel_gnt_p2[0]), .QN(n10329) );
  NAND3X0 U36861 ( .IN1(s10_msel_gnt_p2[2]), .IN2(n4011), .IN3(
        s10_msel_gnt_p2[0]), .QN(n10019) );
  NAND3X0 U36862 ( .IN1(s1_msel_gnt_p2_2_), .IN2(n3606), .IN3(test_so45), .QN(
        n11877) );
  NAND3X0 U36863 ( .IN1(s0_msel_gnt_p2[2]), .IN2(n3561), .IN3(
        s0_msel_gnt_p2[0]), .QN(n11567) );
  NAND3X0 U36864 ( .IN1(test_so76), .IN2(n3966), .IN3(s9_msel_gnt_p2_0_), .QN(
        n9709) );
  NAND3X0 U36865 ( .IN1(s8_msel_gnt_p2_2_), .IN2(n3921), .IN3(
        s8_msel_gnt_p2_0_), .QN(n9398) );
  NAND3X0 U36866 ( .IN1(test_so99), .IN2(n4236), .IN3(s15_msel_gnt_p2_0_), 
        .QN(n14136) );
  NAND3X0 U36867 ( .IN1(s7_msel_gnt_p3[2]), .IN2(n3884), .IN3(
        s7_msel_gnt_p3[0]), .QN(n13929) );
  NAND3X0 U36868 ( .IN1(test_so65), .IN2(n3839), .IN3(s6_msel_gnt_p3_0_), .QN(
        n13620) );
  NAND3X0 U36869 ( .IN1(s14_msel_gnt_p3[2]), .IN2(n4199), .IN3(
        s14_msel_gnt_p3[0]), .QN(n11454) );
  NAND3X0 U36870 ( .IN1(s5_msel_gnt_p3_2_), .IN2(n3794), .IN3(
        s5_msel_gnt_p3_0_), .QN(n13311) );
  NAND3X0 U36871 ( .IN1(s4_msel_gnt_p3_2_), .IN2(n3749), .IN3(test_so57), .QN(
        n13002) );
  NAND3X0 U36872 ( .IN1(s13_msel_gnt_p3[2]), .IN2(n4154), .IN3(
        s13_msel_gnt_p3[0]), .QN(n11145) );
  NAND3X0 U36873 ( .IN1(test_so88), .IN2(n4109), .IN3(s12_msel_gnt_p3_0_), 
        .QN(n10835) );
  NAND3X0 U36874 ( .IN1(s3_msel_gnt_p3[2]), .IN2(n3704), .IN3(
        s3_msel_gnt_p3[0]), .QN(n12693) );
  NAND3X0 U36875 ( .IN1(s2_msel_gnt_p3[2]), .IN2(n3659), .IN3(
        s2_msel_gnt_p3[0]), .QN(n12384) );
  NAND3X0 U36876 ( .IN1(s11_msel_gnt_p3_2_), .IN2(n4064), .IN3(
        s11_msel_gnt_p3_0_), .QN(n10526) );
  NAND3X0 U36877 ( .IN1(s10_msel_gnt_p3_2_), .IN2(n4019), .IN3(test_so80), 
        .QN(n10216) );
  NAND3X0 U36878 ( .IN1(s1_msel_gnt_p3[2]), .IN2(n3614), .IN3(
        s1_msel_gnt_p3[0]), .QN(n12074) );
  NAND3X0 U36879 ( .IN1(test_so42), .IN2(n3569), .IN3(s0_msel_gnt_p3_0_), .QN(
        n11764) );
  NAND3X0 U36880 ( .IN1(s9_msel_gnt_p3[2]), .IN2(n3974), .IN3(
        s9_msel_gnt_p3[0]), .QN(n9906) );
  NAND3X0 U36881 ( .IN1(s8_msel_gnt_p3[2]), .IN2(n3929), .IN3(
        s8_msel_gnt_p3[0]), .QN(n9595) );
  NAND3X0 U36882 ( .IN1(s15_msel_gnt_p3[2]), .IN2(n4244), .IN3(
        s15_msel_gnt_p3[0]), .QN(n14203) );
  NAND3X0 U36883 ( .IN1(s7_msel_gnt_p1[2]), .IN2(n3868), .IN3(
        s7_msel_gnt_p1[0]), .QN(n13863) );
  NAND3X0 U36884 ( .IN1(test_so64), .IN2(n3823), .IN3(s6_msel_gnt_p1_0_), .QN(
        n13554) );
  NAND3X0 U36885 ( .IN1(s14_msel_gnt_p1[2]), .IN2(n4183), .IN3(
        s14_msel_gnt_p1[0]), .QN(n11388) );
  NAND3X0 U36886 ( .IN1(s5_msel_gnt_p1_2_), .IN2(n3778), .IN3(
        s5_msel_gnt_p1_0_), .QN(n13245) );
  NAND3X0 U36887 ( .IN1(s4_msel_gnt_p1_2_), .IN2(n3733), .IN3(test_so56), .QN(
        n12936) );
  NAND3X0 U36888 ( .IN1(s13_msel_gnt_p1[2]), .IN2(n4138), .IN3(
        s13_msel_gnt_p1[0]), .QN(n11079) );
  NAND3X0 U36889 ( .IN1(test_so87), .IN2(n4093), .IN3(s12_msel_gnt_p1_0_), 
        .QN(n10769) );
  NAND3X0 U36890 ( .IN1(s3_msel_gnt_p1[2]), .IN2(n3688), .IN3(
        s3_msel_gnt_p1[0]), .QN(n12627) );
  NAND3X0 U36891 ( .IN1(s2_msel_gnt_p1[2]), .IN2(n3643), .IN3(
        s2_msel_gnt_p1[0]), .QN(n12318) );
  NAND3X0 U36892 ( .IN1(s11_msel_gnt_p1_2_), .IN2(n4048), .IN3(
        s11_msel_gnt_p1_0_), .QN(n10460) );
  NAND3X0 U36893 ( .IN1(s10_msel_gnt_p1_2_), .IN2(n4003), .IN3(test_so79), 
        .QN(n10150) );
  NAND3X0 U36894 ( .IN1(s1_msel_gnt_p1[2]), .IN2(n3598), .IN3(
        s1_msel_gnt_p1[0]), .QN(n12008) );
  NAND3X0 U36895 ( .IN1(test_so41), .IN2(n3553), .IN3(s0_msel_gnt_p1_0_), .QN(
        n11698) );
  NAND3X0 U36896 ( .IN1(s9_msel_gnt_p1[2]), .IN2(n3958), .IN3(
        s9_msel_gnt_p1[0]), .QN(n9840) );
  NAND3X0 U36897 ( .IN1(s8_msel_gnt_p1[2]), .IN2(n3913), .IN3(
        s8_msel_gnt_p1[0]), .QN(n9529) );
  NAND3X0 U36898 ( .IN1(s15_msel_gnt_p1[2]), .IN2(n4228), .IN3(
        s15_msel_gnt_p1[0]), .QN(n13996) );
  ISOLANDX1 U36899 ( .D(m0s7_cyc), .ISO(n13651), .Q(n13847) );
  ISOLANDX1 U36900 ( .D(test_so17), .ISO(n13342), .Q(n13538) );
  ISOLANDX1 U36901 ( .D(m0s14_cyc), .ISO(n11176), .Q(n11372) );
  ISOLANDX1 U36902 ( .D(m0s5_cyc), .ISO(n13033), .Q(n13229) );
  ISOLANDX1 U36903 ( .D(m0s4_cyc), .ISO(n12724), .Q(n12920) );
  ISOLANDX1 U36904 ( .D(test_so18), .ISO(n10867), .Q(n11063) );
  ISOLANDX1 U36905 ( .D(m0s12_cyc), .ISO(n10557), .Q(n10753) );
  ISOLANDX1 U36906 ( .D(m0s3_cyc), .ISO(n12415), .Q(n12611) );
  ISOLANDX1 U36907 ( .D(m0s2_cyc), .ISO(n12106), .Q(n12302) );
  ISOLANDX1 U36908 ( .D(m0s11_cyc), .ISO(n10248), .Q(n10444) );
  ISOLANDX1 U36909 ( .D(m0s10_cyc), .ISO(n9938), .Q(n10134) );
  ISOLANDX1 U36910 ( .D(m0s1_cyc), .ISO(n11796), .Q(n11992) );
  ISOLANDX1 U36911 ( .D(m0s0_cyc), .ISO(n11486), .Q(n11682) );
  ISOLANDX1 U36912 ( .D(m0s9_cyc), .ISO(n9628), .Q(n9824) );
  ISOLANDX1 U36913 ( .D(m0s8_cyc), .ISO(n9317), .Q(n9513) );
  ISOLANDX1 U36914 ( .D(m0s15_cyc), .ISO(n14281), .Q(n13980) );
  AO22X1 U36915 ( .IN1(n14324), .IN2(m7s0_cyc), .IN3(n14325), .IN4(n18769), 
        .Q(n17636) );
  AO22X1 U36916 ( .IN1(n14324), .IN2(m7s1_cyc), .IN3(n14325), .IN4(n17824), 
        .Q(n17637) );
  AO22X1 U36917 ( .IN1(n14324), .IN2(m7s2_cyc), .IN3(n14325), .IN4(n17794), 
        .Q(n17638) );
  AO22X1 U36918 ( .IN1(n14324), .IN2(m7s3_cyc), .IN3(n14325), .IN4(n17793), 
        .Q(n17639) );
  AO22X1 U36919 ( .IN1(n14324), .IN2(m7s4_cyc), .IN3(n14325), .IN4(n17796), 
        .Q(n17640) );
  AO22X1 U36920 ( .IN1(n14324), .IN2(test_so34), .IN3(n14325), .IN4(n17795), 
        .Q(n17641) );
  AO22X1 U36921 ( .IN1(n14324), .IN2(m7s6_cyc), .IN3(n14325), .IN4(n17869), 
        .Q(n17642) );
  AO22X1 U36922 ( .IN1(n14324), .IN2(m7s7_cyc), .IN3(n14325), .IN4(n17882), 
        .Q(n17643) );
  AO22X1 U36923 ( .IN1(n14324), .IN2(m7s8_cyc), .IN3(n14325), .IN4(n17830), 
        .Q(n17644) );
  AO22X1 U36924 ( .IN1(n14324), .IN2(m7s9_cyc), .IN3(n14325), .IN4(n17873), 
        .Q(n17645) );
  AO22X1 U36925 ( .IN1(n14324), .IN2(m7s10_cyc), .IN3(n14325), .IN4(n18793), 
        .Q(n17646) );
  AO22X1 U36926 ( .IN1(n14324), .IN2(test_so35), .IN3(n14325), .IN4(n17820), 
        .Q(n17647) );
  AO22X1 U36927 ( .IN1(n14324), .IN2(m7s12_cyc), .IN3(n14325), .IN4(n17809), 
        .Q(n17648) );
  AO22X1 U36928 ( .IN1(n14324), .IN2(m7s13_cyc), .IN3(n14325), .IN4(n17810), 
        .Q(n17649) );
  AO22X1 U36929 ( .IN1(n14324), .IN2(m7s14_cyc), .IN3(n14325), .IN4(n17817), 
        .Q(n17650) );
  AO22X1 U36930 ( .IN1(n14324), .IN2(m7s15_cyc), .IN3(n14325), .IN4(n17781), 
        .Q(n17651) );
  AO22X1 U36931 ( .IN1(n14326), .IN2(m6s0_cyc), .IN3(n14327), .IN4(n18721), 
        .Q(n17652) );
  AO22X1 U36932 ( .IN1(n14326), .IN2(m6s1_cyc), .IN3(n14327), .IN4(n17859), 
        .Q(n17653) );
  AO22X1 U36933 ( .IN1(n14326), .IN2(m6s2_cyc), .IN3(n14327), .IN4(n17834), 
        .Q(n17654) );
  AO22X1 U36934 ( .IN1(n14326), .IN2(test_so31), .IN3(n14327), .IN4(n18727), 
        .Q(n17655) );
  AO22X1 U36935 ( .IN1(n14326), .IN2(m6s4_cyc), .IN3(n14327), .IN4(n17836), 
        .Q(n17656) );
  AO22X1 U36936 ( .IN1(n14326), .IN2(m6s5_cyc), .IN3(n14327), .IN4(n17835), 
        .Q(n17657) );
  AO22X1 U36937 ( .IN1(n14326), .IN2(m6s6_cyc), .IN3(n14327), .IN4(n18733), 
        .Q(n17658) );
  AO22X1 U36938 ( .IN1(n14326), .IN2(m6s7_cyc), .IN3(n14327), .IN4(n17858), 
        .Q(n17659) );
  AO22X1 U36939 ( .IN1(n14326), .IN2(m6s8_cyc), .IN3(n14327), .IN4(n17865), 
        .Q(n17660) );
  AO22X1 U36940 ( .IN1(n14326), .IN2(test_so32), .IN3(n14327), .IN4(n17877), 
        .Q(n17661) );
  AO22X1 U36941 ( .IN1(n14326), .IN2(m6s10_cyc), .IN3(n14327), .IN4(n18745), 
        .Q(n17662) );
  AO22X1 U36942 ( .IN1(n14326), .IN2(m6s11_cyc), .IN3(n14327), .IN4(n17850), 
        .Q(n17663) );
  AO22X1 U36943 ( .IN1(n14326), .IN2(m6s12_cyc), .IN3(n14327), .IN4(n18757), 
        .Q(n17664) );
  AO22X1 U36944 ( .IN1(n14326), .IN2(m6s13_cyc), .IN3(n14327), .IN4(n17846), 
        .Q(n17665) );
  AO22X1 U36945 ( .IN1(n14326), .IN2(m6s14_cyc), .IN3(n14327), .IN4(n17854), 
        .Q(n17666) );
  AO22X1 U36946 ( .IN1(n14326), .IN2(test_so33), .IN3(n14327), .IN4(n17785), 
        .Q(n17667) );
  AO22X1 U36947 ( .IN1(n14332), .IN2(test_so23), .IN3(n14333), .IN4(n18577), 
        .Q(n17700) );
  AO22X1 U36948 ( .IN1(n14332), .IN2(m3s1_cyc), .IN3(n14333), .IN4(n17825), 
        .Q(n17701) );
  AO22X1 U36949 ( .IN1(n14332), .IN2(m3s2_cyc), .IN3(n14333), .IN4(n17802), 
        .Q(n17702) );
  AO22X1 U36950 ( .IN1(n14332), .IN2(m3s3_cyc), .IN3(n14333), .IN4(n17801), 
        .Q(n17703) );
  AO22X1 U36951 ( .IN1(n14332), .IN2(m3s4_cyc), .IN3(n14333), .IN4(n17804), 
        .Q(n17704) );
  AO22X1 U36952 ( .IN1(n14332), .IN2(m3s5_cyc), .IN3(n14333), .IN4(n17803), 
        .Q(n17705) );
  AO22X1 U36953 ( .IN1(n14332), .IN2(m3s6_cyc), .IN3(n14333), .IN4(n17870), 
        .Q(n17706) );
  AO22X1 U36954 ( .IN1(n14332), .IN2(test_so24), .IN3(n14333), .IN4(n17883), 
        .Q(n17707) );
  AO22X1 U36955 ( .IN1(n14332), .IN2(m3s8_cyc), .IN3(n14333), .IN4(n17832), 
        .Q(n17708) );
  AO22X1 U36956 ( .IN1(n14332), .IN2(m3s9_cyc), .IN3(n14333), .IN4(n17875), 
        .Q(n17709) );
  AO22X1 U36957 ( .IN1(n14332), .IN2(m3s10_cyc), .IN3(n14333), .IN4(n18601), 
        .Q(n17710) );
  AO22X1 U36958 ( .IN1(n14332), .IN2(m3s11_cyc), .IN3(n14333), .IN4(n17822), 
        .Q(n17711) );
  AO22X1 U36959 ( .IN1(n14332), .IN2(m3s12_cyc), .IN3(n14333), .IN4(n17813), 
        .Q(n17712) );
  AO22X1 U36960 ( .IN1(n14332), .IN2(m3s13_cyc), .IN3(n14333), .IN4(n17814), 
        .Q(n17713) );
  AO22X1 U36961 ( .IN1(n14332), .IN2(test_so25), .IN3(n14333), .IN4(n17818), 
        .Q(n17714) );
  AO22X1 U36962 ( .IN1(n14332), .IN2(m3s15_cyc), .IN3(n14333), .IN4(n17783), 
        .Q(n17715) );
  AO22X1 U36963 ( .IN1(n14334), .IN2(m2s0_cyc), .IN3(n14335), .IN4(n18529), 
        .Q(n17716) );
  AO22X1 U36964 ( .IN1(n14334), .IN2(m2s1_cyc), .IN3(n14335), .IN4(n17862), 
        .Q(n17717) );
  AO22X1 U36965 ( .IN1(n14334), .IN2(test_so21), .IN3(n14335), .IN4(n17840), 
        .Q(n17718) );
  AO22X1 U36966 ( .IN1(n14334), .IN2(m2s3_cyc), .IN3(n14335), .IN4(n18535), 
        .Q(n17719) );
  AO22X1 U36967 ( .IN1(n14334), .IN2(m2s4_cyc), .IN3(n14335), .IN4(n17842), 
        .Q(n17720) );
  AO22X1 U36968 ( .IN1(n14334), .IN2(m2s5_cyc), .IN3(n14335), .IN4(n17841), 
        .Q(n17721) );
  AO22X1 U36969 ( .IN1(n14334), .IN2(m2s6_cyc), .IN3(n14335), .IN4(n18541), 
        .Q(n17722) );
  AO22X1 U36970 ( .IN1(n14334), .IN2(m2s7_cyc), .IN3(n14335), .IN4(n17861), 
        .Q(n17723) );
  AO22X1 U36971 ( .IN1(n14334), .IN2(m2s8_cyc), .IN3(n14335), .IN4(n17867), 
        .Q(n17724) );
  AO22X1 U36972 ( .IN1(n14334), .IN2(test_so22), .IN3(n14335), .IN4(n17879), 
        .Q(n17725) );
  AO22X1 U36973 ( .IN1(n14334), .IN2(m2s10_cyc), .IN3(n14335), .IN4(n18553), 
        .Q(n17726) );
  AO22X1 U36974 ( .IN1(n14334), .IN2(m2s11_cyc), .IN3(n14335), .IN4(n17852), 
        .Q(n17727) );
  AO22X1 U36975 ( .IN1(n14334), .IN2(m2s12_cyc), .IN3(n14335), .IN4(n18565), 
        .Q(n17728) );
  AO22X1 U36976 ( .IN1(n14334), .IN2(m2s13_cyc), .IN3(n14335), .IN4(n17848), 
        .Q(n17729) );
  AO22X1 U36977 ( .IN1(n14334), .IN2(m2s14_cyc), .IN3(n14335), .IN4(n17856), 
        .Q(n17730) );
  AO22X1 U36978 ( .IN1(n14334), .IN2(m2s15_cyc), .IN3(n14335), .IN4(n17786), 
        .Q(n17731) );
  AO22X1 U36979 ( .IN1(n14336), .IN2(m1s0_cyc), .IN3(n14337), .IN4(n18481), 
        .Q(n17732) );
  AO22X1 U36980 ( .IN1(n14336), .IN2(m1s1_cyc), .IN3(n14337), .IN4(n17826), 
        .Q(n17733) );
  AO22X1 U36981 ( .IN1(n14336), .IN2(m1s2_cyc), .IN3(n14337), .IN4(n17806), 
        .Q(n17734) );
  AO22X1 U36982 ( .IN1(n14336), .IN2(m1s3_cyc), .IN3(n14337), .IN4(n17805), 
        .Q(n17735) );
  AO22X1 U36983 ( .IN1(n14336), .IN2(test_so19), .IN3(n14337), .IN4(n17808), 
        .Q(n17736) );
  AO22X1 U36984 ( .IN1(n14336), .IN2(m1s5_cyc), .IN3(n14337), .IN4(n17807), 
        .Q(n17737) );
  AO22X1 U36985 ( .IN1(n14336), .IN2(m1s6_cyc), .IN3(n14337), .IN4(n17871), 
        .Q(n17738) );
  AO22X1 U36986 ( .IN1(n14336), .IN2(m1s7_cyc), .IN3(n14337), .IN4(n17884), 
        .Q(n17739) );
  AO22X1 U36987 ( .IN1(n14336), .IN2(m1s8_cyc), .IN3(n14337), .IN4(n17833), 
        .Q(n17740) );
  AO22X1 U36988 ( .IN1(n14336), .IN2(m1s9_cyc), .IN3(n14337), .IN4(n17876), 
        .Q(n17741) );
  AO22X1 U36989 ( .IN1(n14336), .IN2(m1s10_cyc), .IN3(n14337), .IN4(n18505), 
        .Q(n17742) );
  AO22X1 U36990 ( .IN1(n14336), .IN2(test_so20), .IN3(n14337), .IN4(n17823), 
        .Q(n17743) );
  AO22X1 U36991 ( .IN1(n14336), .IN2(m1s12_cyc), .IN3(n14337), .IN4(n17815), 
        .Q(n17744) );
  AO22X1 U36992 ( .IN1(n14336), .IN2(m1s13_cyc), .IN3(n14337), .IN4(n17816), 
        .Q(n17745) );
  AO22X1 U36993 ( .IN1(n14336), .IN2(m1s14_cyc), .IN3(n14337), .IN4(n17819), 
        .Q(n17746) );
  AO22X1 U36994 ( .IN1(n14336), .IN2(m1s15_cyc), .IN3(n14337), .IN4(n17784), 
        .Q(n17747) );
  AO22X1 U36995 ( .IN1(n14338), .IN2(m0s0_cyc), .IN3(n14339), .IN4(n18433), 
        .Q(n17748) );
  AO22X1 U36996 ( .IN1(n14338), .IN2(m0s1_cyc), .IN3(n14339), .IN4(n17864), 
        .Q(n17749) );
  AO22X1 U36997 ( .IN1(n14338), .IN2(m0s2_cyc), .IN3(n14339), .IN4(n17843), 
        .Q(n17750) );
  AO22X1 U36998 ( .IN1(n14338), .IN2(m0s3_cyc), .IN3(n14339), .IN4(n18439), 
        .Q(n17751) );
  AO22X1 U36999 ( .IN1(n14338), .IN2(m0s4_cyc), .IN3(n14339), .IN4(n17845), 
        .Q(n17752) );
  AO22X1 U37000 ( .IN1(n14338), .IN2(m0s5_cyc), .IN3(n14339), .IN4(n17844), 
        .Q(n17753) );
  AO22X1 U37001 ( .IN1(n14338), .IN2(test_so17), .IN3(n14339), .IN4(n18445), 
        .Q(n17754) );
  AO22X1 U37002 ( .IN1(n14338), .IN2(m0s7_cyc), .IN3(n14339), .IN4(n17863), 
        .Q(n17755) );
  AO22X1 U37003 ( .IN1(n14338), .IN2(m0s8_cyc), .IN3(n14339), .IN4(n17868), 
        .Q(n17756) );
  AO22X1 U37004 ( .IN1(n14338), .IN2(m0s9_cyc), .IN3(n14339), .IN4(n17880), 
        .Q(n17757) );
  AO22X1 U37005 ( .IN1(n14338), .IN2(m0s10_cyc), .IN3(n14339), .IN4(n18457), 
        .Q(n17758) );
  AO22X1 U37006 ( .IN1(n14338), .IN2(m0s11_cyc), .IN3(n14339), .IN4(n17853), 
        .Q(n17759) );
  AO22X1 U37007 ( .IN1(n14338), .IN2(m0s12_cyc), .IN3(n14339), .IN4(n18469), 
        .Q(n17760) );
  AO22X1 U37008 ( .IN1(n14338), .IN2(test_so18), .IN3(n14339), .IN4(n17849), 
        .Q(n17761) );
  AO22X1 U37009 ( .IN1(n14338), .IN2(m0s14_cyc), .IN3(n14339), .IN4(n17857), 
        .Q(n17762) );
  AO22X1 U37010 ( .IN1(n14338), .IN2(m0s15_cyc), .IN3(n14339), .IN4(n17787), 
        .Q(n17763) );
  NAND2X0 U37011 ( .IN1(conf15_4_), .IN2(n18086), .QN(n14279) );
  NAND2X0 U37012 ( .IN1(conf15_14_), .IN2(n18189), .QN(n14280) );
  NAND2X0 U37013 ( .IN1(conf15_6_), .IN2(n18087), .QN(n14276) );
  NAND2X0 U37014 ( .IN1(conf15_2_), .IN2(n18088), .QN(n14278) );
  NAND2X0 U37015 ( .IN1(conf15_12_), .IN2(n18190), .QN(n14283) );
  NAND2X0 U37016 ( .IN1(conf7_15_), .IN2(n18032), .QN(n13659) );
  NAND2X0 U37017 ( .IN1(conf7_7_), .IN2(n17965), .QN(n13643) );
  NAND2X0 U37018 ( .IN1(conf6_15_), .IN2(n18201), .QN(n13350) );
  NAND2X0 U37019 ( .IN1(conf6_7_), .IN2(n18102), .QN(n13334) );
  NAND2X0 U37020 ( .IN1(conf14_15_), .IN2(n18202), .QN(n11184) );
  NAND2X0 U37021 ( .IN1(conf14_7_), .IN2(n18103), .QN(n11168) );
  NAND2X0 U37022 ( .IN1(conf5_15_), .IN2(n18049), .QN(n13041) );
  NAND2X0 U37023 ( .IN1(conf5_7_), .IN2(n17993), .QN(n13025) );
  NAND2X0 U37024 ( .IN1(conf4_15_), .IN2(n18217), .QN(n12732) );
  NAND2X0 U37025 ( .IN1(conf4_7_), .IN2(n18130), .QN(n12716) );
  NAND2X0 U37026 ( .IN1(conf13_15_), .IN2(n18050), .QN(n10875) );
  NAND2X0 U37027 ( .IN1(conf13_7_), .IN2(n17994), .QN(n10859) );
  NAND2X0 U37028 ( .IN1(conf12_15_), .IN2(n18218), .QN(n10565) );
  NAND2X0 U37029 ( .IN1(conf12_7_), .IN2(n18131), .QN(n10549) );
  NAND2X0 U37030 ( .IN1(conf3_15_), .IN2(n18033), .QN(n12423) );
  NAND2X0 U37031 ( .IN1(conf3_7_), .IN2(n17966), .QN(n12407) );
  NAND2X0 U37032 ( .IN1(conf2_15_), .IN2(n18203), .QN(n12114) );
  NAND2X0 U37033 ( .IN1(conf2_7_), .IN2(n18104), .QN(n12098) );
  NAND2X0 U37034 ( .IN1(conf11_15_), .IN2(n18051), .QN(n10256) );
  NAND2X0 U37035 ( .IN1(conf11_7_), .IN2(n17995), .QN(n10240) );
  NAND2X0 U37036 ( .IN1(conf10_15_), .IN2(n18219), .QN(n9946) );
  NAND2X0 U37037 ( .IN1(conf10_7_), .IN2(n18132), .QN(n9930) );
  NAND2X0 U37038 ( .IN1(conf1_15_), .IN2(n18052), .QN(n11804) );
  NAND2X0 U37039 ( .IN1(conf1_7_), .IN2(n17996), .QN(n11788) );
  NAND2X0 U37040 ( .IN1(conf0_15_), .IN2(n18220), .QN(n11494) );
  NAND2X0 U37041 ( .IN1(conf0_7_), .IN2(n18133), .QN(n11478) );
  NAND2X0 U37042 ( .IN1(conf9_15_), .IN2(n18034), .QN(n9636) );
  NAND2X0 U37043 ( .IN1(conf9_7_), .IN2(n17967), .QN(n9620) );
  NAND2X0 U37044 ( .IN1(conf8_15_), .IN2(n18204), .QN(n9325) );
  NAND2X0 U37045 ( .IN1(conf8_7_), .IN2(n18105), .QN(n9309) );
  NAND2X0 U37046 ( .IN1(conf7_3_), .IN2(n17968), .QN(n13649) );
  NAND2X0 U37047 ( .IN1(conf7_5_), .IN2(n17969), .QN(n13646) );
  NAND2X0 U37048 ( .IN1(conf6_3_), .IN2(n18106), .QN(n13340) );
  NAND2X0 U37049 ( .IN1(conf6_5_), .IN2(n18107), .QN(n13337) );
  NAND2X0 U37050 ( .IN1(conf14_3_), .IN2(n18108), .QN(n11174) );
  NAND2X0 U37051 ( .IN1(conf14_5_), .IN2(n18109), .QN(n11171) );
  NAND2X0 U37052 ( .IN1(conf5_3_), .IN2(n17997), .QN(n13031) );
  NAND2X0 U37053 ( .IN1(conf5_5_), .IN2(n17998), .QN(n13028) );
  NAND2X0 U37054 ( .IN1(conf4_3_), .IN2(n18134), .QN(n12722) );
  NAND2X0 U37055 ( .IN1(conf4_5_), .IN2(n18135), .QN(n12719) );
  NAND2X0 U37056 ( .IN1(conf13_3_), .IN2(n17999), .QN(n10865) );
  NAND2X0 U37057 ( .IN1(conf13_5_), .IN2(n18000), .QN(n10862) );
  NAND2X0 U37058 ( .IN1(conf12_3_), .IN2(n18136), .QN(n10555) );
  NAND2X0 U37059 ( .IN1(conf12_5_), .IN2(n18137), .QN(n10552) );
  NAND2X0 U37060 ( .IN1(conf3_3_), .IN2(n17970), .QN(n12413) );
  NAND2X0 U37061 ( .IN1(conf3_5_), .IN2(n17971), .QN(n12410) );
  NAND2X0 U37062 ( .IN1(conf2_3_), .IN2(n18110), .QN(n12104) );
  NAND2X0 U37063 ( .IN1(conf2_5_), .IN2(n18111), .QN(n12101) );
  NAND2X0 U37064 ( .IN1(conf11_3_), .IN2(n18001), .QN(n10246) );
  NAND2X0 U37065 ( .IN1(conf11_5_), .IN2(n18002), .QN(n10243) );
  NAND2X0 U37066 ( .IN1(conf10_3_), .IN2(n18138), .QN(n9936) );
  NAND2X0 U37067 ( .IN1(conf10_5_), .IN2(n18139), .QN(n9933) );
  NAND2X0 U37068 ( .IN1(conf1_3_), .IN2(n18003), .QN(n11794) );
  NAND2X0 U37069 ( .IN1(conf1_5_), .IN2(n18004), .QN(n11791) );
  NAND2X0 U37070 ( .IN1(conf0_3_), .IN2(n18140), .QN(n11484) );
  NAND2X0 U37071 ( .IN1(conf0_5_), .IN2(n18141), .QN(n11481) );
  NAND2X0 U37072 ( .IN1(conf9_3_), .IN2(n17972), .QN(n9626) );
  NAND2X0 U37073 ( .IN1(conf9_5_), .IN2(n17973), .QN(n9623) );
  NAND2X0 U37074 ( .IN1(conf8_3_), .IN2(n18112), .QN(n9315) );
  NAND2X0 U37075 ( .IN1(conf8_5_), .IN2(n18113), .QN(n9312) );
  NAND2X0 U37076 ( .IN1(conf7_1_), .IN2(n18021), .QN(n13652) );
  NAND2X0 U37077 ( .IN1(conf6_1_), .IN2(n18142), .QN(n13343) );
  NAND2X0 U37078 ( .IN1(conf14_1_), .IN2(n18143), .QN(n11177) );
  NAND2X0 U37079 ( .IN1(conf5_1_), .IN2(n18025), .QN(n13034) );
  NAND2X0 U37080 ( .IN1(conf4_1_), .IN2(n18146), .QN(n12725) );
  NAND2X0 U37081 ( .IN1(conf13_1_), .IN2(n18026), .QN(n10868) );
  NAND2X0 U37082 ( .IN1(conf12_1_), .IN2(n18147), .QN(n10558) );
  NAND2X0 U37083 ( .IN1(conf3_1_), .IN2(n18022), .QN(n12416) );
  NAND2X0 U37084 ( .IN1(conf2_1_), .IN2(n18144), .QN(n12107) );
  NAND2X0 U37085 ( .IN1(conf11_1_), .IN2(n18027), .QN(n10249) );
  NAND2X0 U37086 ( .IN1(conf10_1_), .IN2(n18148), .QN(n9939) );
  NAND2X0 U37087 ( .IN1(conf1_1_), .IN2(n18028), .QN(n11797) );
  NAND2X0 U37088 ( .IN1(conf0_1_), .IN2(n18149), .QN(n11487) );
  NAND2X0 U37089 ( .IN1(conf9_1_), .IN2(n18023), .QN(n9629) );
  NAND2X0 U37090 ( .IN1(conf8_1_), .IN2(n18145), .QN(n9318) );
  NAND3X0 U37091 ( .IN1(n3884), .IN2(n3885), .IN3(n3883), .QN(n13902) );
  NAND3X0 U37092 ( .IN1(n3839), .IN2(n3840), .IN3(n3838), .QN(n13593) );
  NAND3X0 U37093 ( .IN1(n4199), .IN2(n4200), .IN3(n4198), .QN(n11427) );
  NAND3X0 U37094 ( .IN1(n3794), .IN2(n3795), .IN3(n3793), .QN(n13284) );
  NAND3X0 U37095 ( .IN1(n3749), .IN2(n3750), .IN3(n3748), .QN(n12975) );
  NAND3X0 U37096 ( .IN1(n4154), .IN2(n4155), .IN3(n4153), .QN(n11118) );
  NAND3X0 U37097 ( .IN1(n4109), .IN2(n4110), .IN3(n4108), .QN(n10808) );
  NAND3X0 U37098 ( .IN1(n3704), .IN2(n3705), .IN3(n3703), .QN(n12666) );
  NAND3X0 U37099 ( .IN1(n3659), .IN2(n3660), .IN3(n3658), .QN(n12357) );
  NAND3X0 U37100 ( .IN1(n4064), .IN2(n4065), .IN3(n4063), .QN(n10499) );
  NAND3X0 U37101 ( .IN1(n4019), .IN2(n4020), .IN3(n4018), .QN(n10189) );
  NAND3X0 U37102 ( .IN1(n3614), .IN2(n3615), .IN3(n3613), .QN(n12047) );
  NAND3X0 U37103 ( .IN1(n3569), .IN2(n3570), .IN3(n3568), .QN(n11737) );
  NAND3X0 U37104 ( .IN1(n3974), .IN2(n3975), .IN3(n3973), .QN(n9879) );
  NAND3X0 U37105 ( .IN1(n3929), .IN2(n3930), .IN3(n3928), .QN(n9568) );
  NAND3X0 U37106 ( .IN1(n4228), .IN2(n4229), .IN3(n4227), .QN(n13969) );
  NAND3X0 U37107 ( .IN1(n4244), .IN2(n4245), .IN3(n4243), .QN(n14176) );
  NAND3X0 U37108 ( .IN1(n4236), .IN2(n4237), .IN3(n4235), .QN(n14109) );
  NAND2X0 U37109 ( .IN1(conf7_4_), .IN2(n18089), .QN(n13645) );
  NAND2X0 U37110 ( .IN1(conf7_14_), .IN2(n18191), .QN(n13658) );
  NAND2X0 U37111 ( .IN1(conf7_6_), .IN2(n18090), .QN(n13642) );
  NAND2X0 U37112 ( .IN1(conf6_4_), .IN2(n17977), .QN(n13336) );
  NAND2X0 U37113 ( .IN1(conf6_14_), .IN2(n18037), .QN(n13349) );
  NAND2X0 U37114 ( .IN1(conf6_6_), .IN2(n17978), .QN(n13333) );
  NAND2X0 U37115 ( .IN1(conf14_4_), .IN2(n17979), .QN(n11170) );
  NAND2X0 U37116 ( .IN1(conf14_14_), .IN2(n18038), .QN(n11183) );
  NAND2X0 U37117 ( .IN1(conf14_6_), .IN2(n17980), .QN(n11167) );
  NAND2X0 U37118 ( .IN1(conf5_4_), .IN2(n18114), .QN(n13027) );
  NAND2X0 U37119 ( .IN1(conf5_14_), .IN2(n18205), .QN(n13040) );
  NAND2X0 U37120 ( .IN1(conf5_6_), .IN2(n18115), .QN(n13024) );
  NAND2X0 U37121 ( .IN1(conf4_4_), .IN2(n18005), .QN(n12718) );
  NAND2X0 U37122 ( .IN1(conf4_14_), .IN2(n18053), .QN(n12731) );
  NAND2X0 U37123 ( .IN1(conf4_6_), .IN2(n18006), .QN(n12715) );
  NAND2X0 U37124 ( .IN1(conf13_4_), .IN2(n18116), .QN(n10861) );
  NAND2X0 U37125 ( .IN1(conf13_14_), .IN2(n18206), .QN(n10874) );
  NAND2X0 U37126 ( .IN1(conf13_6_), .IN2(n18117), .QN(n10858) );
  NAND2X0 U37127 ( .IN1(conf12_4_), .IN2(n18007), .QN(n10551) );
  NAND2X0 U37128 ( .IN1(conf12_14_), .IN2(n18054), .QN(n10564) );
  NAND2X0 U37129 ( .IN1(conf12_6_), .IN2(n18008), .QN(n10548) );
  NAND2X0 U37130 ( .IN1(conf3_4_), .IN2(n18091), .QN(n12409) );
  NAND2X0 U37131 ( .IN1(conf3_14_), .IN2(n18192), .QN(n12422) );
  NAND2X0 U37132 ( .IN1(conf3_6_), .IN2(n18092), .QN(n12406) );
  NAND2X0 U37133 ( .IN1(conf2_4_), .IN2(n17981), .QN(n12100) );
  NAND2X0 U37134 ( .IN1(conf2_14_), .IN2(n18039), .QN(n12113) );
  NAND2X0 U37135 ( .IN1(conf2_6_), .IN2(n17982), .QN(n12097) );
  NAND2X0 U37136 ( .IN1(conf11_4_), .IN2(n18118), .QN(n10242) );
  NAND2X0 U37137 ( .IN1(conf11_14_), .IN2(n18207), .QN(n10255) );
  NAND2X0 U37138 ( .IN1(conf11_6_), .IN2(n18119), .QN(n10239) );
  NAND2X0 U37139 ( .IN1(conf10_4_), .IN2(n18009), .QN(n9932) );
  NAND2X0 U37140 ( .IN1(conf10_14_), .IN2(n18055), .QN(n9945) );
  NAND2X0 U37141 ( .IN1(conf10_6_), .IN2(n18010), .QN(n9929) );
  NAND2X0 U37142 ( .IN1(conf1_4_), .IN2(n18120), .QN(n11790) );
  NAND2X0 U37143 ( .IN1(conf1_14_), .IN2(n18208), .QN(n11803) );
  NAND2X0 U37144 ( .IN1(conf1_6_), .IN2(n18121), .QN(n11787) );
  NAND2X0 U37145 ( .IN1(conf0_4_), .IN2(n18011), .QN(n11480) );
  NAND2X0 U37146 ( .IN1(conf0_14_), .IN2(n18056), .QN(n11493) );
  NAND2X0 U37147 ( .IN1(conf0_6_), .IN2(n18012), .QN(n11477) );
  NAND2X0 U37148 ( .IN1(conf9_4_), .IN2(n18093), .QN(n9622) );
  NAND2X0 U37149 ( .IN1(conf9_14_), .IN2(n18193), .QN(n9635) );
  NAND2X0 U37150 ( .IN1(conf9_6_), .IN2(n18094), .QN(n9619) );
  NAND2X0 U37151 ( .IN1(conf8_4_), .IN2(n17983), .QN(n9311) );
  NAND2X0 U37152 ( .IN1(conf8_14_), .IN2(n18040), .QN(n9324) );
  NAND2X0 U37153 ( .IN1(conf8_6_), .IN2(n17984), .QN(n9308) );
  NAND2X0 U37154 ( .IN1(conf7_2_), .IN2(n18095), .QN(n13648) );
  NAND2X0 U37155 ( .IN1(conf6_2_), .IN2(n17985), .QN(n13339) );
  NAND2X0 U37156 ( .IN1(conf14_2_), .IN2(n17986), .QN(n11173) );
  NAND2X0 U37157 ( .IN1(conf5_2_), .IN2(n18122), .QN(n13030) );
  NAND2X0 U37158 ( .IN1(conf4_2_), .IN2(n18013), .QN(n12721) );
  NAND2X0 U37159 ( .IN1(conf13_2_), .IN2(n18123), .QN(n10864) );
  NAND2X0 U37160 ( .IN1(conf12_2_), .IN2(n18014), .QN(n10554) );
  NAND2X0 U37161 ( .IN1(conf3_2_), .IN2(n18096), .QN(n12412) );
  NAND2X0 U37162 ( .IN1(conf2_2_), .IN2(n17987), .QN(n12103) );
  NAND2X0 U37163 ( .IN1(conf11_2_), .IN2(n18124), .QN(n10245) );
  NAND2X0 U37164 ( .IN1(conf10_2_), .IN2(n18015), .QN(n9935) );
  NAND2X0 U37165 ( .IN1(conf1_2_), .IN2(n18125), .QN(n11793) );
  NAND2X0 U37166 ( .IN1(conf0_2_), .IN2(n18016), .QN(n11483) );
  NAND2X0 U37167 ( .IN1(conf9_2_), .IN2(n18097), .QN(n9625) );
  NAND2X0 U37168 ( .IN1(conf8_2_), .IN2(n17988), .QN(n9314) );
  NAND2X0 U37169 ( .IN1(conf7_12_), .IN2(n18194), .QN(n13661) );
  NAND2X0 U37170 ( .IN1(conf6_12_), .IN2(n18041), .QN(n13352) );
  NAND2X0 U37171 ( .IN1(conf14_12_), .IN2(n18042), .QN(n11186) );
  NAND2X0 U37172 ( .IN1(conf5_12_), .IN2(n18209), .QN(n13043) );
  NAND2X0 U37173 ( .IN1(conf4_12_), .IN2(n18057), .QN(n12734) );
  NAND2X0 U37174 ( .IN1(conf13_12_), .IN2(n18210), .QN(n10877) );
  NAND2X0 U37175 ( .IN1(conf12_12_), .IN2(n18058), .QN(n10567) );
  NAND2X0 U37176 ( .IN1(conf3_12_), .IN2(n18195), .QN(n12425) );
  NAND2X0 U37177 ( .IN1(conf2_12_), .IN2(n18043), .QN(n12116) );
  NAND2X0 U37178 ( .IN1(conf11_12_), .IN2(n18211), .QN(n10258) );
  NAND2X0 U37179 ( .IN1(conf10_12_), .IN2(n18059), .QN(n9948) );
  NAND2X0 U37180 ( .IN1(conf1_12_), .IN2(n18212), .QN(n11806) );
  NAND2X0 U37181 ( .IN1(conf0_12_), .IN2(n18060), .QN(n11496) );
  NAND2X0 U37182 ( .IN1(conf9_12_), .IN2(n18196), .QN(n9638) );
  NAND2X0 U37183 ( .IN1(conf8_12_), .IN2(n18044), .QN(n9327) );
  NAND3X0 U37184 ( .IN1(n3868), .IN2(n3869), .IN3(n3867), .QN(n13836) );
  NAND3X0 U37185 ( .IN1(n3876), .IN2(n3877), .IN3(n3875), .QN(n13708) );
  NAND3X0 U37186 ( .IN1(n3823), .IN2(n3824), .IN3(n3822), .QN(n13527) );
  NAND3X0 U37187 ( .IN1(n3831), .IN2(n3832), .IN3(n3830), .QN(n13399) );
  NAND3X0 U37188 ( .IN1(n4183), .IN2(n4184), .IN3(n4182), .QN(n11361) );
  NAND3X0 U37189 ( .IN1(n4191), .IN2(n4192), .IN3(n4190), .QN(n11233) );
  NAND3X0 U37190 ( .IN1(n3778), .IN2(n3779), .IN3(n3777), .QN(n13218) );
  NAND3X0 U37191 ( .IN1(n3786), .IN2(n3787), .IN3(n3785), .QN(n13090) );
  NAND3X0 U37192 ( .IN1(n3733), .IN2(n3734), .IN3(n3732), .QN(n12909) );
  NAND3X0 U37193 ( .IN1(n3741), .IN2(n3742), .IN3(n3740), .QN(n12781) );
  NAND3X0 U37194 ( .IN1(n4138), .IN2(n4139), .IN3(n4137), .QN(n11052) );
  NAND3X0 U37195 ( .IN1(n4146), .IN2(n4147), .IN3(n4145), .QN(n10924) );
  NAND3X0 U37196 ( .IN1(n4093), .IN2(n4094), .IN3(n4092), .QN(n10742) );
  NAND3X0 U37197 ( .IN1(n4101), .IN2(n4102), .IN3(n4100), .QN(n10614) );
  NAND3X0 U37198 ( .IN1(n3688), .IN2(n3689), .IN3(n3687), .QN(n12600) );
  NAND3X0 U37199 ( .IN1(n3696), .IN2(n3697), .IN3(n3695), .QN(n12472) );
  NAND3X0 U37200 ( .IN1(n3643), .IN2(n3644), .IN3(n3642), .QN(n12291) );
  NAND3X0 U37201 ( .IN1(n3651), .IN2(n3652), .IN3(n3650), .QN(n12163) );
  NAND3X0 U37202 ( .IN1(n4048), .IN2(n4049), .IN3(n4047), .QN(n10433) );
  NAND3X0 U37203 ( .IN1(n4056), .IN2(n4057), .IN3(n4055), .QN(n10305) );
  NAND3X0 U37204 ( .IN1(n4003), .IN2(n4004), .IN3(n4002), .QN(n10123) );
  NAND3X0 U37205 ( .IN1(n4011), .IN2(n4012), .IN3(n4010), .QN(n9995) );
  NAND3X0 U37206 ( .IN1(n3598), .IN2(n3599), .IN3(n3597), .QN(n11981) );
  NAND3X0 U37207 ( .IN1(n3606), .IN2(n3607), .IN3(n3605), .QN(n11853) );
  NAND3X0 U37208 ( .IN1(n3553), .IN2(n3554), .IN3(n3552), .QN(n11671) );
  NAND3X0 U37209 ( .IN1(n3561), .IN2(n3562), .IN3(n3560), .QN(n11543) );
  NAND3X0 U37210 ( .IN1(n3958), .IN2(n3959), .IN3(n3957), .QN(n9813) );
  NAND3X0 U37211 ( .IN1(n3966), .IN2(n3967), .IN3(n3965), .QN(n9685) );
  NAND3X0 U37212 ( .IN1(n3913), .IN2(n3914), .IN3(n3912), .QN(n9502) );
  NAND3X0 U37213 ( .IN1(n3921), .IN2(n3922), .IN3(n3920), .QN(n9374) );
  NAND3X0 U37214 ( .IN1(n3884), .IN2(n3885), .IN3(s7_msel_gnt_p3[0]), .QN(
        n13903) );
  NAND3X0 U37215 ( .IN1(n3868), .IN2(n3869), .IN3(s7_msel_gnt_p1[0]), .QN(
        n13837) );
  NAND3X0 U37216 ( .IN1(n3876), .IN2(n3877), .IN3(test_so68), .QN(n13709) );
  NAND3X0 U37217 ( .IN1(n3839), .IN2(n3840), .IN3(s6_msel_gnt_p3_0_), .QN(
        n13594) );
  NAND3X0 U37218 ( .IN1(n3823), .IN2(n3824), .IN3(s6_msel_gnt_p1_0_), .QN(
        n13528) );
  NAND3X0 U37219 ( .IN1(n3831), .IN2(n3832), .IN3(s6_msel_gnt_p2[0]), .QN(
        n13400) );
  NAND3X0 U37220 ( .IN1(n4199), .IN2(n4200), .IN3(s14_msel_gnt_p3[0]), .QN(
        n11428) );
  NAND3X0 U37221 ( .IN1(n4183), .IN2(n4184), .IN3(s14_msel_gnt_p1[0]), .QN(
        n11362) );
  NAND3X0 U37222 ( .IN1(n4191), .IN2(n4192), .IN3(s14_msel_gnt_p2_0_), .QN(
        n11234) );
  NAND3X0 U37223 ( .IN1(n3794), .IN2(n3795), .IN3(s5_msel_gnt_p3_0_), .QN(
        n13285) );
  NAND3X0 U37224 ( .IN1(n3778), .IN2(n3779), .IN3(s5_msel_gnt_p1_0_), .QN(
        n13219) );
  NAND3X0 U37225 ( .IN1(n3786), .IN2(n3787), .IN3(s5_msel_gnt_p2[0]), .QN(
        n13091) );
  NAND3X0 U37226 ( .IN1(n3749), .IN2(n3750), .IN3(test_so57), .QN(n12976) );
  NAND3X0 U37227 ( .IN1(n3733), .IN2(n3734), .IN3(test_so56), .QN(n12910) );
  NAND3X0 U37228 ( .IN1(n3741), .IN2(n3742), .IN3(s4_msel_gnt_p2[0]), .QN(
        n12782) );
  NAND3X0 U37229 ( .IN1(n4154), .IN2(n4155), .IN3(s13_msel_gnt_p3[0]), .QN(
        n11119) );
  NAND3X0 U37230 ( .IN1(n4138), .IN2(n4139), .IN3(s13_msel_gnt_p1[0]), .QN(
        n11053) );
  NAND3X0 U37231 ( .IN1(n4146), .IN2(n4147), .IN3(test_so91), .QN(n10925) );
  NAND3X0 U37232 ( .IN1(n4109), .IN2(n4110), .IN3(s12_msel_gnt_p3_0_), .QN(
        n10809) );
  NAND3X0 U37233 ( .IN1(n4093), .IN2(n4094), .IN3(s12_msel_gnt_p1_0_), .QN(
        n10743) );
  NAND3X0 U37234 ( .IN1(n4101), .IN2(n4102), .IN3(s12_msel_gnt_p2[0]), .QN(
        n10615) );
  NAND3X0 U37235 ( .IN1(n3704), .IN2(n3705), .IN3(s3_msel_gnt_p3[0]), .QN(
        n12667) );
  NAND3X0 U37236 ( .IN1(n3688), .IN2(n3689), .IN3(s3_msel_gnt_p1[0]), .QN(
        n12601) );
  NAND3X0 U37237 ( .IN1(n3696), .IN2(n3697), .IN3(s3_msel_gnt_p2_0_), .QN(
        n12473) );
  NAND3X0 U37238 ( .IN1(n3659), .IN2(n3660), .IN3(s2_msel_gnt_p3[0]), .QN(
        n12358) );
  NAND3X0 U37239 ( .IN1(n3643), .IN2(n3644), .IN3(s2_msel_gnt_p1[0]), .QN(
        n12292) );
  NAND3X0 U37240 ( .IN1(n3651), .IN2(n3652), .IN3(s2_msel_gnt_p2_0_), .QN(
        n12164) );
  NAND3X0 U37241 ( .IN1(n4064), .IN2(n4065), .IN3(s11_msel_gnt_p3_0_), .QN(
        n10500) );
  NAND3X0 U37242 ( .IN1(n4048), .IN2(n4049), .IN3(s11_msel_gnt_p1_0_), .QN(
        n10434) );
  NAND3X0 U37243 ( .IN1(n4056), .IN2(n4057), .IN3(s11_msel_gnt_p2[0]), .QN(
        n10306) );
  NAND3X0 U37244 ( .IN1(n4019), .IN2(n4020), .IN3(test_so80), .QN(n10190) );
  NAND3X0 U37245 ( .IN1(n4003), .IN2(n4004), .IN3(test_so79), .QN(n10124) );
  NAND3X0 U37246 ( .IN1(n4011), .IN2(n4012), .IN3(s10_msel_gnt_p2[0]), .QN(
        n9996) );
  NAND3X0 U37247 ( .IN1(n3614), .IN2(n3615), .IN3(s1_msel_gnt_p3[0]), .QN(
        n12048) );
  NAND3X0 U37248 ( .IN1(n3598), .IN2(n3599), .IN3(s1_msel_gnt_p1[0]), .QN(
        n11982) );
  NAND3X0 U37249 ( .IN1(n3606), .IN2(n3607), .IN3(test_so45), .QN(n11854) );
  NAND3X0 U37250 ( .IN1(n3569), .IN2(n3570), .IN3(s0_msel_gnt_p3_0_), .QN(
        n11738) );
  NAND3X0 U37251 ( .IN1(n3553), .IN2(n3554), .IN3(s0_msel_gnt_p1_0_), .QN(
        n11672) );
  NAND3X0 U37252 ( .IN1(n3561), .IN2(n3562), .IN3(s0_msel_gnt_p2[0]), .QN(
        n11544) );
  NAND3X0 U37253 ( .IN1(n3974), .IN2(n3975), .IN3(s9_msel_gnt_p3[0]), .QN(
        n9880) );
  NAND3X0 U37254 ( .IN1(n3958), .IN2(n3959), .IN3(s9_msel_gnt_p1[0]), .QN(
        n9814) );
  NAND3X0 U37255 ( .IN1(n3966), .IN2(n3967), .IN3(s9_msel_gnt_p2_0_), .QN(
        n9686) );
  NAND3X0 U37256 ( .IN1(n3929), .IN2(n3930), .IN3(s8_msel_gnt_p3[0]), .QN(
        n9569) );
  NAND3X0 U37257 ( .IN1(n3913), .IN2(n3914), .IN3(s8_msel_gnt_p1[0]), .QN(
        n9503) );
  NAND3X0 U37258 ( .IN1(n3921), .IN2(n3922), .IN3(s8_msel_gnt_p2_0_), .QN(
        n9375) );
  NAND3X0 U37259 ( .IN1(n4228), .IN2(n4229), .IN3(s15_msel_gnt_p1[0]), .QN(
        n13970) );
  NAND3X0 U37260 ( .IN1(n4244), .IN2(n4245), .IN3(s15_msel_gnt_p3[0]), .QN(
        n14177) );
  NAND3X0 U37261 ( .IN1(n4236), .IN2(n4237), .IN3(s15_msel_gnt_p2_0_), .QN(
        n14110) );
  NAND2X0 U37262 ( .IN1(conf15_5_), .IN2(n17974), .QN(n14291) );
  NAND2X0 U37263 ( .IN1(conf15_3_), .IN2(n17975), .QN(n14292) );
  NAND2X0 U37264 ( .IN1(conf15_13_), .IN2(n18035), .QN(n14299) );
  NAND2X0 U37265 ( .IN1(conf15_15_), .IN2(n18036), .QN(n14298) );
  NAND2X0 U37266 ( .IN1(conf15_7_), .IN2(n17976), .QN(n14290) );
  NAND2X0 U37267 ( .IN1(conf15_1_), .IN2(n18024), .QN(n14293) );
  NAND2X0 U37268 ( .IN1(test_so16), .IN2(n18098), .QN(n14281) );
  NAND2X0 U37269 ( .IN1(test_so8), .IN2(n18099), .QN(n13651) );
  NAND2X0 U37270 ( .IN1(test_so7), .IN2(n17989), .QN(n13342) );
  NAND2X0 U37271 ( .IN1(test_so15), .IN2(n17990), .QN(n11176) );
  NAND2X0 U37272 ( .IN1(test_so6), .IN2(n18126), .QN(n13033) );
  NAND2X0 U37273 ( .IN1(test_so5), .IN2(n18017), .QN(n12724) );
  NAND2X0 U37274 ( .IN1(test_so14), .IN2(n18127), .QN(n10867) );
  NAND2X0 U37275 ( .IN1(test_so13), .IN2(n18018), .QN(n10557) );
  NAND2X0 U37276 ( .IN1(test_so4), .IN2(n18100), .QN(n12415) );
  NAND2X0 U37277 ( .IN1(test_so3), .IN2(n17991), .QN(n12106) );
  NAND2X0 U37278 ( .IN1(test_so12), .IN2(n18128), .QN(n10248) );
  NAND2X0 U37279 ( .IN1(test_so11), .IN2(n18019), .QN(n9938) );
  NAND2X0 U37280 ( .IN1(test_so2), .IN2(n18129), .QN(n11796) );
  NAND2X0 U37281 ( .IN1(test_so1), .IN2(n18020), .QN(n11486) );
  NAND2X0 U37282 ( .IN1(test_so10), .IN2(n18101), .QN(n9628) );
  NAND2X0 U37283 ( .IN1(test_so9), .IN2(n17992), .QN(n9317) );
  NAND3X0 U37284 ( .IN1(s7_msel_gnt_p3[1]), .IN2(s7_msel_gnt_p3[2]), .IN3(
        s7_msel_gnt_p3[0]), .QN(n13927) );
  NAND3X0 U37285 ( .IN1(s6_msel_gnt_p3_1_), .IN2(test_so65), .IN3(
        s6_msel_gnt_p3_0_), .QN(n13618) );
  NAND3X0 U37286 ( .IN1(s14_msel_gnt_p3[1]), .IN2(s14_msel_gnt_p3[2]), .IN3(
        s14_msel_gnt_p3[0]), .QN(n11452) );
  NAND3X0 U37287 ( .IN1(test_so61), .IN2(s5_msel_gnt_p3_2_), .IN3(
        s5_msel_gnt_p3_0_), .QN(n13309) );
  NAND3X0 U37288 ( .IN1(s4_msel_gnt_p3_1_), .IN2(s4_msel_gnt_p3_2_), .IN3(
        test_so57), .QN(n13000) );
  NAND3X0 U37289 ( .IN1(s13_msel_gnt_p3[1]), .IN2(s13_msel_gnt_p3[2]), .IN3(
        s13_msel_gnt_p3[0]), .QN(n11143) );
  NAND3X0 U37290 ( .IN1(s12_msel_gnt_p3_1_), .IN2(test_so88), .IN3(
        s12_msel_gnt_p3_0_), .QN(n10833) );
  NAND3X0 U37291 ( .IN1(s3_msel_gnt_p3[1]), .IN2(s3_msel_gnt_p3[2]), .IN3(
        s3_msel_gnt_p3[0]), .QN(n12691) );
  NAND3X0 U37292 ( .IN1(s2_msel_gnt_p3[1]), .IN2(s2_msel_gnt_p3[2]), .IN3(
        s2_msel_gnt_p3[0]), .QN(n12382) );
  NAND3X0 U37293 ( .IN1(test_so84), .IN2(s11_msel_gnt_p3_2_), .IN3(
        s11_msel_gnt_p3_0_), .QN(n10524) );
  NAND3X0 U37294 ( .IN1(s10_msel_gnt_p3_1_), .IN2(s10_msel_gnt_p3_2_), .IN3(
        test_so80), .QN(n10214) );
  NAND3X0 U37295 ( .IN1(s1_msel_gnt_p3[1]), .IN2(s1_msel_gnt_p3[2]), .IN3(
        s1_msel_gnt_p3[0]), .QN(n12072) );
  NAND3X0 U37296 ( .IN1(s0_msel_gnt_p3_1_), .IN2(test_so42), .IN3(
        s0_msel_gnt_p3_0_), .QN(n11762) );
  NAND3X0 U37297 ( .IN1(s9_msel_gnt_p3[1]), .IN2(s9_msel_gnt_p3[2]), .IN3(
        s9_msel_gnt_p3[0]), .QN(n9904) );
  NAND3X0 U37298 ( .IN1(s8_msel_gnt_p3[1]), .IN2(s8_msel_gnt_p3[2]), .IN3(
        s8_msel_gnt_p3[0]), .QN(n9593) );
  NAND3X0 U37299 ( .IN1(s15_msel_gnt_p3[1]), .IN2(s15_msel_gnt_p3[2]), .IN3(
        s15_msel_gnt_p3[0]), .QN(n14201) );
  NAND3X0 U37300 ( .IN1(s7_msel_gnt_p2_1_), .IN2(s7_msel_gnt_p2_2_), .IN3(
        test_so68), .QN(n13731) );
  NAND3X0 U37301 ( .IN1(s6_msel_gnt_p2[1]), .IN2(s6_msel_gnt_p2[2]), .IN3(
        s6_msel_gnt_p2[0]), .QN(n13422) );
  NAND3X0 U37302 ( .IN1(test_so95), .IN2(s14_msel_gnt_p2_2_), .IN3(
        s14_msel_gnt_p2_0_), .QN(n11256) );
  NAND3X0 U37303 ( .IN1(s5_msel_gnt_p2[1]), .IN2(s5_msel_gnt_p2[2]), .IN3(
        s5_msel_gnt_p2[0]), .QN(n13113) );
  NAND3X0 U37304 ( .IN1(s4_msel_gnt_p2[1]), .IN2(s4_msel_gnt_p2[2]), .IN3(
        s4_msel_gnt_p2[0]), .QN(n12804) );
  NAND3X0 U37305 ( .IN1(s13_msel_gnt_p2_1_), .IN2(s13_msel_gnt_p2_2_), .IN3(
        test_so91), .QN(n10947) );
  NAND3X0 U37306 ( .IN1(s12_msel_gnt_p2[1]), .IN2(s12_msel_gnt_p2[2]), .IN3(
        s12_msel_gnt_p2[0]), .QN(n10637) );
  NAND3X0 U37307 ( .IN1(s3_msel_gnt_p2_1_), .IN2(test_so53), .IN3(
        s3_msel_gnt_p2_0_), .QN(n12495) );
  NAND3X0 U37308 ( .IN1(test_so49), .IN2(s2_msel_gnt_p2_2_), .IN3(
        s2_msel_gnt_p2_0_), .QN(n12186) );
  NAND3X0 U37309 ( .IN1(s11_msel_gnt_p2[1]), .IN2(s11_msel_gnt_p2[2]), .IN3(
        s11_msel_gnt_p2[0]), .QN(n10328) );
  NAND3X0 U37310 ( .IN1(s10_msel_gnt_p2[1]), .IN2(s10_msel_gnt_p2[2]), .IN3(
        s10_msel_gnt_p2[0]), .QN(n10018) );
  NAND3X0 U37311 ( .IN1(s1_msel_gnt_p2_1_), .IN2(s1_msel_gnt_p2_2_), .IN3(
        test_so45), .QN(n11876) );
  NAND3X0 U37312 ( .IN1(s0_msel_gnt_p2[1]), .IN2(s0_msel_gnt_p2[2]), .IN3(
        s0_msel_gnt_p2[0]), .QN(n11566) );
  NAND3X0 U37313 ( .IN1(s9_msel_gnt_p2_1_), .IN2(test_so76), .IN3(
        s9_msel_gnt_p2_0_), .QN(n9708) );
  NAND3X0 U37314 ( .IN1(test_so72), .IN2(s8_msel_gnt_p2_2_), .IN3(
        s8_msel_gnt_p2_0_), .QN(n9397) );
  NAND3X0 U37315 ( .IN1(s15_msel_gnt_p2_1_), .IN2(test_so99), .IN3(
        s15_msel_gnt_p2_0_), .QN(n14135) );
  NAND3X0 U37316 ( .IN1(s7_msel_gnt_p1[1]), .IN2(s7_msel_gnt_p1[2]), .IN3(
        s7_msel_gnt_p1[0]), .QN(n13862) );
  NAND3X0 U37317 ( .IN1(s6_msel_gnt_p1_1_), .IN2(test_so64), .IN3(
        s6_msel_gnt_p1_0_), .QN(n13553) );
  NAND3X0 U37318 ( .IN1(s14_msel_gnt_p1[1]), .IN2(s14_msel_gnt_p1[2]), .IN3(
        s14_msel_gnt_p1[0]), .QN(n11387) );
  NAND3X0 U37319 ( .IN1(test_so60), .IN2(s5_msel_gnt_p1_2_), .IN3(
        s5_msel_gnt_p1_0_), .QN(n13244) );
  NAND3X0 U37320 ( .IN1(s4_msel_gnt_p1_1_), .IN2(s4_msel_gnt_p1_2_), .IN3(
        test_so56), .QN(n12935) );
  NAND3X0 U37321 ( .IN1(s13_msel_gnt_p1[1]), .IN2(s13_msel_gnt_p1[2]), .IN3(
        s13_msel_gnt_p1[0]), .QN(n11078) );
  NAND3X0 U37322 ( .IN1(s12_msel_gnt_p1_1_), .IN2(test_so87), .IN3(
        s12_msel_gnt_p1_0_), .QN(n10768) );
  NAND3X0 U37323 ( .IN1(s3_msel_gnt_p1[1]), .IN2(s3_msel_gnt_p1[2]), .IN3(
        s3_msel_gnt_p1[0]), .QN(n12626) );
  NAND3X0 U37324 ( .IN1(s2_msel_gnt_p1[1]), .IN2(s2_msel_gnt_p1[2]), .IN3(
        s2_msel_gnt_p1[0]), .QN(n12317) );
  NAND3X0 U37325 ( .IN1(test_so83), .IN2(s11_msel_gnt_p1_2_), .IN3(
        s11_msel_gnt_p1_0_), .QN(n10459) );
  NAND3X0 U37326 ( .IN1(s10_msel_gnt_p1_1_), .IN2(s10_msel_gnt_p1_2_), .IN3(
        test_so79), .QN(n10149) );
  NAND3X0 U37327 ( .IN1(s1_msel_gnt_p1[1]), .IN2(s1_msel_gnt_p1[2]), .IN3(
        s1_msel_gnt_p1[0]), .QN(n12007) );
  NAND3X0 U37328 ( .IN1(s0_msel_gnt_p1_1_), .IN2(test_so41), .IN3(
        s0_msel_gnt_p1_0_), .QN(n11697) );
  NAND3X0 U37329 ( .IN1(s9_msel_gnt_p1[1]), .IN2(s9_msel_gnt_p1[2]), .IN3(
        s9_msel_gnt_p1[0]), .QN(n9839) );
  NAND3X0 U37330 ( .IN1(s8_msel_gnt_p1[1]), .IN2(s8_msel_gnt_p1[2]), .IN3(
        s8_msel_gnt_p1[0]), .QN(n9528) );
  NAND3X0 U37331 ( .IN1(s15_msel_gnt_p1[1]), .IN2(s15_msel_gnt_p1[2]), .IN3(
        s15_msel_gnt_p1[0]), .QN(n13995) );
  NAND4X0 U37332 ( .IN1(m7s7_cyc), .IN2(n13657), .IN3(n13658), .IN4(n13659), 
        .QN(n13656) );
  NAND4X0 U37333 ( .IN1(test_so24), .IN2(n13641), .IN3(n13642), .IN4(n13643), 
        .QN(n13640) );
  NAND4X0 U37334 ( .IN1(m7s6_cyc), .IN2(n13348), .IN3(n13349), .IN4(n13350), 
        .QN(n13347) );
  NAND4X0 U37335 ( .IN1(m3s6_cyc), .IN2(n13332), .IN3(n13333), .IN4(n13334), 
        .QN(n13331) );
  NAND4X0 U37336 ( .IN1(m7s14_cyc), .IN2(n11182), .IN3(n11183), .IN4(n11184), 
        .QN(n11181) );
  NAND4X0 U37337 ( .IN1(test_so25), .IN2(n11166), .IN3(n11167), .IN4(n11168), 
        .QN(n11165) );
  NAND4X0 U37338 ( .IN1(test_so34), .IN2(n13039), .IN3(n13040), .IN4(n13041), 
        .QN(n13038) );
  NAND4X0 U37339 ( .IN1(m3s5_cyc), .IN2(n13023), .IN3(n13024), .IN4(n13025), 
        .QN(n13022) );
  NAND4X0 U37340 ( .IN1(m7s4_cyc), .IN2(n12730), .IN3(n12731), .IN4(n12732), 
        .QN(n12729) );
  NAND4X0 U37341 ( .IN1(m3s4_cyc), .IN2(n12714), .IN3(n12715), .IN4(n12716), 
        .QN(n12713) );
  NAND4X0 U37342 ( .IN1(m7s13_cyc), .IN2(n10873), .IN3(n10874), .IN4(n10875), 
        .QN(n10872) );
  NAND4X0 U37343 ( .IN1(m3s13_cyc), .IN2(n10857), .IN3(n10858), .IN4(n10859), 
        .QN(n10856) );
  NAND4X0 U37344 ( .IN1(m7s12_cyc), .IN2(n10563), .IN3(n10564), .IN4(n10565), 
        .QN(n10562) );
  NAND4X0 U37345 ( .IN1(m3s12_cyc), .IN2(n10547), .IN3(n10548), .IN4(n10549), 
        .QN(n10546) );
  NAND4X0 U37346 ( .IN1(m7s3_cyc), .IN2(n12421), .IN3(n12422), .IN4(n12423), 
        .QN(n12420) );
  NAND4X0 U37347 ( .IN1(m3s3_cyc), .IN2(n12405), .IN3(n12406), .IN4(n12407), 
        .QN(n12404) );
  NAND4X0 U37348 ( .IN1(m7s2_cyc), .IN2(n12112), .IN3(n12113), .IN4(n12114), 
        .QN(n12111) );
  NAND4X0 U37349 ( .IN1(m3s2_cyc), .IN2(n12096), .IN3(n12097), .IN4(n12098), 
        .QN(n12095) );
  NAND4X0 U37350 ( .IN1(test_so35), .IN2(n10254), .IN3(n10255), .IN4(n10256), 
        .QN(n10253) );
  NAND4X0 U37351 ( .IN1(m3s11_cyc), .IN2(n10238), .IN3(n10239), .IN4(n10240), 
        .QN(n10237) );
  NAND4X0 U37352 ( .IN1(m7s10_cyc), .IN2(n9944), .IN3(n9945), .IN4(n9946), 
        .QN(n9943) );
  NAND4X0 U37353 ( .IN1(m3s10_cyc), .IN2(n9928), .IN3(n9929), .IN4(n9930), 
        .QN(n9927) );
  NAND4X0 U37354 ( .IN1(m7s1_cyc), .IN2(n11802), .IN3(n11803), .IN4(n11804), 
        .QN(n11801) );
  NAND4X0 U37355 ( .IN1(m3s1_cyc), .IN2(n11786), .IN3(n11787), .IN4(n11788), 
        .QN(n11785) );
  NAND4X0 U37356 ( .IN1(m7s0_cyc), .IN2(n11492), .IN3(n11493), .IN4(n11494), 
        .QN(n11491) );
  NAND4X0 U37357 ( .IN1(test_so23), .IN2(n11476), .IN3(n11477), .IN4(n11478), 
        .QN(n11475) );
  NAND4X0 U37358 ( .IN1(m7s9_cyc), .IN2(n9634), .IN3(n9635), .IN4(n9636), .QN(
        n9633) );
  NAND4X0 U37359 ( .IN1(m3s9_cyc), .IN2(n9618), .IN3(n9619), .IN4(n9620), .QN(
        n9617) );
  NAND4X0 U37360 ( .IN1(m7s8_cyc), .IN2(n9323), .IN3(n9324), .IN4(n9325), .QN(
        n9322) );
  NAND4X0 U37361 ( .IN1(m3s8_cyc), .IN2(n9307), .IN3(n9308), .IN4(n9309), .QN(
        n9306) );
  NAND4X0 U37362 ( .IN1(m7s15_cyc), .IN2(n14298), .IN3(n14069), .IN4(n14280), 
        .QN(n14297) );
  NAND4X0 U37363 ( .IN1(m3s15_cyc), .IN2(n14290), .IN3(n14073), .IN4(n14276), 
        .QN(n14289) );
  NAND4X0 U37364 ( .IN1(m6s7_cyc), .IN2(n13660), .IN3(n13661), .IN4(n13662), 
        .QN(n13655) );
  NAND4X0 U37365 ( .IN1(m2s7_cyc), .IN2(n13644), .IN3(n13645), .IN4(n13646), 
        .QN(n13639) );
  NAND4X0 U37366 ( .IN1(m6s6_cyc), .IN2(n13351), .IN3(n13352), .IN4(n13353), 
        .QN(n13346) );
  NAND4X0 U37367 ( .IN1(m2s6_cyc), .IN2(n13335), .IN3(n13336), .IN4(n13337), 
        .QN(n13330) );
  NAND4X0 U37368 ( .IN1(m6s14_cyc), .IN2(n11185), .IN3(n11186), .IN4(n11187), 
        .QN(n11180) );
  NAND4X0 U37369 ( .IN1(m2s14_cyc), .IN2(n11169), .IN3(n11170), .IN4(n11171), 
        .QN(n11164) );
  NAND4X0 U37370 ( .IN1(m6s5_cyc), .IN2(n13042), .IN3(n13043), .IN4(n13044), 
        .QN(n13037) );
  NAND4X0 U37371 ( .IN1(m2s5_cyc), .IN2(n13026), .IN3(n13027), .IN4(n13028), 
        .QN(n13021) );
  NAND4X0 U37372 ( .IN1(m6s4_cyc), .IN2(n12733), .IN3(n12734), .IN4(n12735), 
        .QN(n12728) );
  NAND4X0 U37373 ( .IN1(m2s4_cyc), .IN2(n12717), .IN3(n12718), .IN4(n12719), 
        .QN(n12712) );
  NAND4X0 U37374 ( .IN1(m6s13_cyc), .IN2(n10876), .IN3(n10877), .IN4(n10878), 
        .QN(n10871) );
  NAND4X0 U37375 ( .IN1(m2s13_cyc), .IN2(n10860), .IN3(n10861), .IN4(n10862), 
        .QN(n10855) );
  NAND4X0 U37376 ( .IN1(m6s12_cyc), .IN2(n10566), .IN3(n10567), .IN4(n10568), 
        .QN(n10561) );
  NAND4X0 U37377 ( .IN1(m2s12_cyc), .IN2(n10550), .IN3(n10551), .IN4(n10552), 
        .QN(n10545) );
  NAND4X0 U37378 ( .IN1(test_so31), .IN2(n12424), .IN3(n12425), .IN4(n12426), 
        .QN(n12419) );
  NAND4X0 U37379 ( .IN1(m2s3_cyc), .IN2(n12408), .IN3(n12409), .IN4(n12410), 
        .QN(n12403) );
  NAND4X0 U37380 ( .IN1(m6s2_cyc), .IN2(n12115), .IN3(n12116), .IN4(n12117), 
        .QN(n12110) );
  NAND4X0 U37381 ( .IN1(test_so21), .IN2(n12099), .IN3(n12100), .IN4(n12101), 
        .QN(n12094) );
  NAND4X0 U37382 ( .IN1(m6s11_cyc), .IN2(n10257), .IN3(n10258), .IN4(n10259), 
        .QN(n10252) );
  NAND4X0 U37383 ( .IN1(m2s11_cyc), .IN2(n10241), .IN3(n10242), .IN4(n10243), 
        .QN(n10236) );
  NAND4X0 U37384 ( .IN1(m6s10_cyc), .IN2(n9947), .IN3(n9948), .IN4(n9949), 
        .QN(n9942) );
  NAND4X0 U37385 ( .IN1(m2s10_cyc), .IN2(n9931), .IN3(n9932), .IN4(n9933), 
        .QN(n9926) );
  NAND4X0 U37386 ( .IN1(m6s1_cyc), .IN2(n11805), .IN3(n11806), .IN4(n11807), 
        .QN(n11800) );
  NAND4X0 U37387 ( .IN1(m2s1_cyc), .IN2(n11789), .IN3(n11790), .IN4(n11791), 
        .QN(n11784) );
  NAND4X0 U37388 ( .IN1(m6s0_cyc), .IN2(n11495), .IN3(n11496), .IN4(n11497), 
        .QN(n11490) );
  NAND4X0 U37389 ( .IN1(m2s0_cyc), .IN2(n11479), .IN3(n11480), .IN4(n11481), 
        .QN(n11474) );
  NAND4X0 U37390 ( .IN1(test_so32), .IN2(n9637), .IN3(n9638), .IN4(n9639), 
        .QN(n9632) );
  NAND4X0 U37391 ( .IN1(test_so22), .IN2(n9621), .IN3(n9622), .IN4(n9623), 
        .QN(n9616) );
  NAND4X0 U37392 ( .IN1(m6s8_cyc), .IN2(n9326), .IN3(n9327), .IN4(n9328), .QN(
        n9321) );
  NAND4X0 U37393 ( .IN1(m2s8_cyc), .IN2(n9310), .IN3(n9311), .IN4(n9312), .QN(
        n9305) );
  NAND4X0 U37394 ( .IN1(test_so33), .IN2(n14299), .IN3(n14068), .IN4(n14283), 
        .QN(n14296) );
  NAND4X0 U37395 ( .IN1(m2s15_cyc), .IN2(n14291), .IN3(n14072), .IN4(n14279), 
        .QN(n14288) );
  NAND4X0 U37396 ( .IN1(m1s7_cyc), .IN2(n13647), .IN3(n13648), .IN4(n13649), 
        .QN(n13638) );
  NAND4X0 U37397 ( .IN1(m1s6_cyc), .IN2(n13338), .IN3(n13339), .IN4(n13340), 
        .QN(n13329) );
  NAND4X0 U37398 ( .IN1(m1s14_cyc), .IN2(n11172), .IN3(n11173), .IN4(n11174), 
        .QN(n11163) );
  NAND4X0 U37399 ( .IN1(m1s5_cyc), .IN2(n13029), .IN3(n13030), .IN4(n13031), 
        .QN(n13020) );
  NAND4X0 U37400 ( .IN1(test_so19), .IN2(n12720), .IN3(n12721), .IN4(n12722), 
        .QN(n12711) );
  NAND4X0 U37401 ( .IN1(m1s13_cyc), .IN2(n10863), .IN3(n10864), .IN4(n10865), 
        .QN(n10854) );
  NAND4X0 U37402 ( .IN1(m1s12_cyc), .IN2(n10553), .IN3(n10554), .IN4(n10555), 
        .QN(n10544) );
  NAND4X0 U37403 ( .IN1(m1s3_cyc), .IN2(n12411), .IN3(n12412), .IN4(n12413), 
        .QN(n12402) );
  NAND4X0 U37404 ( .IN1(m1s2_cyc), .IN2(n12102), .IN3(n12103), .IN4(n12104), 
        .QN(n12093) );
  NAND4X0 U37405 ( .IN1(test_so20), .IN2(n10244), .IN3(n10245), .IN4(n10246), 
        .QN(n10235) );
  NAND4X0 U37406 ( .IN1(m1s10_cyc), .IN2(n9934), .IN3(n9935), .IN4(n9936), 
        .QN(n9925) );
  NAND4X0 U37407 ( .IN1(m1s1_cyc), .IN2(n11792), .IN3(n11793), .IN4(n11794), 
        .QN(n11783) );
  NAND4X0 U37408 ( .IN1(m1s0_cyc), .IN2(n11482), .IN3(n11483), .IN4(n11484), 
        .QN(n11473) );
  NAND4X0 U37409 ( .IN1(m1s9_cyc), .IN2(n9624), .IN3(n9625), .IN4(n9626), .QN(
        n9615) );
  NAND4X0 U37410 ( .IN1(m1s8_cyc), .IN2(n9313), .IN3(n9314), .IN4(n9315), .QN(
        n9304) );
  NAND4X0 U37411 ( .IN1(m1s15_cyc), .IN2(n14292), .IN3(n14075), .IN4(n14278), 
        .QN(n14287) );
  INVX0 U37412 ( .IN(s1_rty_i), .QN(n2381) );
  INVX0 U37413 ( .IN(s9_rty_i), .QN(n2661) );
  INVX0 U37414 ( .IN(s3_rty_i), .QN(n2451) );
  INVX0 U37415 ( .IN(s10_rty_i), .QN(n2696) );
  INVX0 U37416 ( .IN(s1_err_i), .QN(n2380) );
  INVX0 U37417 ( .IN(s9_err_i), .QN(n2660) );
  INVX0 U37418 ( .IN(s3_err_i), .QN(n2450) );
  INVX0 U37419 ( .IN(s10_err_i), .QN(n2695) );
  INVX0 U37420 ( .IN(s1_ack_i), .QN(n2379) );
  INVX0 U37421 ( .IN(s9_ack_i), .QN(n2659) );
  INVX0 U37422 ( .IN(s3_ack_i), .QN(n2449) );
  INVX0 U37423 ( .IN(s10_ack_i), .QN(n2694) );
  INVX0 U37424 ( .IN(s9_data_i[0]), .QN(n2658) );
  INVX0 U37425 ( .IN(s5_data_i[0]), .QN(n2518) );
  INVX0 U37426 ( .IN(s3_data_i[0]), .QN(n2448) );
  INVX0 U37427 ( .IN(s9_data_i[1]), .QN(n2657) );
  INVX0 U37428 ( .IN(s5_data_i[1]), .QN(n2517) );
  INVX0 U37429 ( .IN(s3_data_i[1]), .QN(n2447) );
  INVX0 U37430 ( .IN(s9_data_i[2]), .QN(n2656) );
  INVX0 U37431 ( .IN(s5_data_i[2]), .QN(n2516) );
  INVX0 U37432 ( .IN(s3_data_i[2]), .QN(n2446) );
  INVX0 U37433 ( .IN(s9_data_i[3]), .QN(n2655) );
  INVX0 U37434 ( .IN(s5_data_i[3]), .QN(n2515) );
  INVX0 U37435 ( .IN(s3_data_i[3]), .QN(n2445) );
  INVX0 U37436 ( .IN(s9_data_i[4]), .QN(n2654) );
  INVX0 U37437 ( .IN(s5_data_i[4]), .QN(n2514) );
  INVX0 U37438 ( .IN(s3_data_i[4]), .QN(n2444) );
  INVX0 U37439 ( .IN(s9_data_i[5]), .QN(n2653) );
  INVX0 U37440 ( .IN(s5_data_i[5]), .QN(n2513) );
  INVX0 U37441 ( .IN(s3_data_i[5]), .QN(n2443) );
  INVX0 U37442 ( .IN(s9_data_i[6]), .QN(n2652) );
  INVX0 U37443 ( .IN(s5_data_i[6]), .QN(n2512) );
  INVX0 U37444 ( .IN(s3_data_i[6]), .QN(n2442) );
  INVX0 U37445 ( .IN(s9_data_i[7]), .QN(n2651) );
  INVX0 U37446 ( .IN(s5_data_i[7]), .QN(n2511) );
  INVX0 U37447 ( .IN(s3_data_i[7]), .QN(n2441) );
  INVX0 U37448 ( .IN(s9_data_i[8]), .QN(n2650) );
  INVX0 U37449 ( .IN(s5_data_i[8]), .QN(n2510) );
  INVX0 U37450 ( .IN(s3_data_i[8]), .QN(n2440) );
  INVX0 U37451 ( .IN(s9_data_i[9]), .QN(n2649) );
  INVX0 U37452 ( .IN(s5_data_i[9]), .QN(n2509) );
  INVX0 U37453 ( .IN(s3_data_i[9]), .QN(n2439) );
  INVX0 U37454 ( .IN(s9_data_i[10]), .QN(n2648) );
  INVX0 U37455 ( .IN(s5_data_i[10]), .QN(n2508) );
  INVX0 U37456 ( .IN(s3_data_i[10]), .QN(n2438) );
  INVX0 U37457 ( .IN(s9_data_i[11]), .QN(n2647) );
  INVX0 U37458 ( .IN(s5_data_i[11]), .QN(n2507) );
  INVX0 U37459 ( .IN(s3_data_i[11]), .QN(n2437) );
  INVX0 U37460 ( .IN(s9_data_i[12]), .QN(n2646) );
  INVX0 U37461 ( .IN(s5_data_i[12]), .QN(n2506) );
  INVX0 U37462 ( .IN(s3_data_i[12]), .QN(n2436) );
  INVX0 U37463 ( .IN(s9_data_i[13]), .QN(n2645) );
  INVX0 U37464 ( .IN(s5_data_i[13]), .QN(n2505) );
  INVX0 U37465 ( .IN(s3_data_i[13]), .QN(n2435) );
  INVX0 U37466 ( .IN(s9_data_i[14]), .QN(n2644) );
  INVX0 U37467 ( .IN(s5_data_i[14]), .QN(n2504) );
  INVX0 U37468 ( .IN(s3_data_i[14]), .QN(n2434) );
  INVX0 U37469 ( .IN(s9_data_i[15]), .QN(n2643) );
  INVX0 U37470 ( .IN(s5_data_i[15]), .QN(n2503) );
  INVX0 U37471 ( .IN(s3_data_i[15]), .QN(n2433) );
  INVX0 U37472 ( .IN(s9_data_i[16]), .QN(n2642) );
  INVX0 U37473 ( .IN(s5_data_i[16]), .QN(n2502) );
  INVX0 U37474 ( .IN(s3_data_i[16]), .QN(n2432) );
  INVX0 U37475 ( .IN(s9_data_i[17]), .QN(n2641) );
  INVX0 U37476 ( .IN(s5_data_i[17]), .QN(n2501) );
  INVX0 U37477 ( .IN(s3_data_i[17]), .QN(n2431) );
  INVX0 U37478 ( .IN(s9_data_i[18]), .QN(n2640) );
  INVX0 U37479 ( .IN(s5_data_i[18]), .QN(n2500) );
  INVX0 U37480 ( .IN(s3_data_i[18]), .QN(n2430) );
  INVX0 U37481 ( .IN(s9_data_i[19]), .QN(n2639) );
  INVX0 U37482 ( .IN(s5_data_i[19]), .QN(n2499) );
  INVX0 U37483 ( .IN(s3_data_i[19]), .QN(n2429) );
  INVX0 U37484 ( .IN(s9_data_i[20]), .QN(n2638) );
  INVX0 U37485 ( .IN(s5_data_i[20]), .QN(n2498) );
  INVX0 U37486 ( .IN(s3_data_i[20]), .QN(n2428) );
  INVX0 U37487 ( .IN(s9_data_i[21]), .QN(n2637) );
  INVX0 U37488 ( .IN(s5_data_i[21]), .QN(n2497) );
  INVX0 U37489 ( .IN(s3_data_i[21]), .QN(n2427) );
  INVX0 U37490 ( .IN(s9_data_i[22]), .QN(n2636) );
  INVX0 U37491 ( .IN(s5_data_i[22]), .QN(n2496) );
  INVX0 U37492 ( .IN(s3_data_i[22]), .QN(n2426) );
  INVX0 U37493 ( .IN(s9_data_i[23]), .QN(n2635) );
  INVX0 U37494 ( .IN(s5_data_i[23]), .QN(n2495) );
  INVX0 U37495 ( .IN(s3_data_i[23]), .QN(n2425) );
  INVX0 U37496 ( .IN(s9_data_i[24]), .QN(n2634) );
  INVX0 U37497 ( .IN(s5_data_i[24]), .QN(n2494) );
  INVX0 U37498 ( .IN(s3_data_i[24]), .QN(n2424) );
  INVX0 U37499 ( .IN(s9_data_i[25]), .QN(n2633) );
  INVX0 U37500 ( .IN(s5_data_i[25]), .QN(n2493) );
  INVX0 U37501 ( .IN(s3_data_i[25]), .QN(n2423) );
  INVX0 U37502 ( .IN(s9_data_i[26]), .QN(n2632) );
  INVX0 U37503 ( .IN(s5_data_i[26]), .QN(n2492) );
  INVX0 U37504 ( .IN(s3_data_i[26]), .QN(n2422) );
  INVX0 U37505 ( .IN(s9_data_i[27]), .QN(n2631) );
  INVX0 U37506 ( .IN(s5_data_i[27]), .QN(n2491) );
  INVX0 U37507 ( .IN(s3_data_i[27]), .QN(n2421) );
  INVX0 U37508 ( .IN(s9_data_i[28]), .QN(n2630) );
  INVX0 U37509 ( .IN(s5_data_i[28]), .QN(n2490) );
  INVX0 U37510 ( .IN(s3_data_i[28]), .QN(n2420) );
  INVX0 U37511 ( .IN(s9_data_i[29]), .QN(n2629) );
  INVX0 U37512 ( .IN(s5_data_i[29]), .QN(n2489) );
  INVX0 U37513 ( .IN(s3_data_i[29]), .QN(n2419) );
  INVX0 U37514 ( .IN(s9_data_i[30]), .QN(n2628) );
  INVX0 U37515 ( .IN(s5_data_i[30]), .QN(n2488) );
  INVX0 U37516 ( .IN(s3_data_i[30]), .QN(n2418) );
  INVX0 U37517 ( .IN(s9_data_i[31]), .QN(n2627) );
  INVX0 U37518 ( .IN(s5_data_i[31]), .QN(n2487) );
  INVX0 U37519 ( .IN(s3_data_i[31]), .QN(n2417) );
  INVX0 U37520 ( .IN(s8_rty_i), .QN(n2626) );
  INVX0 U37521 ( .IN(s2_rty_i), .QN(n2416) );
  INVX0 U37522 ( .IN(s0_rty_i), .QN(n2346) );
  INVX0 U37523 ( .IN(s8_err_i), .QN(n2625) );
  INVX0 U37524 ( .IN(s2_err_i), .QN(n2415) );
  INVX0 U37525 ( .IN(s0_err_i), .QN(n2345) );
  INVX0 U37526 ( .IN(s8_ack_i), .QN(n2624) );
  INVX0 U37527 ( .IN(s2_ack_i), .QN(n2414) );
  INVX0 U37528 ( .IN(s0_ack_i), .QN(n2344) );
  INVX0 U37529 ( .IN(s14_data_i[0]), .QN(n2833) );
  INVX0 U37530 ( .IN(s8_data_i[0]), .QN(n2623) );
  INVX0 U37531 ( .IN(s4_data_i[0]), .QN(n2483) );
  INVX0 U37532 ( .IN(s2_data_i[0]), .QN(n2413) );
  INVX0 U37533 ( .IN(s14_data_i[1]), .QN(n2832) );
  INVX0 U37534 ( .IN(s8_data_i[1]), .QN(n2622) );
  INVX0 U37535 ( .IN(s4_data_i[1]), .QN(n2482) );
  INVX0 U37536 ( .IN(s2_data_i[1]), .QN(n2412) );
  INVX0 U37537 ( .IN(s14_data_i[2]), .QN(n2831) );
  INVX0 U37538 ( .IN(s8_data_i[2]), .QN(n2621) );
  INVX0 U37539 ( .IN(s4_data_i[2]), .QN(n2481) );
  INVX0 U37540 ( .IN(s2_data_i[2]), .QN(n2411) );
  INVX0 U37541 ( .IN(s14_data_i[3]), .QN(n2830) );
  INVX0 U37542 ( .IN(s8_data_i[3]), .QN(n2620) );
  INVX0 U37543 ( .IN(s4_data_i[3]), .QN(n2480) );
  INVX0 U37544 ( .IN(s2_data_i[3]), .QN(n2410) );
  INVX0 U37545 ( .IN(s14_data_i[4]), .QN(n2829) );
  INVX0 U37546 ( .IN(s8_data_i[4]), .QN(n2619) );
  INVX0 U37547 ( .IN(s4_data_i[4]), .QN(n2479) );
  INVX0 U37548 ( .IN(s2_data_i[4]), .QN(n2409) );
  INVX0 U37549 ( .IN(s14_data_i[5]), .QN(n2828) );
  INVX0 U37550 ( .IN(s8_data_i[5]), .QN(n2618) );
  INVX0 U37551 ( .IN(s4_data_i[5]), .QN(n2478) );
  INVX0 U37552 ( .IN(s2_data_i[5]), .QN(n2408) );
  INVX0 U37553 ( .IN(s14_data_i[6]), .QN(n2827) );
  INVX0 U37554 ( .IN(s8_data_i[6]), .QN(n2617) );
  INVX0 U37555 ( .IN(s4_data_i[6]), .QN(n2477) );
  INVX0 U37556 ( .IN(s2_data_i[6]), .QN(n2407) );
  INVX0 U37557 ( .IN(s14_data_i[7]), .QN(n2826) );
  INVX0 U37558 ( .IN(s8_data_i[7]), .QN(n2616) );
  INVX0 U37559 ( .IN(s4_data_i[7]), .QN(n2476) );
  INVX0 U37560 ( .IN(s2_data_i[7]), .QN(n2406) );
  INVX0 U37561 ( .IN(s14_data_i[8]), .QN(n2825) );
  INVX0 U37562 ( .IN(s8_data_i[8]), .QN(n2615) );
  INVX0 U37563 ( .IN(s4_data_i[8]), .QN(n2475) );
  INVX0 U37564 ( .IN(s2_data_i[8]), .QN(n2405) );
  INVX0 U37565 ( .IN(s14_data_i[9]), .QN(n2824) );
  INVX0 U37566 ( .IN(s8_data_i[9]), .QN(n2614) );
  INVX0 U37567 ( .IN(s4_data_i[9]), .QN(n2474) );
  INVX0 U37568 ( .IN(s2_data_i[9]), .QN(n2404) );
  INVX0 U37569 ( .IN(s14_data_i[10]), .QN(n2823) );
  INVX0 U37570 ( .IN(s8_data_i[10]), .QN(n2613) );
  INVX0 U37571 ( .IN(s4_data_i[10]), .QN(n2473) );
  INVX0 U37572 ( .IN(s2_data_i[10]), .QN(n2403) );
  INVX0 U37573 ( .IN(s14_data_i[11]), .QN(n2822) );
  INVX0 U37574 ( .IN(s8_data_i[11]), .QN(n2612) );
  INVX0 U37575 ( .IN(s4_data_i[11]), .QN(n2472) );
  INVX0 U37576 ( .IN(s2_data_i[11]), .QN(n2402) );
  INVX0 U37577 ( .IN(s14_data_i[12]), .QN(n2821) );
  INVX0 U37578 ( .IN(s8_data_i[12]), .QN(n2611) );
  INVX0 U37579 ( .IN(s4_data_i[12]), .QN(n2471) );
  INVX0 U37580 ( .IN(s2_data_i[12]), .QN(n2401) );
  INVX0 U37581 ( .IN(s14_data_i[13]), .QN(n2820) );
  INVX0 U37582 ( .IN(s8_data_i[13]), .QN(n2610) );
  INVX0 U37583 ( .IN(s4_data_i[13]), .QN(n2470) );
  INVX0 U37584 ( .IN(s2_data_i[13]), .QN(n2400) );
  INVX0 U37585 ( .IN(s14_data_i[14]), .QN(n2819) );
  INVX0 U37586 ( .IN(s8_data_i[14]), .QN(n2609) );
  INVX0 U37587 ( .IN(s4_data_i[14]), .QN(n2469) );
  INVX0 U37588 ( .IN(s2_data_i[14]), .QN(n2399) );
  INVX0 U37589 ( .IN(s14_data_i[15]), .QN(n2818) );
  INVX0 U37590 ( .IN(s8_data_i[15]), .QN(n2608) );
  INVX0 U37591 ( .IN(s4_data_i[15]), .QN(n2468) );
  INVX0 U37592 ( .IN(s2_data_i[15]), .QN(n2398) );
  INVX0 U37593 ( .IN(s14_data_i[16]), .QN(n2817) );
  INVX0 U37594 ( .IN(s8_data_i[16]), .QN(n2607) );
  INVX0 U37595 ( .IN(s4_data_i[16]), .QN(n2467) );
  INVX0 U37596 ( .IN(s2_data_i[16]), .QN(n2397) );
  INVX0 U37597 ( .IN(s14_data_i[17]), .QN(n2816) );
  INVX0 U37598 ( .IN(s8_data_i[17]), .QN(n2606) );
  INVX0 U37599 ( .IN(s4_data_i[17]), .QN(n2466) );
  INVX0 U37600 ( .IN(s2_data_i[17]), .QN(n2396) );
  INVX0 U37601 ( .IN(s14_data_i[18]), .QN(n2815) );
  INVX0 U37602 ( .IN(s8_data_i[18]), .QN(n2605) );
  INVX0 U37603 ( .IN(s4_data_i[18]), .QN(n2465) );
  INVX0 U37604 ( .IN(s2_data_i[18]), .QN(n2395) );
  INVX0 U37605 ( .IN(s14_data_i[19]), .QN(n2814) );
  INVX0 U37606 ( .IN(s8_data_i[19]), .QN(n2604) );
  INVX0 U37607 ( .IN(s4_data_i[19]), .QN(n2464) );
  INVX0 U37608 ( .IN(s2_data_i[19]), .QN(n2394) );
  INVX0 U37609 ( .IN(s14_data_i[20]), .QN(n2813) );
  INVX0 U37610 ( .IN(s8_data_i[20]), .QN(n2603) );
  INVX0 U37611 ( .IN(s4_data_i[20]), .QN(n2463) );
  INVX0 U37612 ( .IN(s2_data_i[20]), .QN(n2393) );
  INVX0 U37613 ( .IN(s14_data_i[21]), .QN(n2812) );
  INVX0 U37614 ( .IN(s8_data_i[21]), .QN(n2602) );
  INVX0 U37615 ( .IN(s4_data_i[21]), .QN(n2462) );
  INVX0 U37616 ( .IN(s2_data_i[21]), .QN(n2392) );
  INVX0 U37617 ( .IN(s14_data_i[22]), .QN(n2811) );
  INVX0 U37618 ( .IN(s8_data_i[22]), .QN(n2601) );
  INVX0 U37619 ( .IN(s4_data_i[22]), .QN(n2461) );
  INVX0 U37620 ( .IN(s2_data_i[22]), .QN(n2391) );
  INVX0 U37621 ( .IN(s14_data_i[23]), .QN(n2810) );
  INVX0 U37622 ( .IN(s8_data_i[23]), .QN(n2600) );
  INVX0 U37623 ( .IN(s4_data_i[23]), .QN(n2460) );
  INVX0 U37624 ( .IN(s2_data_i[23]), .QN(n2390) );
  INVX0 U37625 ( .IN(s14_data_i[24]), .QN(n2809) );
  INVX0 U37626 ( .IN(s8_data_i[24]), .QN(n2599) );
  INVX0 U37627 ( .IN(s4_data_i[24]), .QN(n2459) );
  INVX0 U37628 ( .IN(s2_data_i[24]), .QN(n2389) );
  INVX0 U37629 ( .IN(s14_data_i[25]), .QN(n2808) );
  INVX0 U37630 ( .IN(s8_data_i[25]), .QN(n2598) );
  INVX0 U37631 ( .IN(s4_data_i[25]), .QN(n2458) );
  INVX0 U37632 ( .IN(s2_data_i[25]), .QN(n2388) );
  INVX0 U37633 ( .IN(s14_data_i[26]), .QN(n2807) );
  INVX0 U37634 ( .IN(s8_data_i[26]), .QN(n2597) );
  INVX0 U37635 ( .IN(s4_data_i[26]), .QN(n2457) );
  INVX0 U37636 ( .IN(s2_data_i[26]), .QN(n2387) );
  INVX0 U37637 ( .IN(s14_data_i[27]), .QN(n2806) );
  INVX0 U37638 ( .IN(s8_data_i[27]), .QN(n2596) );
  INVX0 U37639 ( .IN(s4_data_i[27]), .QN(n2456) );
  INVX0 U37640 ( .IN(s2_data_i[27]), .QN(n2386) );
  INVX0 U37641 ( .IN(s14_data_i[28]), .QN(n2805) );
  INVX0 U37642 ( .IN(s8_data_i[28]), .QN(n2595) );
  INVX0 U37643 ( .IN(s4_data_i[28]), .QN(n2455) );
  INVX0 U37644 ( .IN(s2_data_i[28]), .QN(n2385) );
  INVX0 U37645 ( .IN(s14_data_i[29]), .QN(n2804) );
  INVX0 U37646 ( .IN(s8_data_i[29]), .QN(n2594) );
  INVX0 U37647 ( .IN(s4_data_i[29]), .QN(n2454) );
  INVX0 U37648 ( .IN(s2_data_i[29]), .QN(n2384) );
  INVX0 U37649 ( .IN(s14_data_i[30]), .QN(n2803) );
  INVX0 U37650 ( .IN(s8_data_i[30]), .QN(n2593) );
  INVX0 U37651 ( .IN(s4_data_i[30]), .QN(n2453) );
  INVX0 U37652 ( .IN(s2_data_i[30]), .QN(n2383) );
  INVX0 U37653 ( .IN(s14_data_i[31]), .QN(n2802) );
  INVX0 U37654 ( .IN(s8_data_i[31]), .QN(n2592) );
  INVX0 U37655 ( .IN(s4_data_i[31]), .QN(n2452) );
  INVX0 U37656 ( .IN(s2_data_i[31]), .QN(n2382) );
  INVX0 U37657 ( .IN(s14_rty_i), .QN(n2836) );
  INVX0 U37658 ( .IN(s7_rty_i), .QN(n2591) );
  INVX0 U37659 ( .IN(s5_rty_i), .QN(n2521) );
  INVX0 U37660 ( .IN(s12_rty_i), .QN(n2766) );
  INVX0 U37661 ( .IN(s14_err_i), .QN(n2835) );
  INVX0 U37662 ( .IN(s7_err_i), .QN(n2590) );
  INVX0 U37663 ( .IN(s5_err_i), .QN(n2520) );
  INVX0 U37664 ( .IN(s12_err_i), .QN(n2765) );
  INVX0 U37665 ( .IN(s14_ack_i), .QN(n2834) );
  INVX0 U37666 ( .IN(s7_ack_i), .QN(n2589) );
  INVX0 U37667 ( .IN(s5_ack_i), .QN(n2519) );
  INVX0 U37668 ( .IN(s12_ack_i), .QN(n2764) );
  INVX0 U37669 ( .IN(s13_data_i[0]), .QN(n2798) );
  INVX0 U37670 ( .IN(s11_data_i[0]), .QN(n2728) );
  INVX0 U37671 ( .IN(s7_data_i[0]), .QN(n2588) );
  INVX0 U37672 ( .IN(s1_data_i[0]), .QN(n2378) );
  INVX0 U37673 ( .IN(s13_data_i[1]), .QN(n2797) );
  INVX0 U37674 ( .IN(s11_data_i[1]), .QN(n2727) );
  INVX0 U37675 ( .IN(s7_data_i[1]), .QN(n2587) );
  INVX0 U37676 ( .IN(s1_data_i[1]), .QN(n2377) );
  INVX0 U37677 ( .IN(s13_data_i[2]), .QN(n2796) );
  INVX0 U37678 ( .IN(s11_data_i[2]), .QN(n2726) );
  INVX0 U37679 ( .IN(s7_data_i[2]), .QN(n2586) );
  INVX0 U37680 ( .IN(s1_data_i[2]), .QN(n2376) );
  INVX0 U37681 ( .IN(s13_data_i[3]), .QN(n2795) );
  INVX0 U37682 ( .IN(s11_data_i[3]), .QN(n2725) );
  INVX0 U37683 ( .IN(s7_data_i[3]), .QN(n2585) );
  INVX0 U37684 ( .IN(s1_data_i[3]), .QN(n2375) );
  INVX0 U37685 ( .IN(s13_data_i[4]), .QN(n2794) );
  INVX0 U37686 ( .IN(s11_data_i[4]), .QN(n2724) );
  INVX0 U37687 ( .IN(s7_data_i[4]), .QN(n2584) );
  INVX0 U37688 ( .IN(s1_data_i[4]), .QN(n2374) );
  INVX0 U37689 ( .IN(s13_data_i[5]), .QN(n2793) );
  INVX0 U37690 ( .IN(s11_data_i[5]), .QN(n2723) );
  INVX0 U37691 ( .IN(s7_data_i[5]), .QN(n2583) );
  INVX0 U37692 ( .IN(s1_data_i[5]), .QN(n2373) );
  INVX0 U37693 ( .IN(s13_data_i[6]), .QN(n2792) );
  INVX0 U37694 ( .IN(s11_data_i[6]), .QN(n2722) );
  INVX0 U37695 ( .IN(s7_data_i[6]), .QN(n2582) );
  INVX0 U37696 ( .IN(s1_data_i[6]), .QN(n2372) );
  INVX0 U37697 ( .IN(s13_data_i[7]), .QN(n2791) );
  INVX0 U37698 ( .IN(s11_data_i[7]), .QN(n2721) );
  INVX0 U37699 ( .IN(s7_data_i[7]), .QN(n2581) );
  INVX0 U37700 ( .IN(s1_data_i[7]), .QN(n2371) );
  INVX0 U37701 ( .IN(s13_data_i[8]), .QN(n2790) );
  INVX0 U37702 ( .IN(s11_data_i[8]), .QN(n2720) );
  INVX0 U37703 ( .IN(s7_data_i[8]), .QN(n2580) );
  INVX0 U37704 ( .IN(s1_data_i[8]), .QN(n2370) );
  INVX0 U37705 ( .IN(s13_data_i[9]), .QN(n2789) );
  INVX0 U37706 ( .IN(s11_data_i[9]), .QN(n2719) );
  INVX0 U37707 ( .IN(s7_data_i[9]), .QN(n2579) );
  INVX0 U37708 ( .IN(s1_data_i[9]), .QN(n2369) );
  INVX0 U37709 ( .IN(s13_data_i[10]), .QN(n2788) );
  INVX0 U37710 ( .IN(s11_data_i[10]), .QN(n2718) );
  INVX0 U37711 ( .IN(s7_data_i[10]), .QN(n2578) );
  INVX0 U37712 ( .IN(s1_data_i[10]), .QN(n2368) );
  INVX0 U37713 ( .IN(s13_data_i[11]), .QN(n2787) );
  INVX0 U37714 ( .IN(s11_data_i[11]), .QN(n2717) );
  INVX0 U37715 ( .IN(s7_data_i[11]), .QN(n2577) );
  INVX0 U37716 ( .IN(s1_data_i[11]), .QN(n2367) );
  INVX0 U37717 ( .IN(s13_data_i[12]), .QN(n2786) );
  INVX0 U37718 ( .IN(s11_data_i[12]), .QN(n2716) );
  INVX0 U37719 ( .IN(s7_data_i[12]), .QN(n2576) );
  INVX0 U37720 ( .IN(s1_data_i[12]), .QN(n2366) );
  INVX0 U37721 ( .IN(s13_data_i[13]), .QN(n2785) );
  INVX0 U37722 ( .IN(s11_data_i[13]), .QN(n2715) );
  INVX0 U37723 ( .IN(s7_data_i[13]), .QN(n2575) );
  INVX0 U37724 ( .IN(s1_data_i[13]), .QN(n2365) );
  INVX0 U37725 ( .IN(s13_data_i[14]), .QN(n2784) );
  INVX0 U37726 ( .IN(s11_data_i[14]), .QN(n2714) );
  INVX0 U37727 ( .IN(s7_data_i[14]), .QN(n2574) );
  INVX0 U37728 ( .IN(s1_data_i[14]), .QN(n2364) );
  INVX0 U37729 ( .IN(s13_data_i[15]), .QN(n2783) );
  INVX0 U37730 ( .IN(s11_data_i[15]), .QN(n2713) );
  INVX0 U37731 ( .IN(s7_data_i[15]), .QN(n2573) );
  INVX0 U37732 ( .IN(s1_data_i[15]), .QN(n2363) );
  INVX0 U37733 ( .IN(s13_data_i[16]), .QN(n2782) );
  INVX0 U37734 ( .IN(s11_data_i[16]), .QN(n2712) );
  INVX0 U37735 ( .IN(s7_data_i[16]), .QN(n2572) );
  INVX0 U37736 ( .IN(s1_data_i[16]), .QN(n2362) );
  INVX0 U37737 ( .IN(s13_data_i[17]), .QN(n2781) );
  INVX0 U37738 ( .IN(s11_data_i[17]), .QN(n2711) );
  INVX0 U37739 ( .IN(s7_data_i[17]), .QN(n2571) );
  INVX0 U37740 ( .IN(s1_data_i[17]), .QN(n2361) );
  INVX0 U37741 ( .IN(s13_data_i[18]), .QN(n2780) );
  INVX0 U37742 ( .IN(s11_data_i[18]), .QN(n2710) );
  INVX0 U37743 ( .IN(s7_data_i[18]), .QN(n2570) );
  INVX0 U37744 ( .IN(s1_data_i[18]), .QN(n2360) );
  INVX0 U37745 ( .IN(s13_data_i[19]), .QN(n2779) );
  INVX0 U37746 ( .IN(s11_data_i[19]), .QN(n2709) );
  INVX0 U37747 ( .IN(s7_data_i[19]), .QN(n2569) );
  INVX0 U37748 ( .IN(s1_data_i[19]), .QN(n2359) );
  INVX0 U37749 ( .IN(s13_data_i[20]), .QN(n2778) );
  INVX0 U37750 ( .IN(s11_data_i[20]), .QN(n2708) );
  INVX0 U37751 ( .IN(s7_data_i[20]), .QN(n2568) );
  INVX0 U37752 ( .IN(s1_data_i[20]), .QN(n2358) );
  INVX0 U37753 ( .IN(s13_data_i[21]), .QN(n2777) );
  INVX0 U37754 ( .IN(s11_data_i[21]), .QN(n2707) );
  INVX0 U37755 ( .IN(s7_data_i[21]), .QN(n2567) );
  INVX0 U37756 ( .IN(s1_data_i[21]), .QN(n2357) );
  INVX0 U37757 ( .IN(s13_data_i[22]), .QN(n2776) );
  INVX0 U37758 ( .IN(s11_data_i[22]), .QN(n2706) );
  INVX0 U37759 ( .IN(s7_data_i[22]), .QN(n2566) );
  INVX0 U37760 ( .IN(s1_data_i[22]), .QN(n2356) );
  INVX0 U37761 ( .IN(s13_data_i[23]), .QN(n2775) );
  INVX0 U37762 ( .IN(s11_data_i[23]), .QN(n2705) );
  INVX0 U37763 ( .IN(s7_data_i[23]), .QN(n2565) );
  INVX0 U37764 ( .IN(s1_data_i[23]), .QN(n2355) );
  INVX0 U37765 ( .IN(s13_data_i[24]), .QN(n2774) );
  INVX0 U37766 ( .IN(s11_data_i[24]), .QN(n2704) );
  INVX0 U37767 ( .IN(s7_data_i[24]), .QN(n2564) );
  INVX0 U37768 ( .IN(s1_data_i[24]), .QN(n2354) );
  INVX0 U37769 ( .IN(s13_data_i[25]), .QN(n2773) );
  INVX0 U37770 ( .IN(s11_data_i[25]), .QN(n2703) );
  INVX0 U37771 ( .IN(s7_data_i[25]), .QN(n2563) );
  INVX0 U37772 ( .IN(s1_data_i[25]), .QN(n2353) );
  INVX0 U37773 ( .IN(s13_data_i[26]), .QN(n2772) );
  INVX0 U37774 ( .IN(s11_data_i[26]), .QN(n2702) );
  INVX0 U37775 ( .IN(s7_data_i[26]), .QN(n2562) );
  INVX0 U37776 ( .IN(s1_data_i[26]), .QN(n2352) );
  INVX0 U37777 ( .IN(s13_data_i[27]), .QN(n2771) );
  INVX0 U37778 ( .IN(s11_data_i[27]), .QN(n2701) );
  INVX0 U37779 ( .IN(s7_data_i[27]), .QN(n2561) );
  INVX0 U37780 ( .IN(s1_data_i[27]), .QN(n2351) );
  INVX0 U37781 ( .IN(s13_data_i[28]), .QN(n2770) );
  INVX0 U37782 ( .IN(s11_data_i[28]), .QN(n2700) );
  INVX0 U37783 ( .IN(s7_data_i[28]), .QN(n2560) );
  INVX0 U37784 ( .IN(s1_data_i[28]), .QN(n2350) );
  INVX0 U37785 ( .IN(s13_data_i[29]), .QN(n2769) );
  INVX0 U37786 ( .IN(s11_data_i[29]), .QN(n2699) );
  INVX0 U37787 ( .IN(s7_data_i[29]), .QN(n2559) );
  INVX0 U37788 ( .IN(s1_data_i[29]), .QN(n2349) );
  INVX0 U37789 ( .IN(s13_data_i[30]), .QN(n2768) );
  INVX0 U37790 ( .IN(s11_data_i[30]), .QN(n2698) );
  INVX0 U37791 ( .IN(s7_data_i[30]), .QN(n2558) );
  INVX0 U37792 ( .IN(s1_data_i[30]), .QN(n2348) );
  INVX0 U37793 ( .IN(s13_data_i[31]), .QN(n2767) );
  INVX0 U37794 ( .IN(s11_data_i[31]), .QN(n2697) );
  INVX0 U37795 ( .IN(s7_data_i[31]), .QN(n2557) );
  INVX0 U37796 ( .IN(s1_data_i[31]), .QN(n2347) );
  INVX0 U37797 ( .IN(s13_rty_i), .QN(n2801) );
  INVX0 U37798 ( .IN(s6_rty_i), .QN(n2556) );
  INVX0 U37799 ( .IN(s4_rty_i), .QN(n2486) );
  INVX0 U37800 ( .IN(s11_rty_i), .QN(n2731) );
  INVX0 U37801 ( .IN(s13_err_i), .QN(n2800) );
  INVX0 U37802 ( .IN(s6_err_i), .QN(n2555) );
  INVX0 U37803 ( .IN(s4_err_i), .QN(n2485) );
  INVX0 U37804 ( .IN(s11_err_i), .QN(n2730) );
  INVX0 U37805 ( .IN(s13_ack_i), .QN(n2799) );
  INVX0 U37806 ( .IN(s6_ack_i), .QN(n2554) );
  INVX0 U37807 ( .IN(s4_ack_i), .QN(n2484) );
  INVX0 U37808 ( .IN(s11_ack_i), .QN(n2729) );
  INVX0 U37809 ( .IN(s12_data_i[0]), .QN(n2763) );
  INVX0 U37810 ( .IN(s10_data_i[0]), .QN(n2693) );
  INVX0 U37811 ( .IN(s6_data_i[0]), .QN(n2553) );
  INVX0 U37812 ( .IN(s0_data_i[0]), .QN(n2343) );
  INVX0 U37813 ( .IN(s12_data_i[1]), .QN(n2762) );
  INVX0 U37814 ( .IN(s10_data_i[1]), .QN(n2692) );
  INVX0 U37815 ( .IN(s6_data_i[1]), .QN(n2552) );
  INVX0 U37816 ( .IN(s0_data_i[1]), .QN(n2342) );
  INVX0 U37817 ( .IN(s12_data_i[2]), .QN(n2761) );
  INVX0 U37818 ( .IN(s10_data_i[2]), .QN(n2691) );
  INVX0 U37819 ( .IN(s6_data_i[2]), .QN(n2551) );
  INVX0 U37820 ( .IN(s0_data_i[2]), .QN(n2341) );
  INVX0 U37821 ( .IN(s12_data_i[3]), .QN(n2760) );
  INVX0 U37822 ( .IN(s10_data_i[3]), .QN(n2690) );
  INVX0 U37823 ( .IN(s6_data_i[3]), .QN(n2550) );
  INVX0 U37824 ( .IN(s0_data_i[3]), .QN(n2340) );
  INVX0 U37825 ( .IN(s12_data_i[4]), .QN(n2759) );
  INVX0 U37826 ( .IN(s10_data_i[4]), .QN(n2689) );
  INVX0 U37827 ( .IN(s6_data_i[4]), .QN(n2549) );
  INVX0 U37828 ( .IN(s0_data_i[4]), .QN(n2339) );
  INVX0 U37829 ( .IN(s12_data_i[5]), .QN(n2758) );
  INVX0 U37830 ( .IN(s10_data_i[5]), .QN(n2688) );
  INVX0 U37831 ( .IN(s6_data_i[5]), .QN(n2548) );
  INVX0 U37832 ( .IN(s0_data_i[5]), .QN(n2338) );
  INVX0 U37833 ( .IN(s12_data_i[6]), .QN(n2757) );
  INVX0 U37834 ( .IN(s10_data_i[6]), .QN(n2687) );
  INVX0 U37835 ( .IN(s6_data_i[6]), .QN(n2547) );
  INVX0 U37836 ( .IN(s0_data_i[6]), .QN(n2337) );
  INVX0 U37837 ( .IN(s12_data_i[7]), .QN(n2756) );
  INVX0 U37838 ( .IN(s10_data_i[7]), .QN(n2686) );
  INVX0 U37839 ( .IN(s6_data_i[7]), .QN(n2546) );
  INVX0 U37840 ( .IN(s0_data_i[7]), .QN(n2336) );
  INVX0 U37841 ( .IN(s12_data_i[8]), .QN(n2755) );
  INVX0 U37842 ( .IN(s10_data_i[8]), .QN(n2685) );
  INVX0 U37843 ( .IN(s6_data_i[8]), .QN(n2545) );
  INVX0 U37844 ( .IN(s0_data_i[8]), .QN(n2335) );
  INVX0 U37845 ( .IN(s12_data_i[9]), .QN(n2754) );
  INVX0 U37846 ( .IN(s10_data_i[9]), .QN(n2684) );
  INVX0 U37847 ( .IN(s6_data_i[9]), .QN(n2544) );
  INVX0 U37848 ( .IN(s0_data_i[9]), .QN(n2334) );
  INVX0 U37849 ( .IN(s12_data_i[10]), .QN(n2753) );
  INVX0 U37850 ( .IN(s10_data_i[10]), .QN(n2683) );
  INVX0 U37851 ( .IN(s6_data_i[10]), .QN(n2543) );
  INVX0 U37852 ( .IN(s0_data_i[10]), .QN(n2333) );
  INVX0 U37853 ( .IN(s12_data_i[11]), .QN(n2752) );
  INVX0 U37854 ( .IN(s10_data_i[11]), .QN(n2682) );
  INVX0 U37855 ( .IN(s6_data_i[11]), .QN(n2542) );
  INVX0 U37856 ( .IN(s0_data_i[11]), .QN(n2332) );
  INVX0 U37857 ( .IN(s12_data_i[12]), .QN(n2751) );
  INVX0 U37858 ( .IN(s10_data_i[12]), .QN(n2681) );
  INVX0 U37859 ( .IN(s6_data_i[12]), .QN(n2541) );
  INVX0 U37860 ( .IN(s0_data_i[12]), .QN(n2331) );
  INVX0 U37861 ( .IN(s12_data_i[13]), .QN(n2750) );
  INVX0 U37862 ( .IN(s10_data_i[13]), .QN(n2680) );
  INVX0 U37863 ( .IN(s6_data_i[13]), .QN(n2540) );
  INVX0 U37864 ( .IN(s0_data_i[13]), .QN(n2330) );
  INVX0 U37865 ( .IN(s12_data_i[14]), .QN(n2749) );
  INVX0 U37866 ( .IN(s10_data_i[14]), .QN(n2679) );
  INVX0 U37867 ( .IN(s6_data_i[14]), .QN(n2539) );
  INVX0 U37868 ( .IN(s0_data_i[14]), .QN(n2329) );
  INVX0 U37869 ( .IN(s12_data_i[15]), .QN(n2748) );
  INVX0 U37870 ( .IN(s10_data_i[15]), .QN(n2678) );
  INVX0 U37871 ( .IN(s6_data_i[15]), .QN(n2538) );
  INVX0 U37872 ( .IN(s0_data_i[15]), .QN(n2328) );
  INVX0 U37873 ( .IN(s12_data_i[16]), .QN(n2747) );
  INVX0 U37874 ( .IN(s10_data_i[16]), .QN(n2677) );
  INVX0 U37875 ( .IN(s6_data_i[16]), .QN(n2537) );
  INVX0 U37876 ( .IN(s0_data_i[16]), .QN(n2327) );
  INVX0 U37877 ( .IN(s12_data_i[17]), .QN(n2746) );
  INVX0 U37878 ( .IN(s10_data_i[17]), .QN(n2676) );
  INVX0 U37879 ( .IN(s6_data_i[17]), .QN(n2536) );
  INVX0 U37880 ( .IN(s0_data_i[17]), .QN(n2326) );
  INVX0 U37881 ( .IN(s12_data_i[18]), .QN(n2745) );
  INVX0 U37882 ( .IN(s10_data_i[18]), .QN(n2675) );
  INVX0 U37883 ( .IN(s6_data_i[18]), .QN(n2535) );
  INVX0 U37884 ( .IN(s0_data_i[18]), .QN(n2325) );
  INVX0 U37885 ( .IN(s12_data_i[19]), .QN(n2744) );
  INVX0 U37886 ( .IN(s10_data_i[19]), .QN(n2674) );
  INVX0 U37887 ( .IN(s6_data_i[19]), .QN(n2534) );
  INVX0 U37888 ( .IN(s0_data_i[19]), .QN(n2324) );
  INVX0 U37889 ( .IN(s12_data_i[20]), .QN(n2743) );
  INVX0 U37890 ( .IN(s10_data_i[20]), .QN(n2673) );
  INVX0 U37891 ( .IN(s6_data_i[20]), .QN(n2533) );
  INVX0 U37892 ( .IN(s0_data_i[20]), .QN(n2323) );
  INVX0 U37893 ( .IN(s12_data_i[21]), .QN(n2742) );
  INVX0 U37894 ( .IN(s10_data_i[21]), .QN(n2672) );
  INVX0 U37895 ( .IN(s6_data_i[21]), .QN(n2532) );
  INVX0 U37896 ( .IN(s0_data_i[21]), .QN(n2322) );
  INVX0 U37897 ( .IN(s12_data_i[22]), .QN(n2741) );
  INVX0 U37898 ( .IN(s10_data_i[22]), .QN(n2671) );
  INVX0 U37899 ( .IN(s6_data_i[22]), .QN(n2531) );
  INVX0 U37900 ( .IN(s0_data_i[22]), .QN(n2321) );
  INVX0 U37901 ( .IN(s12_data_i[23]), .QN(n2740) );
  INVX0 U37902 ( .IN(s10_data_i[23]), .QN(n2670) );
  INVX0 U37903 ( .IN(s6_data_i[23]), .QN(n2530) );
  INVX0 U37904 ( .IN(s0_data_i[23]), .QN(n2320) );
  INVX0 U37905 ( .IN(s12_data_i[24]), .QN(n2739) );
  INVX0 U37906 ( .IN(s10_data_i[24]), .QN(n2669) );
  INVX0 U37907 ( .IN(s6_data_i[24]), .QN(n2529) );
  INVX0 U37908 ( .IN(s0_data_i[24]), .QN(n2319) );
  INVX0 U37909 ( .IN(s12_data_i[25]), .QN(n2738) );
  INVX0 U37910 ( .IN(s10_data_i[25]), .QN(n2668) );
  INVX0 U37911 ( .IN(s6_data_i[25]), .QN(n2528) );
  INVX0 U37912 ( .IN(s0_data_i[25]), .QN(n2318) );
  INVX0 U37913 ( .IN(s12_data_i[26]), .QN(n2737) );
  INVX0 U37914 ( .IN(s10_data_i[26]), .QN(n2667) );
  INVX0 U37915 ( .IN(s6_data_i[26]), .QN(n2527) );
  INVX0 U37916 ( .IN(s0_data_i[26]), .QN(n2317) );
  INVX0 U37917 ( .IN(s12_data_i[27]), .QN(n2736) );
  INVX0 U37918 ( .IN(s10_data_i[27]), .QN(n2666) );
  INVX0 U37919 ( .IN(s6_data_i[27]), .QN(n2526) );
  INVX0 U37920 ( .IN(s0_data_i[27]), .QN(n2316) );
  INVX0 U37921 ( .IN(s12_data_i[28]), .QN(n2735) );
  INVX0 U37922 ( .IN(s10_data_i[28]), .QN(n2665) );
  INVX0 U37923 ( .IN(s6_data_i[28]), .QN(n2525) );
  INVX0 U37924 ( .IN(s0_data_i[28]), .QN(n2315) );
  INVX0 U37925 ( .IN(s12_data_i[29]), .QN(n2734) );
  INVX0 U37926 ( .IN(s10_data_i[29]), .QN(n2664) );
  INVX0 U37927 ( .IN(s6_data_i[29]), .QN(n2524) );
  INVX0 U37928 ( .IN(s0_data_i[29]), .QN(n2314) );
  INVX0 U37929 ( .IN(s12_data_i[30]), .QN(n2733) );
  INVX0 U37930 ( .IN(s10_data_i[30]), .QN(n2663) );
  INVX0 U37931 ( .IN(s6_data_i[30]), .QN(n2523) );
  INVX0 U37932 ( .IN(s0_data_i[30]), .QN(n2313) );
  INVX0 U37933 ( .IN(s12_data_i[31]), .QN(n2732) );
  INVX0 U37934 ( .IN(s10_data_i[31]), .QN(n2662) );
  INVX0 U37935 ( .IN(s6_data_i[31]), .QN(n2522) );
  INVX0 U37936 ( .IN(s0_data_i[31]), .QN(n2312) );
  NBUFFX2 U37937 ( .IN(n4502), .Q(n18430) );
  NAND3X0 U37938 ( .IN1(m5s15_cyc), .IN2(n19711), .IN3(s15_m5_cyc_r), .QN(
        n17102) );
  NAND3X0 U37939 ( .IN1(conf15_11_), .IN2(m5s15_cyc), .IN3(conf15_10_), .QN(
        n14183) );
  NAND3X0 U37940 ( .IN1(conf0_11_), .IN2(m5s0_cyc), .IN3(conf0_10_), .QN(
        n11744) );
  NAND3X0 U37941 ( .IN1(m5s0_cyc), .IN2(n18919), .IN3(s0_m5_cyc_r), .QN(n14487) );
  NAND3X0 U37942 ( .IN1(conf2_11_), .IN2(m5s2_cyc), .IN3(conf2_10_), .QN(
        n12364) );
  NAND3X0 U37943 ( .IN1(m5s2_cyc), .IN2(n19974), .IN3(s2_m5_cyc_r), .QN(n14467) );
  NAND3X0 U37944 ( .IN1(conf4_11_), .IN2(m5s4_cyc), .IN3(conf4_10_), .QN(
        n12982) );
  NAND3X0 U37945 ( .IN1(m5s4_cyc), .IN2(n20237), .IN3(test_so55), .QN(n14447)
         );
  NAND3X0 U37946 ( .IN1(conf7_11_), .IN2(test_so29), .IN3(conf7_10_), .QN(
        n13909) );
  NAND3X0 U37947 ( .IN1(test_so29), .IN2(n20633), .IN3(s7_m5_cyc_r), .QN(
        n14417) );
  NAND3X0 U37948 ( .IN1(conf1_11_), .IN2(test_so28), .IN3(conf1_10_), .QN(
        n12054) );
  NAND3X0 U37949 ( .IN1(test_so28), .IN2(n19843), .IN3(s1_m5_cyc_r), .QN(
        n14477) );
  NAND3X0 U37950 ( .IN1(conf3_11_), .IN2(m5s3_cyc), .IN3(conf3_10_), .QN(
        n12673) );
  NAND3X0 U37951 ( .IN1(m5s3_cyc), .IN2(n20105), .IN3(s3_m5_cyc_r), .QN(n14457) );
  NAND3X0 U37952 ( .IN1(conf5_11_), .IN2(m5s5_cyc), .IN3(conf5_10_), .QN(
        n13291) );
  NAND3X0 U37953 ( .IN1(m5s5_cyc), .IN2(n20369), .IN3(s5_m5_cyc_r), .QN(n14437) );
  OA22X1 U37954 ( .IN1(n14012), .IN2(n14013), .IN3(n14014), .IN4(n3398), .Q(
        n14005) );
  OA221X1 U37955 ( .IN1(n3093), .IN2(n14043), .IN3(n14044), .IN4(n14045), 
        .IN5(n14004), .Q(n14042) );
  OA22X1 U37956 ( .IN1(n14044), .IN2(n14021), .IN3(n14046), .IN4(n14048), .Q(
        n14066) );
  NAND2X0 U37957 ( .IN1(n14012), .IN2(n3254), .QN(n14031) );
  AND2X1 U37958 ( .IN1(n14044), .IN2(n14048), .Q(n14012) );
  NAND3X0 U37959 ( .IN1(conf8_11_), .IN2(m5s8_cyc), .IN3(conf8_10_), .QN(n9575) );
  NAND3X0 U37960 ( .IN1(m5s8_cyc), .IN2(n20765), .IN3(s8_m5_cyc_r), .QN(n14407) );
  NAND2X0 U37961 ( .IN1(n11583), .IN2(n3376), .QN(n11602) );
  AOI21X1 U37962 ( .IN1(n3540), .IN2(n11583), .IN3(n11624), .QN(n11603) );
  AND2X1 U37963 ( .IN1(n11615), .IN2(n11619), .Q(n11583) );
  NAND3X0 U37964 ( .IN1(conf10_11_), .IN2(m5s10_cyc), .IN3(conf10_10_), .QN(
        n10196) );
  NAND3X0 U37965 ( .IN1(m5s10_cyc), .IN2(n19051), .IN3(test_so78), .QN(n14387)
         );
  NAND2X0 U37966 ( .IN1(n12203), .IN2(n3360), .QN(n12222) );
  AOI21X1 U37967 ( .IN1(n3630), .IN2(n12203), .IN3(n12244), .QN(n12223) );
  AND2X1 U37968 ( .IN1(n12235), .IN2(n12239), .Q(n12203) );
  NAND3X0 U37969 ( .IN1(conf12_11_), .IN2(m5s12_cyc), .IN3(conf12_10_), .QN(
        n10815) );
  NAND3X0 U37970 ( .IN1(m5s12_cyc), .IN2(n19315), .IN3(s12_m5_cyc_r), .QN(
        n14367) );
  NAND2X0 U37971 ( .IN1(n12821), .IN2(n3344), .QN(n12840) );
  AOI21X1 U37972 ( .IN1(n3720), .IN2(n12821), .IN3(n12862), .QN(n12841) );
  AND2X1 U37973 ( .IN1(n12853), .IN2(n12857), .Q(n12821) );
  NAND3X0 U37974 ( .IN1(conf14_11_), .IN2(m5s14_cyc), .IN3(conf14_10_), .QN(
        n11434) );
  NAND3X0 U37975 ( .IN1(m5s14_cyc), .IN2(n19579), .IN3(s14_m5_cyc_r), .QN(
        n14347) );
  NAND2X0 U37976 ( .IN1(n13748), .IN2(n3320), .QN(n13767) );
  AOI21X1 U37977 ( .IN1(n3855), .IN2(n13748), .IN3(n13789), .QN(n13768) );
  AND2X1 U37978 ( .IN1(n13780), .IN2(n13784), .Q(n13748) );
  NAND3X0 U37979 ( .IN1(conf9_11_), .IN2(m5s9_cyc), .IN3(conf9_10_), .QN(n9886) );
  NAND3X0 U37980 ( .IN1(m5s9_cyc), .IN2(n20852), .IN3(s9_m5_cyc_r), .QN(n14397) );
  OA22X1 U37981 ( .IN1(n11893), .IN2(n11894), .IN3(n11895), .IN4(n3455), .Q(
        n11886) );
  OA221X1 U37982 ( .IN1(n3179), .IN2(n11924), .IN3(n11925), .IN4(n11926), 
        .IN5(n11885), .Q(n11923) );
  OA22X1 U37983 ( .IN1(n11925), .IN2(n11902), .IN3(n11927), .IN4(n11929), .Q(
        n11947) );
  NAND2X0 U37984 ( .IN1(n11893), .IN2(n3368), .QN(n11912) );
  AND2X1 U37985 ( .IN1(n11925), .IN2(n11929), .Q(n11893) );
  NAND3X0 U37986 ( .IN1(conf11_11_), .IN2(m5s11_cyc), .IN3(conf11_10_), .QN(
        n10506) );
  NAND3X0 U37987 ( .IN1(m5s11_cyc), .IN2(n19183), .IN3(s11_m5_cyc_r), .QN(
        n14377) );
  OA22X1 U37988 ( .IN1(n12512), .IN2(n12513), .IN3(n12514), .IN4(n3447), .Q(
        n12505) );
  OA221X1 U37989 ( .IN1(n3167), .IN2(n12543), .IN3(n12544), .IN4(n12545), 
        .IN5(n12504), .Q(n12542) );
  OA22X1 U37990 ( .IN1(n12544), .IN2(n12521), .IN3(n12546), .IN4(n12548), .Q(
        n12566) );
  NAND2X0 U37991 ( .IN1(n12512), .IN2(n3352), .QN(n12531) );
  AND2X1 U37992 ( .IN1(n12544), .IN2(n12548), .Q(n12512) );
  NAND3X0 U37993 ( .IN1(conf13_11_), .IN2(test_so30), .IN3(conf13_10_), .QN(
        n11125) );
  NAND3X0 U37994 ( .IN1(test_so30), .IN2(n19447), .IN3(s13_m5_cyc_r), .QN(
        n14357) );
  OA22X1 U37995 ( .IN1(n13130), .IN2(n13131), .IN3(n13132), .IN4(n3439), .Q(
        n13123) );
  OA221X1 U37996 ( .IN1(n3155), .IN2(n13161), .IN3(n13162), .IN4(n13163), 
        .IN5(n13122), .Q(n13160) );
  OA22X1 U37997 ( .IN1(n13162), .IN2(n13139), .IN3(n13164), .IN4(n13166), .Q(
        n13184) );
  NAND2X0 U37998 ( .IN1(n13130), .IN2(n3336), .QN(n13149) );
  AND2X1 U37999 ( .IN1(n13162), .IN2(n13166), .Q(n13130) );
  NAND3X0 U38000 ( .IN1(conf6_11_), .IN2(m5s6_cyc), .IN3(conf6_10_), .QN(
        n13600) );
  NAND3X0 U38001 ( .IN1(m5s6_cyc), .IN2(n20501), .IN3(s6_m5_cyc_r), .QN(n14427) );
  AND3X1 U38002 ( .IN1(n14012), .IN2(n3398), .IN3(n14055), .Q(n14057) );
  AO21X1 U38003 ( .IN1(n4217), .IN2(n14044), .IN3(n4214), .Q(n14053) );
  AOI21X1 U38004 ( .IN1(n4215), .IN2(n14012), .IN3(n14053), .QN(n14032) );
  OA22X1 U38005 ( .IN1(n9414), .IN2(n9415), .IN3(n9416), .IN4(n3427), .Q(n9407) );
  OA221X1 U38006 ( .IN1(n3137), .IN2(n9445), .IN3(n9446), .IN4(n9447), .IN5(
        n9406), .Q(n9444) );
  OA22X1 U38007 ( .IN1(n9446), .IN2(n9423), .IN3(n9448), .IN4(n9450), .Q(n9468) );
  AO21X1 U38008 ( .IN1(n3902), .IN2(n9446), .IN3(n3899), .Q(n9455) );
  AND3X1 U38009 ( .IN1(n9414), .IN2(n3427), .IN3(n9457), .Q(n9459) );
  NAND4X0 U38010 ( .IN1(m5s8_cyc), .IN2(n9329), .IN3(n9330), .IN4(n9331), .QN(
        n9320) );
  AO22X1 U38011 ( .IN1(n14328), .IN2(m5s8_cyc), .IN3(n14329), .IN4(n17831), 
        .Q(n17676) );
  AND3X1 U38012 ( .IN1(n9725), .IN2(n3423), .IN3(n9768), .Q(n9770) );
  AO21X1 U38013 ( .IN1(n3947), .IN2(n9757), .IN3(n3944), .Q(n9766) );
  AOI21X1 U38014 ( .IN1(n3945), .IN2(n9725), .IN3(n9766), .QN(n9745) );
  OA22X1 U38015 ( .IN1(n11583), .IN2(n11584), .IN3(n11585), .IN4(n3459), .Q(
        n11576) );
  OA221X1 U38016 ( .IN1(n3185), .IN2(n11614), .IN3(n11615), .IN4(n11616), 
        .IN5(n11575), .Q(n11613) );
  OA22X1 U38017 ( .IN1(n11615), .IN2(n11592), .IN3(n11617), .IN4(n11619), .Q(
        n11637) );
  AO21X1 U38018 ( .IN1(n3542), .IN2(n11615), .IN3(n3539), .Q(n11624) );
  AND3X1 U38019 ( .IN1(n11583), .IN2(n3459), .IN3(n11626), .Q(n11628) );
  NAND4X0 U38020 ( .IN1(m5s0_cyc), .IN2(n11498), .IN3(n11499), .IN4(n11500), 
        .QN(n11489) );
  AO22X1 U38021 ( .IN1(n14328), .IN2(m5s0_cyc), .IN3(n14329), .IN4(n18673), 
        .Q(n17668) );
  AND3X1 U38022 ( .IN1(n11893), .IN2(n3455), .IN3(n11936), .Q(n11938) );
  AO21X1 U38023 ( .IN1(n3587), .IN2(n11925), .IN3(n3584), .Q(n11934) );
  AOI21X1 U38024 ( .IN1(n3585), .IN2(n11893), .IN3(n11934), .QN(n11913) );
  OA22X1 U38025 ( .IN1(n10035), .IN2(n10036), .IN3(n10037), .IN4(n3419), .Q(
        n10028) );
  OA221X1 U38026 ( .IN1(n3125), .IN2(n10066), .IN3(n10067), .IN4(n10068), 
        .IN5(n10027), .Q(n10065) );
  OA22X1 U38027 ( .IN1(n10067), .IN2(n10044), .IN3(n10069), .IN4(n10071), .Q(
        n10089) );
  AO21X1 U38028 ( .IN1(n3992), .IN2(n10067), .IN3(n3989), .Q(n10076) );
  AND3X1 U38029 ( .IN1(n10035), .IN2(n3419), .IN3(n10078), .Q(n10080) );
  NAND4X0 U38030 ( .IN1(m5s10_cyc), .IN2(n9950), .IN3(n9951), .IN4(n9952), 
        .QN(n9941) );
  AO22X1 U38031 ( .IN1(n14328), .IN2(m5s10_cyc), .IN3(n14329), .IN4(n18697), 
        .Q(n17678) );
  AND3X1 U38032 ( .IN1(n10345), .IN2(n3415), .IN3(n10388), .Q(n10390) );
  AO21X1 U38033 ( .IN1(n4037), .IN2(n10377), .IN3(n4034), .Q(n10386) );
  AOI21X1 U38034 ( .IN1(n4035), .IN2(n10345), .IN3(n10386), .QN(n10365) );
  OA22X1 U38035 ( .IN1(n12203), .IN2(n12204), .IN3(n12205), .IN4(n3451), .Q(
        n12196) );
  OA221X1 U38036 ( .IN1(n3173), .IN2(n12234), .IN3(n12235), .IN4(n12236), 
        .IN5(n12195), .Q(n12233) );
  OA22X1 U38037 ( .IN1(n12235), .IN2(n12212), .IN3(n12237), .IN4(n12239), .Q(
        n12257) );
  AO21X1 U38038 ( .IN1(n3632), .IN2(n12235), .IN3(n3629), .Q(n12244) );
  AND3X1 U38039 ( .IN1(n12203), .IN2(n3451), .IN3(n12246), .Q(n12248) );
  NAND4X0 U38040 ( .IN1(m5s2_cyc), .IN2(n12118), .IN3(n12119), .IN4(n12120), 
        .QN(n12109) );
  AO22X1 U38041 ( .IN1(n14328), .IN2(m5s2_cyc), .IN3(n14329), .IN4(n17798), 
        .Q(n17670) );
  AND3X1 U38042 ( .IN1(n12512), .IN2(n3447), .IN3(n12555), .Q(n12557) );
  AO21X1 U38043 ( .IN1(n3677), .IN2(n12544), .IN3(n3674), .Q(n12553) );
  AOI21X1 U38044 ( .IN1(n3675), .IN2(n12512), .IN3(n12553), .QN(n12532) );
  OA22X1 U38045 ( .IN1(n10654), .IN2(n10655), .IN3(n10656), .IN4(n3411), .Q(
        n10647) );
  OA221X1 U38046 ( .IN1(n3113), .IN2(n10685), .IN3(n10686), .IN4(n10687), 
        .IN5(n10646), .Q(n10684) );
  OA22X1 U38047 ( .IN1(n10686), .IN2(n10663), .IN3(n10688), .IN4(n10690), .Q(
        n10708) );
  AO21X1 U38048 ( .IN1(n4082), .IN2(n10686), .IN3(n4079), .Q(n10695) );
  AND3X1 U38049 ( .IN1(n10654), .IN2(n3411), .IN3(n10697), .Q(n10699) );
  NAND4X0 U38050 ( .IN1(m5s12_cyc), .IN2(n10569), .IN3(n10570), .IN4(n10571), 
        .QN(n10560) );
  AO22X1 U38051 ( .IN1(n14328), .IN2(m5s12_cyc), .IN3(n14329), .IN4(n17811), 
        .Q(n17680) );
  AND3X1 U38052 ( .IN1(n10964), .IN2(n3407), .IN3(n11007), .Q(n11009) );
  AO21X1 U38053 ( .IN1(n4127), .IN2(n10996), .IN3(n4124), .Q(n11005) );
  AOI21X1 U38054 ( .IN1(n4125), .IN2(n10964), .IN3(n11005), .QN(n10984) );
  OA22X1 U38055 ( .IN1(n12821), .IN2(n12822), .IN3(n12823), .IN4(n3443), .Q(
        n12814) );
  OA221X1 U38056 ( .IN1(n3161), .IN2(n12852), .IN3(n12853), .IN4(n12854), 
        .IN5(n12813), .Q(n12851) );
  OA22X1 U38057 ( .IN1(n12853), .IN2(n12830), .IN3(n12855), .IN4(n12857), .Q(
        n12875) );
  AO21X1 U38058 ( .IN1(n3722), .IN2(n12853), .IN3(n3719), .Q(n12862) );
  AND3X1 U38059 ( .IN1(n12821), .IN2(n3443), .IN3(n12864), .Q(n12866) );
  NAND4X0 U38060 ( .IN1(m5s4_cyc), .IN2(n12736), .IN3(n12737), .IN4(n12738), 
        .QN(n12727) );
  AO22X1 U38061 ( .IN1(n14328), .IN2(m5s4_cyc), .IN3(n14329), .IN4(n17800), 
        .Q(n17672) );
  AND3X1 U38062 ( .IN1(n13130), .IN2(n3439), .IN3(n13173), .Q(n13175) );
  AO21X1 U38063 ( .IN1(n3767), .IN2(n13162), .IN3(n3764), .Q(n13171) );
  AOI21X1 U38064 ( .IN1(n3765), .IN2(n13130), .IN3(n13171), .QN(n13150) );
  OA22X1 U38065 ( .IN1(n11273), .IN2(n11274), .IN3(n11275), .IN4(n3403), .Q(
        n11266) );
  OA221X1 U38066 ( .IN1(n3101), .IN2(n11304), .IN3(n11305), .IN4(n11306), 
        .IN5(n11265), .Q(n11303) );
  OA22X1 U38067 ( .IN1(n11305), .IN2(n11282), .IN3(n11307), .IN4(n11309), .Q(
        n11327) );
  AO21X1 U38068 ( .IN1(n4172), .IN2(n11305), .IN3(n4169), .Q(n11314) );
  AND3X1 U38069 ( .IN1(n11273), .IN2(n3403), .IN3(n11316), .Q(n11318) );
  NAND4X0 U38070 ( .IN1(m5s14_cyc), .IN2(n11188), .IN3(n11189), .IN4(n11190), 
        .QN(n11179) );
  AO22X1 U38071 ( .IN1(n14328), .IN2(m5s14_cyc), .IN3(n14329), .IN4(n17827), 
        .Q(n17682) );
  AND3X1 U38072 ( .IN1(n13439), .IN2(n3435), .IN3(n13482), .Q(n13484) );
  AO21X1 U38073 ( .IN1(n3812), .IN2(n13471), .IN3(n3809), .Q(n13480) );
  AOI21X1 U38074 ( .IN1(n3810), .IN2(n13439), .IN3(n13480), .QN(n13459) );
  OA22X1 U38075 ( .IN1(n13748), .IN2(n13749), .IN3(n13750), .IN4(n3431), .Q(
        n13741) );
  OA221X1 U38076 ( .IN1(n3143), .IN2(n13779), .IN3(n13780), .IN4(n13781), 
        .IN5(n13740), .Q(n13778) );
  OA22X1 U38077 ( .IN1(n13780), .IN2(n13757), .IN3(n13782), .IN4(n13784), .Q(
        n13802) );
  AO21X1 U38078 ( .IN1(n3857), .IN2(n13780), .IN3(n3854), .Q(n13789) );
  AND3X1 U38079 ( .IN1(n13748), .IN2(n3431), .IN3(n13791), .Q(n13793) );
  NAND4X0 U38080 ( .IN1(test_so29), .IN2(n13663), .IN3(n13664), .IN4(n13665), 
        .QN(n13654) );
  AO22X1 U38081 ( .IN1(n14328), .IN2(test_so29), .IN3(n14329), .IN4(n17828), 
        .Q(n17675) );
  OR2X1 U38082 ( .IN1(n14070), .IN2(n18318), .Q(n14048) );
  NBUFFX2 U38083 ( .IN(m4s9_cyc), .Q(n18320) );
  NBUFFX2 U38084 ( .IN(m4s2_cyc), .Q(n18325) );
  NBUFFX2 U38085 ( .IN(m4s3_cyc), .Q(n18326) );
  NBUFFX2 U38086 ( .IN(m4s14_cyc), .Q(n18331) );
  NBUFFX2 U38087 ( .IN(m4s6_cyc), .Q(n18332) );
  NBUFFX2 U38088 ( .IN(m4s7_cyc), .Q(n18333) );
endmodule

